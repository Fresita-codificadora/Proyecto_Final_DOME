-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Oct 31 2024 19:51:41

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "anda_plis_2" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of anda_plis_2
entity anda_plis_2 is
port (
    leds : out std_logic_vector(13 downto 0);
    swit : in std_logic_vector(10 downto 0);
    uart_tx_o : out std_logic;
    uart_rx_i : in std_logic;
    clk : in std_logic;
    reset : in std_logic);
end anda_plis_2;

-- Architecture of anda_plis_2
-- View name is \INTERFACE\
architecture \INTERFACE\ of anda_plis_2 is

signal \N__39656\ : std_logic;
signal \N__39655\ : std_logic;
signal \N__39654\ : std_logic;
signal \N__39645\ : std_logic;
signal \N__39644\ : std_logic;
signal \N__39643\ : std_logic;
signal \N__39636\ : std_logic;
signal \N__39635\ : std_logic;
signal \N__39634\ : std_logic;
signal \N__39627\ : std_logic;
signal \N__39626\ : std_logic;
signal \N__39625\ : std_logic;
signal \N__39618\ : std_logic;
signal \N__39617\ : std_logic;
signal \N__39616\ : std_logic;
signal \N__39609\ : std_logic;
signal \N__39608\ : std_logic;
signal \N__39607\ : std_logic;
signal \N__39600\ : std_logic;
signal \N__39599\ : std_logic;
signal \N__39598\ : std_logic;
signal \N__39591\ : std_logic;
signal \N__39590\ : std_logic;
signal \N__39589\ : std_logic;
signal \N__39582\ : std_logic;
signal \N__39581\ : std_logic;
signal \N__39580\ : std_logic;
signal \N__39573\ : std_logic;
signal \N__39572\ : std_logic;
signal \N__39571\ : std_logic;
signal \N__39564\ : std_logic;
signal \N__39563\ : std_logic;
signal \N__39562\ : std_logic;
signal \N__39555\ : std_logic;
signal \N__39554\ : std_logic;
signal \N__39553\ : std_logic;
signal \N__39546\ : std_logic;
signal \N__39545\ : std_logic;
signal \N__39544\ : std_logic;
signal \N__39537\ : std_logic;
signal \N__39536\ : std_logic;
signal \N__39535\ : std_logic;
signal \N__39528\ : std_logic;
signal \N__39527\ : std_logic;
signal \N__39526\ : std_logic;
signal \N__39519\ : std_logic;
signal \N__39518\ : std_logic;
signal \N__39517\ : std_logic;
signal \N__39510\ : std_logic;
signal \N__39509\ : std_logic;
signal \N__39508\ : std_logic;
signal \N__39501\ : std_logic;
signal \N__39500\ : std_logic;
signal \N__39499\ : std_logic;
signal \N__39492\ : std_logic;
signal \N__39491\ : std_logic;
signal \N__39490\ : std_logic;
signal \N__39483\ : std_logic;
signal \N__39482\ : std_logic;
signal \N__39481\ : std_logic;
signal \N__39474\ : std_logic;
signal \N__39473\ : std_logic;
signal \N__39472\ : std_logic;
signal \N__39465\ : std_logic;
signal \N__39464\ : std_logic;
signal \N__39463\ : std_logic;
signal \N__39456\ : std_logic;
signal \N__39455\ : std_logic;
signal \N__39454\ : std_logic;
signal \N__39447\ : std_logic;
signal \N__39446\ : std_logic;
signal \N__39445\ : std_logic;
signal \N__39438\ : std_logic;
signal \N__39437\ : std_logic;
signal \N__39436\ : std_logic;
signal \N__39429\ : std_logic;
signal \N__39428\ : std_logic;
signal \N__39427\ : std_logic;
signal \N__39420\ : std_logic;
signal \N__39419\ : std_logic;
signal \N__39418\ : std_logic;
signal \N__39411\ : std_logic;
signal \N__39410\ : std_logic;
signal \N__39409\ : std_logic;
signal \N__39402\ : std_logic;
signal \N__39401\ : std_logic;
signal \N__39400\ : std_logic;
signal \N__39383\ : std_logic;
signal \N__39380\ : std_logic;
signal \N__39377\ : std_logic;
signal \N__39376\ : std_logic;
signal \N__39373\ : std_logic;
signal \N__39370\ : std_logic;
signal \N__39369\ : std_logic;
signal \N__39366\ : std_logic;
signal \N__39363\ : std_logic;
signal \N__39360\ : std_logic;
signal \N__39359\ : std_logic;
signal \N__39356\ : std_logic;
signal \N__39351\ : std_logic;
signal \N__39350\ : std_logic;
signal \N__39349\ : std_logic;
signal \N__39346\ : std_logic;
signal \N__39343\ : std_logic;
signal \N__39340\ : std_logic;
signal \N__39337\ : std_logic;
signal \N__39334\ : std_logic;
signal \N__39323\ : std_logic;
signal \N__39322\ : std_logic;
signal \N__39319\ : std_logic;
signal \N__39318\ : std_logic;
signal \N__39317\ : std_logic;
signal \N__39316\ : std_logic;
signal \N__39313\ : std_logic;
signal \N__39310\ : std_logic;
signal \N__39307\ : std_logic;
signal \N__39306\ : std_logic;
signal \N__39305\ : std_logic;
signal \N__39304\ : std_logic;
signal \N__39303\ : std_logic;
signal \N__39300\ : std_logic;
signal \N__39297\ : std_logic;
signal \N__39294\ : std_logic;
signal \N__39289\ : std_logic;
signal \N__39286\ : std_logic;
signal \N__39283\ : std_logic;
signal \N__39280\ : std_logic;
signal \N__39277\ : std_logic;
signal \N__39274\ : std_logic;
signal \N__39273\ : std_logic;
signal \N__39270\ : std_logic;
signal \N__39267\ : std_logic;
signal \N__39264\ : std_logic;
signal \N__39261\ : std_logic;
signal \N__39258\ : std_logic;
signal \N__39255\ : std_logic;
signal \N__39252\ : std_logic;
signal \N__39249\ : std_logic;
signal \N__39246\ : std_logic;
signal \N__39243\ : std_logic;
signal \N__39242\ : std_logic;
signal \N__39237\ : std_logic;
signal \N__39228\ : std_logic;
signal \N__39227\ : std_logic;
signal \N__39226\ : std_logic;
signal \N__39223\ : std_logic;
signal \N__39220\ : std_logic;
signal \N__39217\ : std_logic;
signal \N__39214\ : std_logic;
signal \N__39209\ : std_logic;
signal \N__39204\ : std_logic;
signal \N__39199\ : std_logic;
signal \N__39188\ : std_logic;
signal \N__39187\ : std_logic;
signal \N__39184\ : std_logic;
signal \N__39181\ : std_logic;
signal \N__39178\ : std_logic;
signal \N__39175\ : std_logic;
signal \N__39172\ : std_logic;
signal \N__39169\ : std_logic;
signal \N__39166\ : std_logic;
signal \N__39163\ : std_logic;
signal \N__39160\ : std_logic;
signal \N__39157\ : std_logic;
signal \N__39154\ : std_logic;
signal \N__39151\ : std_logic;
signal \N__39146\ : std_logic;
signal \N__39143\ : std_logic;
signal \N__39140\ : std_logic;
signal \N__39139\ : std_logic;
signal \N__39138\ : std_logic;
signal \N__39135\ : std_logic;
signal \N__39132\ : std_logic;
signal \N__39129\ : std_logic;
signal \N__39124\ : std_logic;
signal \N__39123\ : std_logic;
signal \N__39122\ : std_logic;
signal \N__39119\ : std_logic;
signal \N__39116\ : std_logic;
signal \N__39113\ : std_logic;
signal \N__39110\ : std_logic;
signal \N__39101\ : std_logic;
signal \N__39100\ : std_logic;
signal \N__39097\ : std_logic;
signal \N__39094\ : std_logic;
signal \N__39091\ : std_logic;
signal \N__39088\ : std_logic;
signal \N__39085\ : std_logic;
signal \N__39082\ : std_logic;
signal \N__39081\ : std_logic;
signal \N__39080\ : std_logic;
signal \N__39079\ : std_logic;
signal \N__39076\ : std_logic;
signal \N__39073\ : std_logic;
signal \N__39070\ : std_logic;
signal \N__39069\ : std_logic;
signal \N__39068\ : std_logic;
signal \N__39065\ : std_logic;
signal \N__39062\ : std_logic;
signal \N__39059\ : std_logic;
signal \N__39058\ : std_logic;
signal \N__39053\ : std_logic;
signal \N__39050\ : std_logic;
signal \N__39049\ : std_logic;
signal \N__39046\ : std_logic;
signal \N__39041\ : std_logic;
signal \N__39038\ : std_logic;
signal \N__39035\ : std_logic;
signal \N__39034\ : std_logic;
signal \N__39031\ : std_logic;
signal \N__39028\ : std_logic;
signal \N__39027\ : std_logic;
signal \N__39026\ : std_logic;
signal \N__39023\ : std_logic;
signal \N__39018\ : std_logic;
signal \N__39013\ : std_logic;
signal \N__39010\ : std_logic;
signal \N__39007\ : std_logic;
signal \N__39004\ : std_logic;
signal \N__39001\ : std_logic;
signal \N__38998\ : std_logic;
signal \N__38995\ : std_logic;
signal \N__38992\ : std_logic;
signal \N__38987\ : std_logic;
signal \N__38980\ : std_logic;
signal \N__38969\ : std_logic;
signal \N__38968\ : std_logic;
signal \N__38965\ : std_logic;
signal \N__38962\ : std_logic;
signal \N__38959\ : std_logic;
signal \N__38956\ : std_logic;
signal \N__38953\ : std_logic;
signal \N__38950\ : std_logic;
signal \N__38947\ : std_logic;
signal \N__38944\ : std_logic;
signal \N__38941\ : std_logic;
signal \N__38938\ : std_logic;
signal \N__38935\ : std_logic;
signal \N__38932\ : std_logic;
signal \N__38927\ : std_logic;
signal \N__38924\ : std_logic;
signal \N__38921\ : std_logic;
signal \N__38918\ : std_logic;
signal \N__38917\ : std_logic;
signal \N__38914\ : std_logic;
signal \N__38911\ : std_logic;
signal \N__38910\ : std_logic;
signal \N__38909\ : std_logic;
signal \N__38906\ : std_logic;
signal \N__38905\ : std_logic;
signal \N__38902\ : std_logic;
signal \N__38899\ : std_logic;
signal \N__38896\ : std_logic;
signal \N__38893\ : std_logic;
signal \N__38890\ : std_logic;
signal \N__38887\ : std_logic;
signal \N__38884\ : std_logic;
signal \N__38881\ : std_logic;
signal \N__38870\ : std_logic;
signal \N__38867\ : std_logic;
signal \N__38866\ : std_logic;
signal \N__38863\ : std_logic;
signal \N__38862\ : std_logic;
signal \N__38861\ : std_logic;
signal \N__38860\ : std_logic;
signal \N__38857\ : std_logic;
signal \N__38854\ : std_logic;
signal \N__38851\ : std_logic;
signal \N__38848\ : std_logic;
signal \N__38847\ : std_logic;
signal \N__38844\ : std_logic;
signal \N__38843\ : std_logic;
signal \N__38840\ : std_logic;
signal \N__38837\ : std_logic;
signal \N__38836\ : std_logic;
signal \N__38833\ : std_logic;
signal \N__38830\ : std_logic;
signal \N__38829\ : std_logic;
signal \N__38828\ : std_logic;
signal \N__38825\ : std_logic;
signal \N__38822\ : std_logic;
signal \N__38819\ : std_logic;
signal \N__38814\ : std_logic;
signal \N__38811\ : std_logic;
signal \N__38808\ : std_logic;
signal \N__38805\ : std_logic;
signal \N__38802\ : std_logic;
signal \N__38799\ : std_logic;
signal \N__38794\ : std_logic;
signal \N__38793\ : std_logic;
signal \N__38790\ : std_logic;
signal \N__38785\ : std_logic;
signal \N__38782\ : std_logic;
signal \N__38779\ : std_logic;
signal \N__38772\ : std_logic;
signal \N__38769\ : std_logic;
signal \N__38756\ : std_logic;
signal \N__38755\ : std_logic;
signal \N__38752\ : std_logic;
signal \N__38749\ : std_logic;
signal \N__38746\ : std_logic;
signal \N__38743\ : std_logic;
signal \N__38740\ : std_logic;
signal \N__38737\ : std_logic;
signal \N__38734\ : std_logic;
signal \N__38731\ : std_logic;
signal \N__38728\ : std_logic;
signal \N__38725\ : std_logic;
signal \N__38722\ : std_logic;
signal \N__38719\ : std_logic;
signal \N__38714\ : std_logic;
signal \N__38711\ : std_logic;
signal \N__38708\ : std_logic;
signal \N__38707\ : std_logic;
signal \N__38704\ : std_logic;
signal \N__38701\ : std_logic;
signal \N__38698\ : std_logic;
signal \N__38697\ : std_logic;
signal \N__38694\ : std_logic;
signal \N__38693\ : std_logic;
signal \N__38692\ : std_logic;
signal \N__38689\ : std_logic;
signal \N__38686\ : std_logic;
signal \N__38683\ : std_logic;
signal \N__38680\ : std_logic;
signal \N__38677\ : std_logic;
signal \N__38666\ : std_logic;
signal \N__38665\ : std_logic;
signal \N__38664\ : std_logic;
signal \N__38661\ : std_logic;
signal \N__38660\ : std_logic;
signal \N__38657\ : std_logic;
signal \N__38656\ : std_logic;
signal \N__38653\ : std_logic;
signal \N__38650\ : std_logic;
signal \N__38647\ : std_logic;
signal \N__38646\ : std_logic;
signal \N__38643\ : std_logic;
signal \N__38642\ : std_logic;
signal \N__38641\ : std_logic;
signal \N__38640\ : std_logic;
signal \N__38637\ : std_logic;
signal \N__38634\ : std_logic;
signal \N__38629\ : std_logic;
signal \N__38626\ : std_logic;
signal \N__38625\ : std_logic;
signal \N__38622\ : std_logic;
signal \N__38619\ : std_logic;
signal \N__38616\ : std_logic;
signal \N__38613\ : std_logic;
signal \N__38610\ : std_logic;
signal \N__38607\ : std_logic;
signal \N__38604\ : std_logic;
signal \N__38603\ : std_logic;
signal \N__38600\ : std_logic;
signal \N__38597\ : std_logic;
signal \N__38594\ : std_logic;
signal \N__38591\ : std_logic;
signal \N__38588\ : std_logic;
signal \N__38587\ : std_logic;
signal \N__38584\ : std_logic;
signal \N__38579\ : std_logic;
signal \N__38576\ : std_logic;
signal \N__38575\ : std_logic;
signal \N__38574\ : std_logic;
signal \N__38573\ : std_logic;
signal \N__38570\ : std_logic;
signal \N__38567\ : std_logic;
signal \N__38564\ : std_logic;
signal \N__38559\ : std_logic;
signal \N__38556\ : std_logic;
signal \N__38553\ : std_logic;
signal \N__38548\ : std_logic;
signal \N__38545\ : std_logic;
signal \N__38540\ : std_logic;
signal \N__38537\ : std_logic;
signal \N__38534\ : std_logic;
signal \N__38523\ : std_logic;
signal \N__38510\ : std_logic;
signal \N__38509\ : std_logic;
signal \N__38506\ : std_logic;
signal \N__38503\ : std_logic;
signal \N__38500\ : std_logic;
signal \N__38497\ : std_logic;
signal \N__38494\ : std_logic;
signal \N__38491\ : std_logic;
signal \N__38488\ : std_logic;
signal \N__38485\ : std_logic;
signal \N__38482\ : std_logic;
signal \N__38479\ : std_logic;
signal \N__38476\ : std_logic;
signal \N__38473\ : std_logic;
signal \N__38468\ : std_logic;
signal \N__38467\ : std_logic;
signal \N__38466\ : std_logic;
signal \N__38465\ : std_logic;
signal \N__38464\ : std_logic;
signal \N__38463\ : std_logic;
signal \N__38462\ : std_logic;
signal \N__38461\ : std_logic;
signal \N__38460\ : std_logic;
signal \N__38459\ : std_logic;
signal \N__38458\ : std_logic;
signal \N__38447\ : std_logic;
signal \N__38434\ : std_logic;
signal \N__38429\ : std_logic;
signal \N__38426\ : std_logic;
signal \N__38423\ : std_logic;
signal \N__38422\ : std_logic;
signal \N__38419\ : std_logic;
signal \N__38416\ : std_logic;
signal \N__38413\ : std_logic;
signal \N__38412\ : std_logic;
signal \N__38409\ : std_logic;
signal \N__38408\ : std_logic;
signal \N__38407\ : std_logic;
signal \N__38404\ : std_logic;
signal \N__38401\ : std_logic;
signal \N__38398\ : std_logic;
signal \N__38395\ : std_logic;
signal \N__38392\ : std_logic;
signal \N__38381\ : std_logic;
signal \N__38378\ : std_logic;
signal \N__38377\ : std_logic;
signal \N__38374\ : std_logic;
signal \N__38371\ : std_logic;
signal \N__38370\ : std_logic;
signal \N__38369\ : std_logic;
signal \N__38366\ : std_logic;
signal \N__38363\ : std_logic;
signal \N__38360\ : std_logic;
signal \N__38359\ : std_logic;
signal \N__38356\ : std_logic;
signal \N__38355\ : std_logic;
signal \N__38352\ : std_logic;
signal \N__38349\ : std_logic;
signal \N__38346\ : std_logic;
signal \N__38343\ : std_logic;
signal \N__38342\ : std_logic;
signal \N__38339\ : std_logic;
signal \N__38338\ : std_logic;
signal \N__38337\ : std_logic;
signal \N__38334\ : std_logic;
signal \N__38331\ : std_logic;
signal \N__38328\ : std_logic;
signal \N__38327\ : std_logic;
signal \N__38326\ : std_logic;
signal \N__38323\ : std_logic;
signal \N__38320\ : std_logic;
signal \N__38317\ : std_logic;
signal \N__38314\ : std_logic;
signal \N__38313\ : std_logic;
signal \N__38310\ : std_logic;
signal \N__38307\ : std_logic;
signal \N__38300\ : std_logic;
signal \N__38297\ : std_logic;
signal \N__38294\ : std_logic;
signal \N__38289\ : std_logic;
signal \N__38284\ : std_logic;
signal \N__38281\ : std_logic;
signal \N__38264\ : std_logic;
signal \N__38263\ : std_logic;
signal \N__38262\ : std_logic;
signal \N__38261\ : std_logic;
signal \N__38260\ : std_logic;
signal \N__38259\ : std_logic;
signal \N__38248\ : std_logic;
signal \N__38247\ : std_logic;
signal \N__38246\ : std_logic;
signal \N__38245\ : std_logic;
signal \N__38244\ : std_logic;
signal \N__38243\ : std_logic;
signal \N__38242\ : std_logic;
signal \N__38239\ : std_logic;
signal \N__38236\ : std_logic;
signal \N__38231\ : std_logic;
signal \N__38222\ : std_logic;
signal \N__38219\ : std_logic;
signal \N__38212\ : std_logic;
signal \N__38209\ : std_logic;
signal \N__38206\ : std_logic;
signal \N__38203\ : std_logic;
signal \N__38198\ : std_logic;
signal \N__38197\ : std_logic;
signal \N__38194\ : std_logic;
signal \N__38191\ : std_logic;
signal \N__38188\ : std_logic;
signal \N__38185\ : std_logic;
signal \N__38182\ : std_logic;
signal \N__38179\ : std_logic;
signal \N__38176\ : std_logic;
signal \N__38173\ : std_logic;
signal \N__38170\ : std_logic;
signal \N__38167\ : std_logic;
signal \N__38164\ : std_logic;
signal \N__38161\ : std_logic;
signal \N__38156\ : std_logic;
signal \N__38155\ : std_logic;
signal \N__38152\ : std_logic;
signal \N__38151\ : std_logic;
signal \N__38150\ : std_logic;
signal \N__38145\ : std_logic;
signal \N__38140\ : std_logic;
signal \N__38139\ : std_logic;
signal \N__38138\ : std_logic;
signal \N__38137\ : std_logic;
signal \N__38136\ : std_logic;
signal \N__38135\ : std_logic;
signal \N__38134\ : std_logic;
signal \N__38133\ : std_logic;
signal \N__38132\ : std_logic;
signal \N__38131\ : std_logic;
signal \N__38130\ : std_logic;
signal \N__38129\ : std_logic;
signal \N__38128\ : std_logic;
signal \N__38125\ : std_logic;
signal \N__38124\ : std_logic;
signal \N__38123\ : std_logic;
signal \N__38120\ : std_logic;
signal \N__38119\ : std_logic;
signal \N__38118\ : std_logic;
signal \N__38117\ : std_logic;
signal \N__38116\ : std_logic;
signal \N__38115\ : std_logic;
signal \N__38114\ : std_logic;
signal \N__38113\ : std_logic;
signal \N__38112\ : std_logic;
signal \N__38111\ : std_logic;
signal \N__38110\ : std_logic;
signal \N__38109\ : std_logic;
signal \N__38108\ : std_logic;
signal \N__38107\ : std_logic;
signal \N__38106\ : std_logic;
signal \N__38105\ : std_logic;
signal \N__38104\ : std_logic;
signal \N__38103\ : std_logic;
signal \N__38102\ : std_logic;
signal \N__38101\ : std_logic;
signal \N__38100\ : std_logic;
signal \N__38099\ : std_logic;
signal \N__38098\ : std_logic;
signal \N__38097\ : std_logic;
signal \N__38096\ : std_logic;
signal \N__38095\ : std_logic;
signal \N__38094\ : std_logic;
signal \N__38093\ : std_logic;
signal \N__38092\ : std_logic;
signal \N__38091\ : std_logic;
signal \N__38090\ : std_logic;
signal \N__38089\ : std_logic;
signal \N__38088\ : std_logic;
signal \N__38087\ : std_logic;
signal \N__38086\ : std_logic;
signal \N__38085\ : std_logic;
signal \N__38084\ : std_logic;
signal \N__38083\ : std_logic;
signal \N__38082\ : std_logic;
signal \N__38081\ : std_logic;
signal \N__38080\ : std_logic;
signal \N__38079\ : std_logic;
signal \N__38078\ : std_logic;
signal \N__38077\ : std_logic;
signal \N__38076\ : std_logic;
signal \N__38075\ : std_logic;
signal \N__38074\ : std_logic;
signal \N__38073\ : std_logic;
signal \N__38072\ : std_logic;
signal \N__38071\ : std_logic;
signal \N__38070\ : std_logic;
signal \N__38069\ : std_logic;
signal \N__38068\ : std_logic;
signal \N__38067\ : std_logic;
signal \N__38066\ : std_logic;
signal \N__38065\ : std_logic;
signal \N__38064\ : std_logic;
signal \N__38063\ : std_logic;
signal \N__38062\ : std_logic;
signal \N__38061\ : std_logic;
signal \N__38060\ : std_logic;
signal \N__38059\ : std_logic;
signal \N__38058\ : std_logic;
signal \N__38057\ : std_logic;
signal \N__38056\ : std_logic;
signal \N__38055\ : std_logic;
signal \N__38054\ : std_logic;
signal \N__38053\ : std_logic;
signal \N__38052\ : std_logic;
signal \N__38051\ : std_logic;
signal \N__38050\ : std_logic;
signal \N__38049\ : std_logic;
signal \N__38048\ : std_logic;
signal \N__38047\ : std_logic;
signal \N__38046\ : std_logic;
signal \N__38045\ : std_logic;
signal \N__38044\ : std_logic;
signal \N__38043\ : std_logic;
signal \N__38042\ : std_logic;
signal \N__38041\ : std_logic;
signal \N__38040\ : std_logic;
signal \N__37847\ : std_logic;
signal \N__37844\ : std_logic;
signal \N__37841\ : std_logic;
signal \N__37840\ : std_logic;
signal \N__37837\ : std_logic;
signal \N__37836\ : std_logic;
signal \N__37835\ : std_logic;
signal \N__37832\ : std_logic;
signal \N__37831\ : std_logic;
signal \N__37830\ : std_logic;
signal \N__37827\ : std_logic;
signal \N__37824\ : std_logic;
signal \N__37823\ : std_logic;
signal \N__37820\ : std_logic;
signal \N__37819\ : std_logic;
signal \N__37814\ : std_logic;
signal \N__37813\ : std_logic;
signal \N__37810\ : std_logic;
signal \N__37809\ : std_logic;
signal \N__37808\ : std_logic;
signal \N__37807\ : std_logic;
signal \N__37802\ : std_logic;
signal \N__37799\ : std_logic;
signal \N__37794\ : std_logic;
signal \N__37793\ : std_logic;
signal \N__37792\ : std_logic;
signal \N__37791\ : std_logic;
signal \N__37790\ : std_logic;
signal \N__37789\ : std_logic;
signal \N__37786\ : std_logic;
signal \N__37783\ : std_logic;
signal \N__37778\ : std_logic;
signal \N__37773\ : std_logic;
signal \N__37766\ : std_logic;
signal \N__37763\ : std_logic;
signal \N__37760\ : std_logic;
signal \N__37759\ : std_logic;
signal \N__37754\ : std_logic;
signal \N__37753\ : std_logic;
signal \N__37750\ : std_logic;
signal \N__37741\ : std_logic;
signal \N__37734\ : std_logic;
signal \N__37733\ : std_logic;
signal \N__37732\ : std_logic;
signal \N__37729\ : std_logic;
signal \N__37728\ : std_logic;
signal \N__37725\ : std_logic;
signal \N__37722\ : std_logic;
signal \N__37719\ : std_logic;
signal \N__37716\ : std_logic;
signal \N__37713\ : std_logic;
signal \N__37710\ : std_logic;
signal \N__37709\ : std_logic;
signal \N__37706\ : std_logic;
signal \N__37701\ : std_logic;
signal \N__37698\ : std_logic;
signal \N__37695\ : std_logic;
signal \N__37692\ : std_logic;
signal \N__37685\ : std_logic;
signal \N__37682\ : std_logic;
signal \N__37681\ : std_logic;
signal \N__37680\ : std_logic;
signal \N__37679\ : std_logic;
signal \N__37678\ : std_logic;
signal \N__37673\ : std_logic;
signal \N__37664\ : std_logic;
signal \N__37661\ : std_logic;
signal \N__37658\ : std_logic;
signal \N__37653\ : std_logic;
signal \N__37650\ : std_logic;
signal \N__37637\ : std_logic;
signal \N__37634\ : std_logic;
signal \N__37631\ : std_logic;
signal \N__37628\ : std_logic;
signal \N__37627\ : std_logic;
signal \N__37626\ : std_logic;
signal \N__37623\ : std_logic;
signal \N__37620\ : std_logic;
signal \N__37617\ : std_logic;
signal \N__37614\ : std_logic;
signal \N__37611\ : std_logic;
signal \N__37608\ : std_logic;
signal \N__37605\ : std_logic;
signal \N__37602\ : std_logic;
signal \N__37599\ : std_logic;
signal \N__37598\ : std_logic;
signal \N__37597\ : std_logic;
signal \N__37594\ : std_logic;
signal \N__37591\ : std_logic;
signal \N__37588\ : std_logic;
signal \N__37585\ : std_logic;
signal \N__37582\ : std_logic;
signal \N__37573\ : std_logic;
signal \N__37570\ : std_logic;
signal \N__37567\ : std_logic;
signal \N__37562\ : std_logic;
signal \N__37561\ : std_logic;
signal \N__37560\ : std_logic;
signal \N__37557\ : std_logic;
signal \N__37554\ : std_logic;
signal \N__37551\ : std_logic;
signal \N__37550\ : std_logic;
signal \N__37549\ : std_logic;
signal \N__37548\ : std_logic;
signal \N__37547\ : std_logic;
signal \N__37546\ : std_logic;
signal \N__37545\ : std_logic;
signal \N__37544\ : std_logic;
signal \N__37543\ : std_logic;
signal \N__37540\ : std_logic;
signal \N__37537\ : std_logic;
signal \N__37532\ : std_logic;
signal \N__37531\ : std_logic;
signal \N__37530\ : std_logic;
signal \N__37527\ : std_logic;
signal \N__37524\ : std_logic;
signal \N__37521\ : std_logic;
signal \N__37516\ : std_logic;
signal \N__37511\ : std_logic;
signal \N__37510\ : std_logic;
signal \N__37509\ : std_logic;
signal \N__37504\ : std_logic;
signal \N__37503\ : std_logic;
signal \N__37502\ : std_logic;
signal \N__37499\ : std_logic;
signal \N__37498\ : std_logic;
signal \N__37497\ : std_logic;
signal \N__37496\ : std_logic;
signal \N__37491\ : std_logic;
signal \N__37480\ : std_logic;
signal \N__37479\ : std_logic;
signal \N__37474\ : std_logic;
signal \N__37471\ : std_logic;
signal \N__37468\ : std_logic;
signal \N__37467\ : std_logic;
signal \N__37466\ : std_logic;
signal \N__37465\ : std_logic;
signal \N__37462\ : std_logic;
signal \N__37461\ : std_logic;
signal \N__37460\ : std_logic;
signal \N__37459\ : std_logic;
signal \N__37456\ : std_logic;
signal \N__37453\ : std_logic;
signal \N__37450\ : std_logic;
signal \N__37449\ : std_logic;
signal \N__37446\ : std_logic;
signal \N__37441\ : std_logic;
signal \N__37438\ : std_logic;
signal \N__37431\ : std_logic;
signal \N__37426\ : std_logic;
signal \N__37423\ : std_logic;
signal \N__37420\ : std_logic;
signal \N__37415\ : std_logic;
signal \N__37412\ : std_logic;
signal \N__37407\ : std_logic;
signal \N__37406\ : std_logic;
signal \N__37405\ : std_logic;
signal \N__37404\ : std_logic;
signal \N__37401\ : std_logic;
signal \N__37398\ : std_logic;
signal \N__37397\ : std_logic;
signal \N__37396\ : std_logic;
signal \N__37393\ : std_logic;
signal \N__37390\ : std_logic;
signal \N__37385\ : std_logic;
signal \N__37384\ : std_logic;
signal \N__37381\ : std_logic;
signal \N__37370\ : std_logic;
signal \N__37365\ : std_logic;
signal \N__37362\ : std_logic;
signal \N__37359\ : std_logic;
signal \N__37356\ : std_logic;
signal \N__37351\ : std_logic;
signal \N__37348\ : std_logic;
signal \N__37343\ : std_logic;
signal \N__37340\ : std_logic;
signal \N__37335\ : std_logic;
signal \N__37316\ : std_logic;
signal \N__37313\ : std_logic;
signal \N__37310\ : std_logic;
signal \N__37307\ : std_logic;
signal \N__37304\ : std_logic;
signal \N__37303\ : std_logic;
signal \N__37302\ : std_logic;
signal \N__37301\ : std_logic;
signal \N__37300\ : std_logic;
signal \N__37299\ : std_logic;
signal \N__37298\ : std_logic;
signal \N__37297\ : std_logic;
signal \N__37296\ : std_logic;
signal \N__37293\ : std_logic;
signal \N__37292\ : std_logic;
signal \N__37289\ : std_logic;
signal \N__37288\ : std_logic;
signal \N__37287\ : std_logic;
signal \N__37286\ : std_logic;
signal \N__37285\ : std_logic;
signal \N__37284\ : std_logic;
signal \N__37283\ : std_logic;
signal \N__37282\ : std_logic;
signal \N__37273\ : std_logic;
signal \N__37266\ : std_logic;
signal \N__37265\ : std_logic;
signal \N__37264\ : std_logic;
signal \N__37263\ : std_logic;
signal \N__37260\ : std_logic;
signal \N__37257\ : std_logic;
signal \N__37256\ : std_logic;
signal \N__37253\ : std_logic;
signal \N__37250\ : std_logic;
signal \N__37249\ : std_logic;
signal \N__37246\ : std_logic;
signal \N__37243\ : std_logic;
signal \N__37242\ : std_logic;
signal \N__37239\ : std_logic;
signal \N__37236\ : std_logic;
signal \N__37235\ : std_logic;
signal \N__37232\ : std_logic;
signal \N__37231\ : std_logic;
signal \N__37228\ : std_logic;
signal \N__37227\ : std_logic;
signal \N__37226\ : std_logic;
signal \N__37221\ : std_logic;
signal \N__37218\ : std_logic;
signal \N__37217\ : std_logic;
signal \N__37214\ : std_logic;
signal \N__37213\ : std_logic;
signal \N__37212\ : std_logic;
signal \N__37209\ : std_logic;
signal \N__37206\ : std_logic;
signal \N__37203\ : std_logic;
signal \N__37200\ : std_logic;
signal \N__37199\ : std_logic;
signal \N__37198\ : std_logic;
signal \N__37195\ : std_logic;
signal \N__37192\ : std_logic;
signal \N__37189\ : std_logic;
signal \N__37184\ : std_logic;
signal \N__37181\ : std_logic;
signal \N__37176\ : std_logic;
signal \N__37173\ : std_logic;
signal \N__37170\ : std_logic;
signal \N__37167\ : std_logic;
signal \N__37164\ : std_logic;
signal \N__37161\ : std_logic;
signal \N__37160\ : std_logic;
signal \N__37159\ : std_logic;
signal \N__37158\ : std_logic;
signal \N__37157\ : std_logic;
signal \N__37156\ : std_logic;
signal \N__37155\ : std_logic;
signal \N__37154\ : std_logic;
signal \N__37153\ : std_logic;
signal \N__37152\ : std_logic;
signal \N__37151\ : std_logic;
signal \N__37148\ : std_logic;
signal \N__37143\ : std_logic;
signal \N__37140\ : std_logic;
signal \N__37137\ : std_logic;
signal \N__37134\ : std_logic;
signal \N__37133\ : std_logic;
signal \N__37130\ : std_logic;
signal \N__37129\ : std_logic;
signal \N__37126\ : std_logic;
signal \N__37119\ : std_logic;
signal \N__37116\ : std_logic;
signal \N__37113\ : std_logic;
signal \N__37112\ : std_logic;
signal \N__37107\ : std_logic;
signal \N__37100\ : std_logic;
signal \N__37095\ : std_logic;
signal \N__37090\ : std_logic;
signal \N__37085\ : std_logic;
signal \N__37082\ : std_logic;
signal \N__37079\ : std_logic;
signal \N__37076\ : std_logic;
signal \N__37073\ : std_logic;
signal \N__37070\ : std_logic;
signal \N__37067\ : std_logic;
signal \N__37064\ : std_logic;
signal \N__37063\ : std_logic;
signal \N__37060\ : std_logic;
signal \N__37057\ : std_logic;
signal \N__37056\ : std_logic;
signal \N__37053\ : std_logic;
signal \N__37050\ : std_logic;
signal \N__37047\ : std_logic;
signal \N__37044\ : std_logic;
signal \N__37039\ : std_logic;
signal \N__37036\ : std_logic;
signal \N__37033\ : std_logic;
signal \N__37030\ : std_logic;
signal \N__37029\ : std_logic;
signal \N__37026\ : std_logic;
signal \N__37019\ : std_logic;
signal \N__37016\ : std_logic;
signal \N__37015\ : std_logic;
signal \N__37014\ : std_logic;
signal \N__37013\ : std_logic;
signal \N__37012\ : std_logic;
signal \N__37009\ : std_logic;
signal \N__37004\ : std_logic;
signal \N__36997\ : std_logic;
signal \N__36996\ : std_logic;
signal \N__36991\ : std_logic;
signal \N__36984\ : std_logic;
signal \N__36975\ : std_logic;
signal \N__36970\ : std_logic;
signal \N__36967\ : std_logic;
signal \N__36960\ : std_logic;
signal \N__36957\ : std_logic;
signal \N__36952\ : std_logic;
signal \N__36949\ : std_logic;
signal \N__36942\ : std_logic;
signal \N__36939\ : std_logic;
signal \N__36938\ : std_logic;
signal \N__36935\ : std_logic;
signal \N__36932\ : std_logic;
signal \N__36929\ : std_logic;
signal \N__36922\ : std_logic;
signal \N__36921\ : std_logic;
signal \N__36918\ : std_logic;
signal \N__36915\ : std_logic;
signal \N__36908\ : std_logic;
signal \N__36905\ : std_logic;
signal \N__36900\ : std_logic;
signal \N__36891\ : std_logic;
signal \N__36888\ : std_logic;
signal \N__36883\ : std_logic;
signal \N__36880\ : std_logic;
signal \N__36877\ : std_logic;
signal \N__36874\ : std_logic;
signal \N__36871\ : std_logic;
signal \N__36868\ : std_logic;
signal \N__36865\ : std_logic;
signal \N__36862\ : std_logic;
signal \N__36859\ : std_logic;
signal \N__36854\ : std_logic;
signal \N__36851\ : std_logic;
signal \N__36848\ : std_logic;
signal \N__36847\ : std_logic;
signal \N__36844\ : std_logic;
signal \N__36841\ : std_logic;
signal \N__36838\ : std_logic;
signal \N__36837\ : std_logic;
signal \N__36836\ : std_logic;
signal \N__36831\ : std_logic;
signal \N__36826\ : std_logic;
signal \N__36819\ : std_logic;
signal \N__36816\ : std_logic;
signal \N__36809\ : std_logic;
signal \N__36806\ : std_logic;
signal \N__36803\ : std_logic;
signal \N__36788\ : std_logic;
signal \N__36787\ : std_logic;
signal \N__36784\ : std_logic;
signal \N__36781\ : std_logic;
signal \N__36780\ : std_logic;
signal \N__36777\ : std_logic;
signal \N__36776\ : std_logic;
signal \N__36773\ : std_logic;
signal \N__36770\ : std_logic;
signal \N__36767\ : std_logic;
signal \N__36764\ : std_logic;
signal \N__36759\ : std_logic;
signal \N__36752\ : std_logic;
signal \N__36751\ : std_logic;
signal \N__36748\ : std_logic;
signal \N__36747\ : std_logic;
signal \N__36746\ : std_logic;
signal \N__36745\ : std_logic;
signal \N__36742\ : std_logic;
signal \N__36739\ : std_logic;
signal \N__36738\ : std_logic;
signal \N__36735\ : std_logic;
signal \N__36732\ : std_logic;
signal \N__36729\ : std_logic;
signal \N__36728\ : std_logic;
signal \N__36727\ : std_logic;
signal \N__36726\ : std_logic;
signal \N__36723\ : std_logic;
signal \N__36720\ : std_logic;
signal \N__36717\ : std_logic;
signal \N__36714\ : std_logic;
signal \N__36711\ : std_logic;
signal \N__36710\ : std_logic;
signal \N__36707\ : std_logic;
signal \N__36704\ : std_logic;
signal \N__36701\ : std_logic;
signal \N__36698\ : std_logic;
signal \N__36697\ : std_logic;
signal \N__36692\ : std_logic;
signal \N__36689\ : std_logic;
signal \N__36684\ : std_logic;
signal \N__36681\ : std_logic;
signal \N__36674\ : std_logic;
signal \N__36671\ : std_logic;
signal \N__36668\ : std_logic;
signal \N__36665\ : std_logic;
signal \N__36662\ : std_logic;
signal \N__36657\ : std_logic;
signal \N__36652\ : std_logic;
signal \N__36649\ : std_logic;
signal \N__36644\ : std_logic;
signal \N__36641\ : std_logic;
signal \N__36638\ : std_logic;
signal \N__36629\ : std_logic;
signal \N__36626\ : std_logic;
signal \N__36625\ : std_logic;
signal \N__36622\ : std_logic;
signal \N__36619\ : std_logic;
signal \N__36616\ : std_logic;
signal \N__36613\ : std_logic;
signal \N__36610\ : std_logic;
signal \N__36607\ : std_logic;
signal \N__36604\ : std_logic;
signal \N__36601\ : std_logic;
signal \N__36598\ : std_logic;
signal \N__36595\ : std_logic;
signal \N__36592\ : std_logic;
signal \N__36589\ : std_logic;
signal \N__36586\ : std_logic;
signal \N__36581\ : std_logic;
signal \N__36580\ : std_logic;
signal \N__36577\ : std_logic;
signal \N__36574\ : std_logic;
signal \N__36573\ : std_logic;
signal \N__36572\ : std_logic;
signal \N__36571\ : std_logic;
signal \N__36570\ : std_logic;
signal \N__36569\ : std_logic;
signal \N__36566\ : std_logic;
signal \N__36565\ : std_logic;
signal \N__36562\ : std_logic;
signal \N__36559\ : std_logic;
signal \N__36556\ : std_logic;
signal \N__36553\ : std_logic;
signal \N__36550\ : std_logic;
signal \N__36547\ : std_logic;
signal \N__36544\ : std_logic;
signal \N__36541\ : std_logic;
signal \N__36536\ : std_logic;
signal \N__36531\ : std_logic;
signal \N__36528\ : std_logic;
signal \N__36527\ : std_logic;
signal \N__36524\ : std_logic;
signal \N__36523\ : std_logic;
signal \N__36520\ : std_logic;
signal \N__36513\ : std_logic;
signal \N__36512\ : std_logic;
signal \N__36509\ : std_logic;
signal \N__36506\ : std_logic;
signal \N__36503\ : std_logic;
signal \N__36500\ : std_logic;
signal \N__36499\ : std_logic;
signal \N__36496\ : std_logic;
signal \N__36493\ : std_logic;
signal \N__36490\ : std_logic;
signal \N__36481\ : std_logic;
signal \N__36478\ : std_logic;
signal \N__36467\ : std_logic;
signal \N__36464\ : std_logic;
signal \N__36463\ : std_logic;
signal \N__36460\ : std_logic;
signal \N__36457\ : std_logic;
signal \N__36454\ : std_logic;
signal \N__36453\ : std_logic;
signal \N__36450\ : std_logic;
signal \N__36449\ : std_logic;
signal \N__36448\ : std_logic;
signal \N__36445\ : std_logic;
signal \N__36442\ : std_logic;
signal \N__36439\ : std_logic;
signal \N__36436\ : std_logic;
signal \N__36433\ : std_logic;
signal \N__36422\ : std_logic;
signal \N__36421\ : std_logic;
signal \N__36418\ : std_logic;
signal \N__36415\ : std_logic;
signal \N__36412\ : std_logic;
signal \N__36409\ : std_logic;
signal \N__36406\ : std_logic;
signal \N__36403\ : std_logic;
signal \N__36400\ : std_logic;
signal \N__36397\ : std_logic;
signal \N__36394\ : std_logic;
signal \N__36391\ : std_logic;
signal \N__36388\ : std_logic;
signal \N__36385\ : std_logic;
signal \N__36382\ : std_logic;
signal \N__36377\ : std_logic;
signal \N__36376\ : std_logic;
signal \N__36375\ : std_logic;
signal \N__36372\ : std_logic;
signal \N__36369\ : std_logic;
signal \N__36368\ : std_logic;
signal \N__36367\ : std_logic;
signal \N__36364\ : std_logic;
signal \N__36363\ : std_logic;
signal \N__36360\ : std_logic;
signal \N__36359\ : std_logic;
signal \N__36358\ : std_logic;
signal \N__36357\ : std_logic;
signal \N__36354\ : std_logic;
signal \N__36351\ : std_logic;
signal \N__36348\ : std_logic;
signal \N__36347\ : std_logic;
signal \N__36344\ : std_logic;
signal \N__36341\ : std_logic;
signal \N__36338\ : std_logic;
signal \N__36337\ : std_logic;
signal \N__36334\ : std_logic;
signal \N__36331\ : std_logic;
signal \N__36328\ : std_logic;
signal \N__36325\ : std_logic;
signal \N__36322\ : std_logic;
signal \N__36319\ : std_logic;
signal \N__36316\ : std_logic;
signal \N__36313\ : std_logic;
signal \N__36310\ : std_logic;
signal \N__36309\ : std_logic;
signal \N__36306\ : std_logic;
signal \N__36303\ : std_logic;
signal \N__36296\ : std_logic;
signal \N__36293\ : std_logic;
signal \N__36286\ : std_logic;
signal \N__36283\ : std_logic;
signal \N__36280\ : std_logic;
signal \N__36277\ : std_logic;
signal \N__36270\ : std_logic;
signal \N__36257\ : std_logic;
signal \N__36254\ : std_logic;
signal \N__36251\ : std_logic;
signal \N__36248\ : std_logic;
signal \N__36247\ : std_logic;
signal \N__36246\ : std_logic;
signal \N__36243\ : std_logic;
signal \N__36240\ : std_logic;
signal \N__36237\ : std_logic;
signal \N__36236\ : std_logic;
signal \N__36233\ : std_logic;
signal \N__36230\ : std_logic;
signal \N__36227\ : std_logic;
signal \N__36224\ : std_logic;
signal \N__36219\ : std_logic;
signal \N__36214\ : std_logic;
signal \N__36209\ : std_logic;
signal \N__36208\ : std_logic;
signal \N__36205\ : std_logic;
signal \N__36202\ : std_logic;
signal \N__36199\ : std_logic;
signal \N__36196\ : std_logic;
signal \N__36193\ : std_logic;
signal \N__36190\ : std_logic;
signal \N__36187\ : std_logic;
signal \N__36184\ : std_logic;
signal \N__36181\ : std_logic;
signal \N__36178\ : std_logic;
signal \N__36175\ : std_logic;
signal \N__36172\ : std_logic;
signal \N__36169\ : std_logic;
signal \N__36164\ : std_logic;
signal \N__36161\ : std_logic;
signal \N__36158\ : std_logic;
signal \N__36155\ : std_logic;
signal \N__36154\ : std_logic;
signal \N__36151\ : std_logic;
signal \N__36148\ : std_logic;
signal \N__36147\ : std_logic;
signal \N__36146\ : std_logic;
signal \N__36143\ : std_logic;
signal \N__36140\ : std_logic;
signal \N__36137\ : std_logic;
signal \N__36134\ : std_logic;
signal \N__36127\ : std_logic;
signal \N__36122\ : std_logic;
signal \N__36121\ : std_logic;
signal \N__36118\ : std_logic;
signal \N__36115\ : std_logic;
signal \N__36114\ : std_logic;
signal \N__36113\ : std_logic;
signal \N__36110\ : std_logic;
signal \N__36107\ : std_logic;
signal \N__36104\ : std_logic;
signal \N__36103\ : std_logic;
signal \N__36100\ : std_logic;
signal \N__36097\ : std_logic;
signal \N__36096\ : std_logic;
signal \N__36093\ : std_logic;
signal \N__36092\ : std_logic;
signal \N__36089\ : std_logic;
signal \N__36086\ : std_logic;
signal \N__36083\ : std_logic;
signal \N__36080\ : std_logic;
signal \N__36077\ : std_logic;
signal \N__36076\ : std_logic;
signal \N__36073\ : std_logic;
signal \N__36070\ : std_logic;
signal \N__36067\ : std_logic;
signal \N__36064\ : std_logic;
signal \N__36057\ : std_logic;
signal \N__36054\ : std_logic;
signal \N__36051\ : std_logic;
signal \N__36050\ : std_logic;
signal \N__36045\ : std_logic;
signal \N__36044\ : std_logic;
signal \N__36043\ : std_logic;
signal \N__36040\ : std_logic;
signal \N__36037\ : std_logic;
signal \N__36034\ : std_logic;
signal \N__36031\ : std_logic;
signal \N__36028\ : std_logic;
signal \N__36025\ : std_logic;
signal \N__36022\ : std_logic;
signal \N__36019\ : std_logic;
signal \N__36012\ : std_logic;
signal \N__35999\ : std_logic;
signal \N__35998\ : std_logic;
signal \N__35995\ : std_logic;
signal \N__35992\ : std_logic;
signal \N__35989\ : std_logic;
signal \N__35986\ : std_logic;
signal \N__35983\ : std_logic;
signal \N__35980\ : std_logic;
signal \N__35977\ : std_logic;
signal \N__35974\ : std_logic;
signal \N__35971\ : std_logic;
signal \N__35968\ : std_logic;
signal \N__35965\ : std_logic;
signal \N__35962\ : std_logic;
signal \N__35959\ : std_logic;
signal \N__35954\ : std_logic;
signal \N__35953\ : std_logic;
signal \N__35952\ : std_logic;
signal \N__35949\ : std_logic;
signal \N__35946\ : std_logic;
signal \N__35943\ : std_logic;
signal \N__35940\ : std_logic;
signal \N__35939\ : std_logic;
signal \N__35938\ : std_logic;
signal \N__35937\ : std_logic;
signal \N__35934\ : std_logic;
signal \N__35933\ : std_logic;
signal \N__35930\ : std_logic;
signal \N__35927\ : std_logic;
signal \N__35924\ : std_logic;
signal \N__35921\ : std_logic;
signal \N__35920\ : std_logic;
signal \N__35919\ : std_logic;
signal \N__35916\ : std_logic;
signal \N__35915\ : std_logic;
signal \N__35912\ : std_logic;
signal \N__35911\ : std_logic;
signal \N__35910\ : std_logic;
signal \N__35907\ : std_logic;
signal \N__35904\ : std_logic;
signal \N__35897\ : std_logic;
signal \N__35892\ : std_logic;
signal \N__35889\ : std_logic;
signal \N__35886\ : std_logic;
signal \N__35883\ : std_logic;
signal \N__35880\ : std_logic;
signal \N__35877\ : std_logic;
signal \N__35874\ : std_logic;
signal \N__35871\ : std_logic;
signal \N__35866\ : std_logic;
signal \N__35863\ : std_logic;
signal \N__35860\ : std_logic;
signal \N__35857\ : std_logic;
signal \N__35854\ : std_logic;
signal \N__35847\ : std_logic;
signal \N__35844\ : std_logic;
signal \N__35831\ : std_logic;
signal \N__35828\ : std_logic;
signal \N__35827\ : std_logic;
signal \N__35824\ : std_logic;
signal \N__35823\ : std_logic;
signal \N__35820\ : std_logic;
signal \N__35819\ : std_logic;
signal \N__35816\ : std_logic;
signal \N__35813\ : std_logic;
signal \N__35812\ : std_logic;
signal \N__35809\ : std_logic;
signal \N__35806\ : std_logic;
signal \N__35803\ : std_logic;
signal \N__35800\ : std_logic;
signal \N__35797\ : std_logic;
signal \N__35792\ : std_logic;
signal \N__35789\ : std_logic;
signal \N__35786\ : std_logic;
signal \N__35783\ : std_logic;
signal \N__35780\ : std_logic;
signal \N__35771\ : std_logic;
signal \N__35770\ : std_logic;
signal \N__35767\ : std_logic;
signal \N__35764\ : std_logic;
signal \N__35761\ : std_logic;
signal \N__35758\ : std_logic;
signal \N__35755\ : std_logic;
signal \N__35752\ : std_logic;
signal \N__35749\ : std_logic;
signal \N__35746\ : std_logic;
signal \N__35743\ : std_logic;
signal \N__35740\ : std_logic;
signal \N__35737\ : std_logic;
signal \N__35734\ : std_logic;
signal \N__35731\ : std_logic;
signal \N__35726\ : std_logic;
signal \N__35723\ : std_logic;
signal \N__35722\ : std_logic;
signal \N__35719\ : std_logic;
signal \N__35716\ : std_logic;
signal \N__35715\ : std_logic;
signal \N__35712\ : std_logic;
signal \N__35711\ : std_logic;
signal \N__35710\ : std_logic;
signal \N__35707\ : std_logic;
signal \N__35706\ : std_logic;
signal \N__35705\ : std_logic;
signal \N__35702\ : std_logic;
signal \N__35701\ : std_logic;
signal \N__35700\ : std_logic;
signal \N__35697\ : std_logic;
signal \N__35694\ : std_logic;
signal \N__35691\ : std_logic;
signal \N__35690\ : std_logic;
signal \N__35687\ : std_logic;
signal \N__35684\ : std_logic;
signal \N__35683\ : std_logic;
signal \N__35682\ : std_logic;
signal \N__35679\ : std_logic;
signal \N__35676\ : std_logic;
signal \N__35673\ : std_logic;
signal \N__35670\ : std_logic;
signal \N__35669\ : std_logic;
signal \N__35664\ : std_logic;
signal \N__35661\ : std_logic;
signal \N__35658\ : std_logic;
signal \N__35655\ : std_logic;
signal \N__35652\ : std_logic;
signal \N__35649\ : std_logic;
signal \N__35646\ : std_logic;
signal \N__35641\ : std_logic;
signal \N__35636\ : std_logic;
signal \N__35633\ : std_logic;
signal \N__35626\ : std_logic;
signal \N__35621\ : std_logic;
signal \N__35618\ : std_logic;
signal \N__35615\ : std_logic;
signal \N__35608\ : std_logic;
signal \N__35605\ : std_logic;
signal \N__35594\ : std_logic;
signal \N__35591\ : std_logic;
signal \N__35588\ : std_logic;
signal \N__35585\ : std_logic;
signal \N__35584\ : std_logic;
signal \N__35581\ : std_logic;
signal \N__35578\ : std_logic;
signal \N__35577\ : std_logic;
signal \N__35572\ : std_logic;
signal \N__35571\ : std_logic;
signal \N__35570\ : std_logic;
signal \N__35567\ : std_logic;
signal \N__35564\ : std_logic;
signal \N__35561\ : std_logic;
signal \N__35558\ : std_logic;
signal \N__35549\ : std_logic;
signal \N__35548\ : std_logic;
signal \N__35545\ : std_logic;
signal \N__35542\ : std_logic;
signal \N__35539\ : std_logic;
signal \N__35536\ : std_logic;
signal \N__35533\ : std_logic;
signal \N__35530\ : std_logic;
signal \N__35527\ : std_logic;
signal \N__35524\ : std_logic;
signal \N__35521\ : std_logic;
signal \N__35518\ : std_logic;
signal \N__35515\ : std_logic;
signal \N__35512\ : std_logic;
signal \N__35509\ : std_logic;
signal \N__35504\ : std_logic;
signal \N__35501\ : std_logic;
signal \N__35500\ : std_logic;
signal \N__35497\ : std_logic;
signal \N__35494\ : std_logic;
signal \N__35493\ : std_logic;
signal \N__35488\ : std_logic;
signal \N__35485\ : std_logic;
signal \N__35484\ : std_logic;
signal \N__35479\ : std_logic;
signal \N__35476\ : std_logic;
signal \N__35473\ : std_logic;
signal \N__35470\ : std_logic;
signal \N__35467\ : std_logic;
signal \N__35462\ : std_logic;
signal \N__35459\ : std_logic;
signal \N__35456\ : std_logic;
signal \N__35453\ : std_logic;
signal \N__35450\ : std_logic;
signal \N__35447\ : std_logic;
signal \N__35444\ : std_logic;
signal \N__35441\ : std_logic;
signal \N__35438\ : std_logic;
signal \N__35435\ : std_logic;
signal \N__35432\ : std_logic;
signal \N__35429\ : std_logic;
signal \N__35426\ : std_logic;
signal \N__35423\ : std_logic;
signal \N__35420\ : std_logic;
signal \N__35417\ : std_logic;
signal \N__35414\ : std_logic;
signal \N__35411\ : std_logic;
signal \N__35410\ : std_logic;
signal \N__35407\ : std_logic;
signal \N__35404\ : std_logic;
signal \N__35401\ : std_logic;
signal \N__35398\ : std_logic;
signal \N__35395\ : std_logic;
signal \N__35392\ : std_logic;
signal \N__35389\ : std_logic;
signal \N__35386\ : std_logic;
signal \N__35383\ : std_logic;
signal \N__35380\ : std_logic;
signal \N__35377\ : std_logic;
signal \N__35374\ : std_logic;
signal \N__35371\ : std_logic;
signal \N__35368\ : std_logic;
signal \N__35365\ : std_logic;
signal \N__35362\ : std_logic;
signal \N__35359\ : std_logic;
signal \N__35356\ : std_logic;
signal \N__35353\ : std_logic;
signal \N__35350\ : std_logic;
signal \N__35347\ : std_logic;
signal \N__35344\ : std_logic;
signal \N__35341\ : std_logic;
signal \N__35338\ : std_logic;
signal \N__35335\ : std_logic;
signal \N__35330\ : std_logic;
signal \N__35327\ : std_logic;
signal \N__35326\ : std_logic;
signal \N__35323\ : std_logic;
signal \N__35322\ : std_logic;
signal \N__35319\ : std_logic;
signal \N__35316\ : std_logic;
signal \N__35315\ : std_logic;
signal \N__35312\ : std_logic;
signal \N__35309\ : std_logic;
signal \N__35306\ : std_logic;
signal \N__35303\ : std_logic;
signal \N__35300\ : std_logic;
signal \N__35297\ : std_logic;
signal \N__35294\ : std_logic;
signal \N__35291\ : std_logic;
signal \N__35288\ : std_logic;
signal \N__35285\ : std_logic;
signal \N__35280\ : std_logic;
signal \N__35277\ : std_logic;
signal \N__35270\ : std_logic;
signal \N__35267\ : std_logic;
signal \N__35264\ : std_logic;
signal \N__35261\ : std_logic;
signal \N__35258\ : std_logic;
signal \N__35255\ : std_logic;
signal \N__35252\ : std_logic;
signal \N__35249\ : std_logic;
signal \N__35246\ : std_logic;
signal \N__35243\ : std_logic;
signal \N__35242\ : std_logic;
signal \N__35241\ : std_logic;
signal \N__35240\ : std_logic;
signal \N__35239\ : std_logic;
signal \N__35238\ : std_logic;
signal \N__35237\ : std_logic;
signal \N__35228\ : std_logic;
signal \N__35223\ : std_logic;
signal \N__35220\ : std_logic;
signal \N__35219\ : std_logic;
signal \N__35218\ : std_logic;
signal \N__35217\ : std_logic;
signal \N__35216\ : std_logic;
signal \N__35215\ : std_logic;
signal \N__35210\ : std_logic;
signal \N__35209\ : std_logic;
signal \N__35208\ : std_logic;
signal \N__35207\ : std_logic;
signal \N__35204\ : std_logic;
signal \N__35197\ : std_logic;
signal \N__35196\ : std_logic;
signal \N__35193\ : std_logic;
signal \N__35190\ : std_logic;
signal \N__35189\ : std_logic;
signal \N__35188\ : std_logic;
signal \N__35187\ : std_logic;
signal \N__35186\ : std_logic;
signal \N__35185\ : std_logic;
signal \N__35182\ : std_logic;
signal \N__35179\ : std_logic;
signal \N__35176\ : std_logic;
signal \N__35173\ : std_logic;
signal \N__35172\ : std_logic;
signal \N__35167\ : std_logic;
signal \N__35166\ : std_logic;
signal \N__35163\ : std_logic;
signal \N__35160\ : std_logic;
signal \N__35157\ : std_logic;
signal \N__35148\ : std_logic;
signal \N__35145\ : std_logic;
signal \N__35140\ : std_logic;
signal \N__35137\ : std_logic;
signal \N__35134\ : std_logic;
signal \N__35131\ : std_logic;
signal \N__35128\ : std_logic;
signal \N__35125\ : std_logic;
signal \N__35122\ : std_logic;
signal \N__35119\ : std_logic;
signal \N__35116\ : std_logic;
signal \N__35113\ : std_logic;
signal \N__35108\ : std_logic;
signal \N__35105\ : std_logic;
signal \N__35100\ : std_logic;
signal \N__35095\ : std_logic;
signal \N__35092\ : std_logic;
signal \N__35075\ : std_logic;
signal \N__35072\ : std_logic;
signal \N__35069\ : std_logic;
signal \N__35066\ : std_logic;
signal \N__35063\ : std_logic;
signal \N__35060\ : std_logic;
signal \N__35057\ : std_logic;
signal \N__35056\ : std_logic;
signal \N__35053\ : std_logic;
signal \N__35050\ : std_logic;
signal \N__35047\ : std_logic;
signal \N__35044\ : std_logic;
signal \N__35041\ : std_logic;
signal \N__35038\ : std_logic;
signal \N__35035\ : std_logic;
signal \N__35032\ : std_logic;
signal \N__35029\ : std_logic;
signal \N__35026\ : std_logic;
signal \N__35023\ : std_logic;
signal \N__35020\ : std_logic;
signal \N__35017\ : std_logic;
signal \N__35014\ : std_logic;
signal \N__35011\ : std_logic;
signal \N__35008\ : std_logic;
signal \N__35005\ : std_logic;
signal \N__35002\ : std_logic;
signal \N__34999\ : std_logic;
signal \N__34996\ : std_logic;
signal \N__34993\ : std_logic;
signal \N__34990\ : std_logic;
signal \N__34987\ : std_logic;
signal \N__34984\ : std_logic;
signal \N__34979\ : std_logic;
signal \N__34976\ : std_logic;
signal \N__34975\ : std_logic;
signal \N__34974\ : std_logic;
signal \N__34973\ : std_logic;
signal \N__34970\ : std_logic;
signal \N__34967\ : std_logic;
signal \N__34966\ : std_logic;
signal \N__34963\ : std_logic;
signal \N__34960\ : std_logic;
signal \N__34957\ : std_logic;
signal \N__34954\ : std_logic;
signal \N__34951\ : std_logic;
signal \N__34948\ : std_logic;
signal \N__34945\ : std_logic;
signal \N__34942\ : std_logic;
signal \N__34939\ : std_logic;
signal \N__34936\ : std_logic;
signal \N__34931\ : std_logic;
signal \N__34928\ : std_logic;
signal \N__34921\ : std_logic;
signal \N__34916\ : std_logic;
signal \N__34913\ : std_logic;
signal \N__34910\ : std_logic;
signal \N__34909\ : std_logic;
signal \N__34908\ : std_logic;
signal \N__34907\ : std_logic;
signal \N__34904\ : std_logic;
signal \N__34903\ : std_logic;
signal \N__34900\ : std_logic;
signal \N__34897\ : std_logic;
signal \N__34894\ : std_logic;
signal \N__34891\ : std_logic;
signal \N__34888\ : std_logic;
signal \N__34885\ : std_logic;
signal \N__34874\ : std_logic;
signal \N__34871\ : std_logic;
signal \N__34870\ : std_logic;
signal \N__34867\ : std_logic;
signal \N__34866\ : std_logic;
signal \N__34865\ : std_logic;
signal \N__34862\ : std_logic;
signal \N__34859\ : std_logic;
signal \N__34856\ : std_logic;
signal \N__34853\ : std_logic;
signal \N__34844\ : std_logic;
signal \N__34841\ : std_logic;
signal \N__34840\ : std_logic;
signal \N__34839\ : std_logic;
signal \N__34838\ : std_logic;
signal \N__34835\ : std_logic;
signal \N__34832\ : std_logic;
signal \N__34829\ : std_logic;
signal \N__34826\ : std_logic;
signal \N__34825\ : std_logic;
signal \N__34822\ : std_logic;
signal \N__34819\ : std_logic;
signal \N__34816\ : std_logic;
signal \N__34813\ : std_logic;
signal \N__34810\ : std_logic;
signal \N__34807\ : std_logic;
signal \N__34804\ : std_logic;
signal \N__34801\ : std_logic;
signal \N__34798\ : std_logic;
signal \N__34795\ : std_logic;
signal \N__34792\ : std_logic;
signal \N__34787\ : std_logic;
signal \N__34782\ : std_logic;
signal \N__34775\ : std_logic;
signal \N__34772\ : std_logic;
signal \N__34769\ : std_logic;
signal \N__34766\ : std_logic;
signal \N__34765\ : std_logic;
signal \N__34764\ : std_logic;
signal \N__34763\ : std_logic;
signal \N__34762\ : std_logic;
signal \N__34761\ : std_logic;
signal \N__34758\ : std_logic;
signal \N__34755\ : std_logic;
signal \N__34752\ : std_logic;
signal \N__34747\ : std_logic;
signal \N__34746\ : std_logic;
signal \N__34745\ : std_logic;
signal \N__34742\ : std_logic;
signal \N__34741\ : std_logic;
signal \N__34738\ : std_logic;
signal \N__34731\ : std_logic;
signal \N__34728\ : std_logic;
signal \N__34727\ : std_logic;
signal \N__34726\ : std_logic;
signal \N__34725\ : std_logic;
signal \N__34722\ : std_logic;
signal \N__34719\ : std_logic;
signal \N__34716\ : std_logic;
signal \N__34713\ : std_logic;
signal \N__34710\ : std_logic;
signal \N__34707\ : std_logic;
signal \N__34706\ : std_logic;
signal \N__34703\ : std_logic;
signal \N__34698\ : std_logic;
signal \N__34695\ : std_logic;
signal \N__34694\ : std_logic;
signal \N__34691\ : std_logic;
signal \N__34688\ : std_logic;
signal \N__34681\ : std_logic;
signal \N__34676\ : std_logic;
signal \N__34673\ : std_logic;
signal \N__34670\ : std_logic;
signal \N__34667\ : std_logic;
signal \N__34652\ : std_logic;
signal \N__34649\ : std_logic;
signal \N__34646\ : std_logic;
signal \N__34643\ : std_logic;
signal \N__34642\ : std_logic;
signal \N__34639\ : std_logic;
signal \N__34636\ : std_logic;
signal \N__34633\ : std_logic;
signal \N__34630\ : std_logic;
signal \N__34629\ : std_logic;
signal \N__34628\ : std_logic;
signal \N__34627\ : std_logic;
signal \N__34626\ : std_logic;
signal \N__34625\ : std_logic;
signal \N__34624\ : std_logic;
signal \N__34623\ : std_logic;
signal \N__34620\ : std_logic;
signal \N__34617\ : std_logic;
signal \N__34610\ : std_logic;
signal \N__34607\ : std_logic;
signal \N__34604\ : std_logic;
signal \N__34599\ : std_logic;
signal \N__34592\ : std_logic;
signal \N__34589\ : std_logic;
signal \N__34588\ : std_logic;
signal \N__34583\ : std_logic;
signal \N__34582\ : std_logic;
signal \N__34579\ : std_logic;
signal \N__34576\ : std_logic;
signal \N__34573\ : std_logic;
signal \N__34570\ : std_logic;
signal \N__34567\ : std_logic;
signal \N__34556\ : std_logic;
signal \N__34553\ : std_logic;
signal \N__34550\ : std_logic;
signal \N__34549\ : std_logic;
signal \N__34546\ : std_logic;
signal \N__34545\ : std_logic;
signal \N__34542\ : std_logic;
signal \N__34539\ : std_logic;
signal \N__34536\ : std_logic;
signal \N__34529\ : std_logic;
signal \N__34528\ : std_logic;
signal \N__34527\ : std_logic;
signal \N__34526\ : std_logic;
signal \N__34525\ : std_logic;
signal \N__34524\ : std_logic;
signal \N__34523\ : std_logic;
signal \N__34522\ : std_logic;
signal \N__34521\ : std_logic;
signal \N__34520\ : std_logic;
signal \N__34519\ : std_logic;
signal \N__34518\ : std_logic;
signal \N__34517\ : std_logic;
signal \N__34516\ : std_logic;
signal \N__34515\ : std_logic;
signal \N__34514\ : std_logic;
signal \N__34513\ : std_logic;
signal \N__34512\ : std_logic;
signal \N__34511\ : std_logic;
signal \N__34510\ : std_logic;
signal \N__34509\ : std_logic;
signal \N__34508\ : std_logic;
signal \N__34507\ : std_logic;
signal \N__34506\ : std_logic;
signal \N__34505\ : std_logic;
signal \N__34504\ : std_logic;
signal \N__34503\ : std_logic;
signal \N__34502\ : std_logic;
signal \N__34501\ : std_logic;
signal \N__34500\ : std_logic;
signal \N__34499\ : std_logic;
signal \N__34498\ : std_logic;
signal \N__34497\ : std_logic;
signal \N__34496\ : std_logic;
signal \N__34495\ : std_logic;
signal \N__34494\ : std_logic;
signal \N__34493\ : std_logic;
signal \N__34492\ : std_logic;
signal \N__34491\ : std_logic;
signal \N__34490\ : std_logic;
signal \N__34489\ : std_logic;
signal \N__34488\ : std_logic;
signal \N__34487\ : std_logic;
signal \N__34486\ : std_logic;
signal \N__34485\ : std_logic;
signal \N__34484\ : std_logic;
signal \N__34483\ : std_logic;
signal \N__34482\ : std_logic;
signal \N__34481\ : std_logic;
signal \N__34480\ : std_logic;
signal \N__34479\ : std_logic;
signal \N__34478\ : std_logic;
signal \N__34477\ : std_logic;
signal \N__34476\ : std_logic;
signal \N__34475\ : std_logic;
signal \N__34474\ : std_logic;
signal \N__34473\ : std_logic;
signal \N__34472\ : std_logic;
signal \N__34471\ : std_logic;
signal \N__34470\ : std_logic;
signal \N__34469\ : std_logic;
signal \N__34468\ : std_logic;
signal \N__34467\ : std_logic;
signal \N__34466\ : std_logic;
signal \N__34465\ : std_logic;
signal \N__34464\ : std_logic;
signal \N__34463\ : std_logic;
signal \N__34462\ : std_logic;
signal \N__34461\ : std_logic;
signal \N__34460\ : std_logic;
signal \N__34459\ : std_logic;
signal \N__34458\ : std_logic;
signal \N__34457\ : std_logic;
signal \N__34456\ : std_logic;
signal \N__34455\ : std_logic;
signal \N__34454\ : std_logic;
signal \N__34453\ : std_logic;
signal \N__34452\ : std_logic;
signal \N__34451\ : std_logic;
signal \N__34450\ : std_logic;
signal \N__34449\ : std_logic;
signal \N__34448\ : std_logic;
signal \N__34447\ : std_logic;
signal \N__34446\ : std_logic;
signal \N__34445\ : std_logic;
signal \N__34444\ : std_logic;
signal \N__34443\ : std_logic;
signal \N__34442\ : std_logic;
signal \N__34441\ : std_logic;
signal \N__34440\ : std_logic;
signal \N__34439\ : std_logic;
signal \N__34438\ : std_logic;
signal \N__34437\ : std_logic;
signal \N__34436\ : std_logic;
signal \N__34435\ : std_logic;
signal \N__34434\ : std_logic;
signal \N__34433\ : std_logic;
signal \N__34432\ : std_logic;
signal \N__34431\ : std_logic;
signal \N__34430\ : std_logic;
signal \N__34429\ : std_logic;
signal \N__34428\ : std_logic;
signal \N__34427\ : std_logic;
signal \N__34426\ : std_logic;
signal \N__34425\ : std_logic;
signal \N__34424\ : std_logic;
signal \N__34423\ : std_logic;
signal \N__34422\ : std_logic;
signal \N__34421\ : std_logic;
signal \N__34420\ : std_logic;
signal \N__34419\ : std_logic;
signal \N__34418\ : std_logic;
signal \N__34417\ : std_logic;
signal \N__34416\ : std_logic;
signal \N__34415\ : std_logic;
signal \N__34414\ : std_logic;
signal \N__34413\ : std_logic;
signal \N__34412\ : std_logic;
signal \N__34411\ : std_logic;
signal \N__34410\ : std_logic;
signal \N__34409\ : std_logic;
signal \N__34408\ : std_logic;
signal \N__34407\ : std_logic;
signal \N__34406\ : std_logic;
signal \N__34405\ : std_logic;
signal \N__34404\ : std_logic;
signal \N__34403\ : std_logic;
signal \N__34402\ : std_logic;
signal \N__34401\ : std_logic;
signal \N__34400\ : std_logic;
signal \N__34399\ : std_logic;
signal \N__34398\ : std_logic;
signal \N__34397\ : std_logic;
signal \N__34396\ : std_logic;
signal \N__34395\ : std_logic;
signal \N__34394\ : std_logic;
signal \N__34393\ : std_logic;
signal \N__34392\ : std_logic;
signal \N__34391\ : std_logic;
signal \N__34390\ : std_logic;
signal \N__34389\ : std_logic;
signal \N__34388\ : std_logic;
signal \N__34387\ : std_logic;
signal \N__34386\ : std_logic;
signal \N__34385\ : std_logic;
signal \N__34384\ : std_logic;
signal \N__34383\ : std_logic;
signal \N__34382\ : std_logic;
signal \N__34381\ : std_logic;
signal \N__34380\ : std_logic;
signal \N__34379\ : std_logic;
signal \N__34378\ : std_logic;
signal \N__34377\ : std_logic;
signal \N__34376\ : std_logic;
signal \N__34375\ : std_logic;
signal \N__34374\ : std_logic;
signal \N__34373\ : std_logic;
signal \N__34372\ : std_logic;
signal \N__34371\ : std_logic;
signal \N__34052\ : std_logic;
signal \N__34049\ : std_logic;
signal \N__34046\ : std_logic;
signal \N__34043\ : std_logic;
signal \N__34040\ : std_logic;
signal \N__34037\ : std_logic;
signal \N__34034\ : std_logic;
signal \N__34031\ : std_logic;
signal \N__34028\ : std_logic;
signal \N__34025\ : std_logic;
signal \N__34022\ : std_logic;
signal \N__34019\ : std_logic;
signal \N__34016\ : std_logic;
signal \N__34013\ : std_logic;
signal \N__34010\ : std_logic;
signal \N__34009\ : std_logic;
signal \N__34006\ : std_logic;
signal \N__34003\ : std_logic;
signal \N__34000\ : std_logic;
signal \N__33997\ : std_logic;
signal \N__33994\ : std_logic;
signal \N__33991\ : std_logic;
signal \N__33988\ : std_logic;
signal \N__33985\ : std_logic;
signal \N__33982\ : std_logic;
signal \N__33979\ : std_logic;
signal \N__33976\ : std_logic;
signal \N__33973\ : std_logic;
signal \N__33970\ : std_logic;
signal \N__33967\ : std_logic;
signal \N__33964\ : std_logic;
signal \N__33961\ : std_logic;
signal \N__33958\ : std_logic;
signal \N__33955\ : std_logic;
signal \N__33952\ : std_logic;
signal \N__33949\ : std_logic;
signal \N__33946\ : std_logic;
signal \N__33943\ : std_logic;
signal \N__33940\ : std_logic;
signal \N__33937\ : std_logic;
signal \N__33934\ : std_logic;
signal \N__33929\ : std_logic;
signal \N__33926\ : std_logic;
signal \N__33923\ : std_logic;
signal \N__33920\ : std_logic;
signal \N__33917\ : std_logic;
signal \N__33914\ : std_logic;
signal \N__33911\ : std_logic;
signal \N__33908\ : std_logic;
signal \N__33905\ : std_logic;
signal \N__33902\ : std_logic;
signal \N__33899\ : std_logic;
signal \N__33896\ : std_logic;
signal \N__33893\ : std_logic;
signal \N__33892\ : std_logic;
signal \N__33889\ : std_logic;
signal \N__33886\ : std_logic;
signal \N__33883\ : std_logic;
signal \N__33880\ : std_logic;
signal \N__33877\ : std_logic;
signal \N__33874\ : std_logic;
signal \N__33871\ : std_logic;
signal \N__33868\ : std_logic;
signal \N__33865\ : std_logic;
signal \N__33862\ : std_logic;
signal \N__33859\ : std_logic;
signal \N__33856\ : std_logic;
signal \N__33853\ : std_logic;
signal \N__33850\ : std_logic;
signal \N__33847\ : std_logic;
signal \N__33844\ : std_logic;
signal \N__33841\ : std_logic;
signal \N__33838\ : std_logic;
signal \N__33835\ : std_logic;
signal \N__33832\ : std_logic;
signal \N__33829\ : std_logic;
signal \N__33826\ : std_logic;
signal \N__33823\ : std_logic;
signal \N__33820\ : std_logic;
signal \N__33817\ : std_logic;
signal \N__33812\ : std_logic;
signal \N__33809\ : std_logic;
signal \N__33806\ : std_logic;
signal \N__33803\ : std_logic;
signal \N__33800\ : std_logic;
signal \N__33797\ : std_logic;
signal \N__33794\ : std_logic;
signal \N__33791\ : std_logic;
signal \N__33788\ : std_logic;
signal \N__33785\ : std_logic;
signal \N__33782\ : std_logic;
signal \N__33779\ : std_logic;
signal \N__33778\ : std_logic;
signal \N__33775\ : std_logic;
signal \N__33772\ : std_logic;
signal \N__33769\ : std_logic;
signal \N__33766\ : std_logic;
signal \N__33763\ : std_logic;
signal \N__33760\ : std_logic;
signal \N__33757\ : std_logic;
signal \N__33754\ : std_logic;
signal \N__33751\ : std_logic;
signal \N__33748\ : std_logic;
signal \N__33745\ : std_logic;
signal \N__33742\ : std_logic;
signal \N__33739\ : std_logic;
signal \N__33736\ : std_logic;
signal \N__33733\ : std_logic;
signal \N__33730\ : std_logic;
signal \N__33727\ : std_logic;
signal \N__33724\ : std_logic;
signal \N__33721\ : std_logic;
signal \N__33718\ : std_logic;
signal \N__33715\ : std_logic;
signal \N__33712\ : std_logic;
signal \N__33709\ : std_logic;
signal \N__33706\ : std_logic;
signal \N__33703\ : std_logic;
signal \N__33698\ : std_logic;
signal \N__33695\ : std_logic;
signal \N__33692\ : std_logic;
signal \N__33689\ : std_logic;
signal \N__33686\ : std_logic;
signal \N__33683\ : std_logic;
signal \N__33682\ : std_logic;
signal \N__33679\ : std_logic;
signal \N__33676\ : std_logic;
signal \N__33673\ : std_logic;
signal \N__33670\ : std_logic;
signal \N__33669\ : std_logic;
signal \N__33664\ : std_logic;
signal \N__33661\ : std_logic;
signal \N__33658\ : std_logic;
signal \N__33655\ : std_logic;
signal \N__33652\ : std_logic;
signal \N__33649\ : std_logic;
signal \N__33648\ : std_logic;
signal \N__33645\ : std_logic;
signal \N__33642\ : std_logic;
signal \N__33639\ : std_logic;
signal \N__33632\ : std_logic;
signal \N__33629\ : std_logic;
signal \N__33626\ : std_logic;
signal \N__33623\ : std_logic;
signal \N__33620\ : std_logic;
signal \N__33617\ : std_logic;
signal \N__33614\ : std_logic;
signal \N__33611\ : std_logic;
signal \N__33608\ : std_logic;
signal \N__33605\ : std_logic;
signal \N__33602\ : std_logic;
signal \N__33599\ : std_logic;
signal \N__33596\ : std_logic;
signal \N__33593\ : std_logic;
signal \N__33590\ : std_logic;
signal \N__33589\ : std_logic;
signal \N__33586\ : std_logic;
signal \N__33583\ : std_logic;
signal \N__33580\ : std_logic;
signal \N__33577\ : std_logic;
signal \N__33574\ : std_logic;
signal \N__33571\ : std_logic;
signal \N__33568\ : std_logic;
signal \N__33565\ : std_logic;
signal \N__33562\ : std_logic;
signal \N__33559\ : std_logic;
signal \N__33556\ : std_logic;
signal \N__33553\ : std_logic;
signal \N__33550\ : std_logic;
signal \N__33547\ : std_logic;
signal \N__33544\ : std_logic;
signal \N__33541\ : std_logic;
signal \N__33538\ : std_logic;
signal \N__33535\ : std_logic;
signal \N__33532\ : std_logic;
signal \N__33529\ : std_logic;
signal \N__33526\ : std_logic;
signal \N__33523\ : std_logic;
signal \N__33520\ : std_logic;
signal \N__33517\ : std_logic;
signal \N__33512\ : std_logic;
signal \N__33509\ : std_logic;
signal \N__33506\ : std_logic;
signal \N__33503\ : std_logic;
signal \N__33500\ : std_logic;
signal \N__33497\ : std_logic;
signal \N__33494\ : std_logic;
signal \N__33491\ : std_logic;
signal \N__33488\ : std_logic;
signal \N__33485\ : std_logic;
signal \N__33482\ : std_logic;
signal \N__33479\ : std_logic;
signal \N__33476\ : std_logic;
signal \N__33475\ : std_logic;
signal \N__33472\ : std_logic;
signal \N__33469\ : std_logic;
signal \N__33466\ : std_logic;
signal \N__33463\ : std_logic;
signal \N__33460\ : std_logic;
signal \N__33457\ : std_logic;
signal \N__33454\ : std_logic;
signal \N__33451\ : std_logic;
signal \N__33448\ : std_logic;
signal \N__33445\ : std_logic;
signal \N__33442\ : std_logic;
signal \N__33439\ : std_logic;
signal \N__33436\ : std_logic;
signal \N__33433\ : std_logic;
signal \N__33430\ : std_logic;
signal \N__33427\ : std_logic;
signal \N__33424\ : std_logic;
signal \N__33421\ : std_logic;
signal \N__33418\ : std_logic;
signal \N__33415\ : std_logic;
signal \N__33412\ : std_logic;
signal \N__33409\ : std_logic;
signal \N__33406\ : std_logic;
signal \N__33403\ : std_logic;
signal \N__33398\ : std_logic;
signal \N__33397\ : std_logic;
signal \N__33394\ : std_logic;
signal \N__33391\ : std_logic;
signal \N__33388\ : std_logic;
signal \N__33385\ : std_logic;
signal \N__33382\ : std_logic;
signal \N__33381\ : std_logic;
signal \N__33380\ : std_logic;
signal \N__33375\ : std_logic;
signal \N__33372\ : std_logic;
signal \N__33369\ : std_logic;
signal \N__33366\ : std_logic;
signal \N__33361\ : std_logic;
signal \N__33356\ : std_logic;
signal \N__33353\ : std_logic;
signal \N__33350\ : std_logic;
signal \N__33347\ : std_logic;
signal \N__33344\ : std_logic;
signal \N__33341\ : std_logic;
signal \N__33338\ : std_logic;
signal \N__33337\ : std_logic;
signal \N__33336\ : std_logic;
signal \N__33333\ : std_logic;
signal \N__33330\ : std_logic;
signal \N__33329\ : std_logic;
signal \N__33326\ : std_logic;
signal \N__33325\ : std_logic;
signal \N__33322\ : std_logic;
signal \N__33319\ : std_logic;
signal \N__33316\ : std_logic;
signal \N__33313\ : std_logic;
signal \N__33310\ : std_logic;
signal \N__33305\ : std_logic;
signal \N__33302\ : std_logic;
signal \N__33297\ : std_logic;
signal \N__33294\ : std_logic;
signal \N__33291\ : std_logic;
signal \N__33288\ : std_logic;
signal \N__33285\ : std_logic;
signal \N__33280\ : std_logic;
signal \N__33275\ : std_logic;
signal \N__33272\ : std_logic;
signal \N__33269\ : std_logic;
signal \N__33266\ : std_logic;
signal \N__33263\ : std_logic;
signal \N__33260\ : std_logic;
signal \N__33257\ : std_logic;
signal \N__33256\ : std_logic;
signal \N__33255\ : std_logic;
signal \N__33254\ : std_logic;
signal \N__33251\ : std_logic;
signal \N__33248\ : std_logic;
signal \N__33245\ : std_logic;
signal \N__33244\ : std_logic;
signal \N__33241\ : std_logic;
signal \N__33238\ : std_logic;
signal \N__33235\ : std_logic;
signal \N__33232\ : std_logic;
signal \N__33229\ : std_logic;
signal \N__33226\ : std_logic;
signal \N__33223\ : std_logic;
signal \N__33218\ : std_logic;
signal \N__33215\ : std_logic;
signal \N__33212\ : std_logic;
signal \N__33207\ : std_logic;
signal \N__33200\ : std_logic;
signal \N__33197\ : std_logic;
signal \N__33194\ : std_logic;
signal \N__33191\ : std_logic;
signal \N__33188\ : std_logic;
signal \N__33187\ : std_logic;
signal \N__33184\ : std_logic;
signal \N__33181\ : std_logic;
signal \N__33180\ : std_logic;
signal \N__33177\ : std_logic;
signal \N__33174\ : std_logic;
signal \N__33171\ : std_logic;
signal \N__33168\ : std_logic;
signal \N__33167\ : std_logic;
signal \N__33164\ : std_logic;
signal \N__33159\ : std_logic;
signal \N__33156\ : std_logic;
signal \N__33153\ : std_logic;
signal \N__33146\ : std_logic;
signal \N__33143\ : std_logic;
signal \N__33140\ : std_logic;
signal \N__33139\ : std_logic;
signal \N__33136\ : std_logic;
signal \N__33135\ : std_logic;
signal \N__33132\ : std_logic;
signal \N__33131\ : std_logic;
signal \N__33128\ : std_logic;
signal \N__33125\ : std_logic;
signal \N__33124\ : std_logic;
signal \N__33121\ : std_logic;
signal \N__33118\ : std_logic;
signal \N__33115\ : std_logic;
signal \N__33112\ : std_logic;
signal \N__33109\ : std_logic;
signal \N__33106\ : std_logic;
signal \N__33103\ : std_logic;
signal \N__33100\ : std_logic;
signal \N__33097\ : std_logic;
signal \N__33094\ : std_logic;
signal \N__33089\ : std_logic;
signal \N__33084\ : std_logic;
signal \N__33081\ : std_logic;
signal \N__33078\ : std_logic;
signal \N__33071\ : std_logic;
signal \N__33068\ : std_logic;
signal \N__33065\ : std_logic;
signal \N__33062\ : std_logic;
signal \N__33061\ : std_logic;
signal \N__33058\ : std_logic;
signal \N__33055\ : std_logic;
signal \N__33054\ : std_logic;
signal \N__33051\ : std_logic;
signal \N__33050\ : std_logic;
signal \N__33047\ : std_logic;
signal \N__33044\ : std_logic;
signal \N__33041\ : std_logic;
signal \N__33038\ : std_logic;
signal \N__33035\ : std_logic;
signal \N__33030\ : std_logic;
signal \N__33027\ : std_logic;
signal \N__33020\ : std_logic;
signal \N__33019\ : std_logic;
signal \N__33016\ : std_logic;
signal \N__33015\ : std_logic;
signal \N__33014\ : std_logic;
signal \N__33011\ : std_logic;
signal \N__33010\ : std_logic;
signal \N__33007\ : std_logic;
signal \N__33004\ : std_logic;
signal \N__33001\ : std_logic;
signal \N__32998\ : std_logic;
signal \N__32995\ : std_logic;
signal \N__32992\ : std_logic;
signal \N__32989\ : std_logic;
signal \N__32986\ : std_logic;
signal \N__32983\ : std_logic;
signal \N__32980\ : std_logic;
signal \N__32975\ : std_logic;
signal \N__32966\ : std_logic;
signal \N__32965\ : std_logic;
signal \N__32964\ : std_logic;
signal \N__32963\ : std_logic;
signal \N__32960\ : std_logic;
signal \N__32959\ : std_logic;
signal \N__32958\ : std_logic;
signal \N__32955\ : std_logic;
signal \N__32952\ : std_logic;
signal \N__32949\ : std_logic;
signal \N__32946\ : std_logic;
signal \N__32943\ : std_logic;
signal \N__32940\ : std_logic;
signal \N__32937\ : std_logic;
signal \N__32934\ : std_logic;
signal \N__32931\ : std_logic;
signal \N__32930\ : std_logic;
signal \N__32925\ : std_logic;
signal \N__32922\ : std_logic;
signal \N__32919\ : std_logic;
signal \N__32914\ : std_logic;
signal \N__32911\ : std_logic;
signal \N__32900\ : std_logic;
signal \N__32899\ : std_logic;
signal \N__32898\ : std_logic;
signal \N__32897\ : std_logic;
signal \N__32896\ : std_logic;
signal \N__32893\ : std_logic;
signal \N__32890\ : std_logic;
signal \N__32885\ : std_logic;
signal \N__32882\ : std_logic;
signal \N__32873\ : std_logic;
signal \N__32872\ : std_logic;
signal \N__32869\ : std_logic;
signal \N__32866\ : std_logic;
signal \N__32863\ : std_logic;
signal \N__32860\ : std_logic;
signal \N__32859\ : std_logic;
signal \N__32854\ : std_logic;
signal \N__32853\ : std_logic;
signal \N__32850\ : std_logic;
signal \N__32847\ : std_logic;
signal \N__32844\ : std_logic;
signal \N__32841\ : std_logic;
signal \N__32836\ : std_logic;
signal \N__32833\ : std_logic;
signal \N__32830\ : std_logic;
signal \N__32825\ : std_logic;
signal \N__32822\ : std_logic;
signal \N__32819\ : std_logic;
signal \N__32816\ : std_logic;
signal \N__32813\ : std_logic;
signal \N__32810\ : std_logic;
signal \N__32807\ : std_logic;
signal \N__32804\ : std_logic;
signal \N__32801\ : std_logic;
signal \N__32798\ : std_logic;
signal \N__32795\ : std_logic;
signal \N__32792\ : std_logic;
signal \N__32789\ : std_logic;
signal \N__32786\ : std_logic;
signal \N__32785\ : std_logic;
signal \N__32782\ : std_logic;
signal \N__32779\ : std_logic;
signal \N__32776\ : std_logic;
signal \N__32773\ : std_logic;
signal \N__32770\ : std_logic;
signal \N__32767\ : std_logic;
signal \N__32764\ : std_logic;
signal \N__32761\ : std_logic;
signal \N__32758\ : std_logic;
signal \N__32755\ : std_logic;
signal \N__32752\ : std_logic;
signal \N__32749\ : std_logic;
signal \N__32746\ : std_logic;
signal \N__32743\ : std_logic;
signal \N__32740\ : std_logic;
signal \N__32737\ : std_logic;
signal \N__32734\ : std_logic;
signal \N__32731\ : std_logic;
signal \N__32728\ : std_logic;
signal \N__32725\ : std_logic;
signal \N__32722\ : std_logic;
signal \N__32719\ : std_logic;
signal \N__32716\ : std_logic;
signal \N__32713\ : std_logic;
signal \N__32710\ : std_logic;
signal \N__32705\ : std_logic;
signal \N__32702\ : std_logic;
signal \N__32699\ : std_logic;
signal \N__32696\ : std_logic;
signal \N__32693\ : std_logic;
signal \N__32690\ : std_logic;
signal \N__32687\ : std_logic;
signal \N__32684\ : std_logic;
signal \N__32681\ : std_logic;
signal \N__32678\ : std_logic;
signal \N__32675\ : std_logic;
signal \N__32672\ : std_logic;
signal \N__32669\ : std_logic;
signal \N__32666\ : std_logic;
signal \N__32663\ : std_logic;
signal \N__32660\ : std_logic;
signal \N__32657\ : std_logic;
signal \N__32656\ : std_logic;
signal \N__32653\ : std_logic;
signal \N__32652\ : std_logic;
signal \N__32649\ : std_logic;
signal \N__32646\ : std_logic;
signal \N__32643\ : std_logic;
signal \N__32636\ : std_logic;
signal \N__32633\ : std_logic;
signal \N__32630\ : std_logic;
signal \N__32627\ : std_logic;
signal \N__32624\ : std_logic;
signal \N__32623\ : std_logic;
signal \N__32620\ : std_logic;
signal \N__32619\ : std_logic;
signal \N__32616\ : std_logic;
signal \N__32613\ : std_logic;
signal \N__32610\ : std_logic;
signal \N__32603\ : std_logic;
signal \N__32600\ : std_logic;
signal \N__32599\ : std_logic;
signal \N__32596\ : std_logic;
signal \N__32593\ : std_logic;
signal \N__32590\ : std_logic;
signal \N__32587\ : std_logic;
signal \N__32586\ : std_logic;
signal \N__32583\ : std_logic;
signal \N__32580\ : std_logic;
signal \N__32577\ : std_logic;
signal \N__32572\ : std_logic;
signal \N__32567\ : std_logic;
signal \N__32564\ : std_logic;
signal \N__32561\ : std_logic;
signal \N__32558\ : std_logic;
signal \N__32555\ : std_logic;
signal \N__32552\ : std_logic;
signal \N__32549\ : std_logic;
signal \N__32546\ : std_logic;
signal \N__32545\ : std_logic;
signal \N__32544\ : std_logic;
signal \N__32543\ : std_logic;
signal \N__32542\ : std_logic;
signal \N__32541\ : std_logic;
signal \N__32540\ : std_logic;
signal \N__32539\ : std_logic;
signal \N__32538\ : std_logic;
signal \N__32537\ : std_logic;
signal \N__32536\ : std_logic;
signal \N__32535\ : std_logic;
signal \N__32530\ : std_logic;
signal \N__32525\ : std_logic;
signal \N__32522\ : std_logic;
signal \N__32517\ : std_logic;
signal \N__32514\ : std_logic;
signal \N__32511\ : std_logic;
signal \N__32506\ : std_logic;
signal \N__32503\ : std_logic;
signal \N__32500\ : std_logic;
signal \N__32497\ : std_logic;
signal \N__32494\ : std_logic;
signal \N__32485\ : std_logic;
signal \N__32482\ : std_logic;
signal \N__32477\ : std_logic;
signal \N__32474\ : std_logic;
signal \N__32465\ : std_logic;
signal \N__32462\ : std_logic;
signal \N__32459\ : std_logic;
signal \N__32458\ : std_logic;
signal \N__32455\ : std_logic;
signal \N__32452\ : std_logic;
signal \N__32449\ : std_logic;
signal \N__32448\ : std_logic;
signal \N__32445\ : std_logic;
signal \N__32442\ : std_logic;
signal \N__32439\ : std_logic;
signal \N__32438\ : std_logic;
signal \N__32435\ : std_logic;
signal \N__32434\ : std_logic;
signal \N__32429\ : std_logic;
signal \N__32426\ : std_logic;
signal \N__32423\ : std_logic;
signal \N__32420\ : std_logic;
signal \N__32417\ : std_logic;
signal \N__32408\ : std_logic;
signal \N__32407\ : std_logic;
signal \N__32406\ : std_logic;
signal \N__32405\ : std_logic;
signal \N__32402\ : std_logic;
signal \N__32399\ : std_logic;
signal \N__32398\ : std_logic;
signal \N__32397\ : std_logic;
signal \N__32396\ : std_logic;
signal \N__32395\ : std_logic;
signal \N__32394\ : std_logic;
signal \N__32393\ : std_logic;
signal \N__32392\ : std_logic;
signal \N__32391\ : std_logic;
signal \N__32386\ : std_logic;
signal \N__32383\ : std_logic;
signal \N__32380\ : std_logic;
signal \N__32377\ : std_logic;
signal \N__32374\ : std_logic;
signal \N__32369\ : std_logic;
signal \N__32366\ : std_logic;
signal \N__32359\ : std_logic;
signal \N__32350\ : std_logic;
signal \N__32349\ : std_logic;
signal \N__32344\ : std_logic;
signal \N__32341\ : std_logic;
signal \N__32336\ : std_logic;
signal \N__32333\ : std_logic;
signal \N__32324\ : std_logic;
signal \N__32321\ : std_logic;
signal \N__32318\ : std_logic;
signal \N__32315\ : std_logic;
signal \N__32312\ : std_logic;
signal \N__32309\ : std_logic;
signal \N__32306\ : std_logic;
signal \N__32305\ : std_logic;
signal \N__32302\ : std_logic;
signal \N__32301\ : std_logic;
signal \N__32298\ : std_logic;
signal \N__32295\ : std_logic;
signal \N__32292\ : std_logic;
signal \N__32285\ : std_logic;
signal \N__32284\ : std_logic;
signal \N__32283\ : std_logic;
signal \N__32282\ : std_logic;
signal \N__32279\ : std_logic;
signal \N__32276\ : std_logic;
signal \N__32273\ : std_logic;
signal \N__32270\ : std_logic;
signal \N__32267\ : std_logic;
signal \N__32264\ : std_logic;
signal \N__32261\ : std_logic;
signal \N__32258\ : std_logic;
signal \N__32255\ : std_logic;
signal \N__32252\ : std_logic;
signal \N__32249\ : std_logic;
signal \N__32246\ : std_logic;
signal \N__32241\ : std_logic;
signal \N__32236\ : std_logic;
signal \N__32231\ : std_logic;
signal \N__32230\ : std_logic;
signal \N__32229\ : std_logic;
signal \N__32226\ : std_logic;
signal \N__32223\ : std_logic;
signal \N__32220\ : std_logic;
signal \N__32215\ : std_logic;
signal \N__32210\ : std_logic;
signal \N__32209\ : std_logic;
signal \N__32206\ : std_logic;
signal \N__32205\ : std_logic;
signal \N__32204\ : std_logic;
signal \N__32201\ : std_logic;
signal \N__32198\ : std_logic;
signal \N__32195\ : std_logic;
signal \N__32192\ : std_logic;
signal \N__32189\ : std_logic;
signal \N__32186\ : std_logic;
signal \N__32183\ : std_logic;
signal \N__32180\ : std_logic;
signal \N__32177\ : std_logic;
signal \N__32172\ : std_logic;
signal \N__32169\ : std_logic;
signal \N__32166\ : std_logic;
signal \N__32163\ : std_logic;
signal \N__32160\ : std_logic;
signal \N__32153\ : std_logic;
signal \N__32152\ : std_logic;
signal \N__32151\ : std_logic;
signal \N__32148\ : std_logic;
signal \N__32145\ : std_logic;
signal \N__32142\ : std_logic;
signal \N__32139\ : std_logic;
signal \N__32132\ : std_logic;
signal \N__32131\ : std_logic;
signal \N__32128\ : std_logic;
signal \N__32125\ : std_logic;
signal \N__32124\ : std_logic;
signal \N__32121\ : std_logic;
signal \N__32118\ : std_logic;
signal \N__32117\ : std_logic;
signal \N__32114\ : std_logic;
signal \N__32111\ : std_logic;
signal \N__32108\ : std_logic;
signal \N__32105\ : std_logic;
signal \N__32102\ : std_logic;
signal \N__32099\ : std_logic;
signal \N__32096\ : std_logic;
signal \N__32093\ : std_logic;
signal \N__32084\ : std_logic;
signal \N__32083\ : std_logic;
signal \N__32082\ : std_logic;
signal \N__32079\ : std_logic;
signal \N__32076\ : std_logic;
signal \N__32073\ : std_logic;
signal \N__32070\ : std_logic;
signal \N__32065\ : std_logic;
signal \N__32060\ : std_logic;
signal \N__32059\ : std_logic;
signal \N__32056\ : std_logic;
signal \N__32053\ : std_logic;
signal \N__32052\ : std_logic;
signal \N__32051\ : std_logic;
signal \N__32048\ : std_logic;
signal \N__32045\ : std_logic;
signal \N__32042\ : std_logic;
signal \N__32039\ : std_logic;
signal \N__32036\ : std_logic;
signal \N__32033\ : std_logic;
signal \N__32030\ : std_logic;
signal \N__32027\ : std_logic;
signal \N__32026\ : std_logic;
signal \N__32025\ : std_logic;
signal \N__32024\ : std_logic;
signal \N__32021\ : std_logic;
signal \N__32016\ : std_logic;
signal \N__32013\ : std_logic;
signal \N__32008\ : std_logic;
signal \N__32005\ : std_logic;
signal \N__31994\ : std_logic;
signal \N__31993\ : std_logic;
signal \N__31990\ : std_logic;
signal \N__31989\ : std_logic;
signal \N__31986\ : std_logic;
signal \N__31985\ : std_logic;
signal \N__31982\ : std_logic;
signal \N__31979\ : std_logic;
signal \N__31976\ : std_logic;
signal \N__31973\ : std_logic;
signal \N__31966\ : std_logic;
signal \N__31963\ : std_logic;
signal \N__31958\ : std_logic;
signal \N__31955\ : std_logic;
signal \N__31954\ : std_logic;
signal \N__31951\ : std_logic;
signal \N__31950\ : std_logic;
signal \N__31947\ : std_logic;
signal \N__31946\ : std_logic;
signal \N__31943\ : std_logic;
signal \N__31940\ : std_logic;
signal \N__31937\ : std_logic;
signal \N__31934\ : std_logic;
signal \N__31931\ : std_logic;
signal \N__31928\ : std_logic;
signal \N__31919\ : std_logic;
signal \N__31918\ : std_logic;
signal \N__31917\ : std_logic;
signal \N__31914\ : std_logic;
signal \N__31909\ : std_logic;
signal \N__31908\ : std_logic;
signal \N__31907\ : std_logic;
signal \N__31906\ : std_logic;
signal \N__31905\ : std_logic;
signal \N__31904\ : std_logic;
signal \N__31903\ : std_logic;
signal \N__31902\ : std_logic;
signal \N__31901\ : std_logic;
signal \N__31900\ : std_logic;
signal \N__31899\ : std_logic;
signal \N__31898\ : std_logic;
signal \N__31897\ : std_logic;
signal \N__31896\ : std_logic;
signal \N__31895\ : std_logic;
signal \N__31894\ : std_logic;
signal \N__31889\ : std_logic;
signal \N__31876\ : std_logic;
signal \N__31873\ : std_logic;
signal \N__31864\ : std_logic;
signal \N__31859\ : std_logic;
signal \N__31858\ : std_logic;
signal \N__31853\ : std_logic;
signal \N__31848\ : std_logic;
signal \N__31843\ : std_logic;
signal \N__31840\ : std_logic;
signal \N__31837\ : std_logic;
signal \N__31834\ : std_logic;
signal \N__31833\ : std_logic;
signal \N__31832\ : std_logic;
signal \N__31831\ : std_logic;
signal \N__31828\ : std_logic;
signal \N__31825\ : std_logic;
signal \N__31820\ : std_logic;
signal \N__31817\ : std_logic;
signal \N__31814\ : std_logic;
signal \N__31809\ : std_logic;
signal \N__31802\ : std_logic;
signal \N__31795\ : std_logic;
signal \N__31792\ : std_logic;
signal \N__31789\ : std_logic;
signal \N__31786\ : std_logic;
signal \N__31781\ : std_logic;
signal \N__31780\ : std_logic;
signal \N__31777\ : std_logic;
signal \N__31776\ : std_logic;
signal \N__31773\ : std_logic;
signal \N__31772\ : std_logic;
signal \N__31769\ : std_logic;
signal \N__31766\ : std_logic;
signal \N__31763\ : std_logic;
signal \N__31760\ : std_logic;
signal \N__31757\ : std_logic;
signal \N__31754\ : std_logic;
signal \N__31751\ : std_logic;
signal \N__31748\ : std_logic;
signal \N__31745\ : std_logic;
signal \N__31742\ : std_logic;
signal \N__31737\ : std_logic;
signal \N__31730\ : std_logic;
signal \N__31727\ : std_logic;
signal \N__31726\ : std_logic;
signal \N__31723\ : std_logic;
signal \N__31720\ : std_logic;
signal \N__31719\ : std_logic;
signal \N__31718\ : std_logic;
signal \N__31715\ : std_logic;
signal \N__31712\ : std_logic;
signal \N__31709\ : std_logic;
signal \N__31706\ : std_logic;
signal \N__31703\ : std_logic;
signal \N__31700\ : std_logic;
signal \N__31697\ : std_logic;
signal \N__31688\ : std_logic;
signal \N__31687\ : std_logic;
signal \N__31686\ : std_logic;
signal \N__31683\ : std_logic;
signal \N__31680\ : std_logic;
signal \N__31677\ : std_logic;
signal \N__31674\ : std_logic;
signal \N__31673\ : std_logic;
signal \N__31672\ : std_logic;
signal \N__31671\ : std_logic;
signal \N__31668\ : std_logic;
signal \N__31667\ : std_logic;
signal \N__31666\ : std_logic;
signal \N__31663\ : std_logic;
signal \N__31660\ : std_logic;
signal \N__31657\ : std_logic;
signal \N__31654\ : std_logic;
signal \N__31651\ : std_logic;
signal \N__31648\ : std_logic;
signal \N__31645\ : std_logic;
signal \N__31642\ : std_logic;
signal \N__31639\ : std_logic;
signal \N__31634\ : std_logic;
signal \N__31631\ : std_logic;
signal \N__31626\ : std_logic;
signal \N__31623\ : std_logic;
signal \N__31622\ : std_logic;
signal \N__31619\ : std_logic;
signal \N__31614\ : std_logic;
signal \N__31613\ : std_logic;
signal \N__31610\ : std_logic;
signal \N__31605\ : std_logic;
signal \N__31604\ : std_logic;
signal \N__31601\ : std_logic;
signal \N__31598\ : std_logic;
signal \N__31595\ : std_logic;
signal \N__31592\ : std_logic;
signal \N__31587\ : std_logic;
signal \N__31584\ : std_logic;
signal \N__31571\ : std_logic;
signal \N__31570\ : std_logic;
signal \N__31567\ : std_logic;
signal \N__31564\ : std_logic;
signal \N__31563\ : std_logic;
signal \N__31562\ : std_logic;
signal \N__31559\ : std_logic;
signal \N__31556\ : std_logic;
signal \N__31553\ : std_logic;
signal \N__31550\ : std_logic;
signal \N__31543\ : std_logic;
signal \N__31540\ : std_logic;
signal \N__31537\ : std_logic;
signal \N__31534\ : std_logic;
signal \N__31529\ : std_logic;
signal \N__31526\ : std_logic;
signal \N__31525\ : std_logic;
signal \N__31522\ : std_logic;
signal \N__31519\ : std_logic;
signal \N__31518\ : std_logic;
signal \N__31515\ : std_logic;
signal \N__31514\ : std_logic;
signal \N__31511\ : std_logic;
signal \N__31508\ : std_logic;
signal \N__31505\ : std_logic;
signal \N__31502\ : std_logic;
signal \N__31499\ : std_logic;
signal \N__31490\ : std_logic;
signal \N__31489\ : std_logic;
signal \N__31488\ : std_logic;
signal \N__31487\ : std_logic;
signal \N__31484\ : std_logic;
signal \N__31483\ : std_logic;
signal \N__31480\ : std_logic;
signal \N__31477\ : std_logic;
signal \N__31474\ : std_logic;
signal \N__31471\ : std_logic;
signal \N__31468\ : std_logic;
signal \N__31465\ : std_logic;
signal \N__31462\ : std_logic;
signal \N__31459\ : std_logic;
signal \N__31450\ : std_logic;
signal \N__31445\ : std_logic;
signal \N__31442\ : std_logic;
signal \N__31439\ : std_logic;
signal \N__31438\ : std_logic;
signal \N__31435\ : std_logic;
signal \N__31432\ : std_logic;
signal \N__31427\ : std_logic;
signal \N__31426\ : std_logic;
signal \N__31423\ : std_logic;
signal \N__31420\ : std_logic;
signal \N__31415\ : std_logic;
signal \N__31412\ : std_logic;
signal \N__31409\ : std_logic;
signal \N__31406\ : std_logic;
signal \N__31403\ : std_logic;
signal \N__31400\ : std_logic;
signal \N__31397\ : std_logic;
signal \N__31396\ : std_logic;
signal \N__31395\ : std_logic;
signal \N__31394\ : std_logic;
signal \N__31391\ : std_logic;
signal \N__31388\ : std_logic;
signal \N__31385\ : std_logic;
signal \N__31382\ : std_logic;
signal \N__31377\ : std_logic;
signal \N__31374\ : std_logic;
signal \N__31371\ : std_logic;
signal \N__31368\ : std_logic;
signal \N__31363\ : std_logic;
signal \N__31360\ : std_logic;
signal \N__31357\ : std_logic;
signal \N__31352\ : std_logic;
signal \N__31351\ : std_logic;
signal \N__31350\ : std_logic;
signal \N__31347\ : std_logic;
signal \N__31346\ : std_logic;
signal \N__31343\ : std_logic;
signal \N__31340\ : std_logic;
signal \N__31337\ : std_logic;
signal \N__31334\ : std_logic;
signal \N__31331\ : std_logic;
signal \N__31330\ : std_logic;
signal \N__31327\ : std_logic;
signal \N__31322\ : std_logic;
signal \N__31319\ : std_logic;
signal \N__31316\ : std_logic;
signal \N__31311\ : std_logic;
signal \N__31304\ : std_logic;
signal \N__31301\ : std_logic;
signal \N__31300\ : std_logic;
signal \N__31299\ : std_logic;
signal \N__31296\ : std_logic;
signal \N__31293\ : std_logic;
signal \N__31290\ : std_logic;
signal \N__31287\ : std_logic;
signal \N__31284\ : std_logic;
signal \N__31283\ : std_logic;
signal \N__31282\ : std_logic;
signal \N__31279\ : std_logic;
signal \N__31276\ : std_logic;
signal \N__31273\ : std_logic;
signal \N__31268\ : std_logic;
signal \N__31265\ : std_logic;
signal \N__31256\ : std_logic;
signal \N__31255\ : std_logic;
signal \N__31252\ : std_logic;
signal \N__31249\ : std_logic;
signal \N__31246\ : std_logic;
signal \N__31245\ : std_logic;
signal \N__31242\ : std_logic;
signal \N__31241\ : std_logic;
signal \N__31238\ : std_logic;
signal \N__31235\ : std_logic;
signal \N__31232\ : std_logic;
signal \N__31229\ : std_logic;
signal \N__31224\ : std_logic;
signal \N__31223\ : std_logic;
signal \N__31220\ : std_logic;
signal \N__31217\ : std_logic;
signal \N__31214\ : std_logic;
signal \N__31211\ : std_logic;
signal \N__31202\ : std_logic;
signal \N__31199\ : std_logic;
signal \N__31196\ : std_logic;
signal \N__31195\ : std_logic;
signal \N__31192\ : std_logic;
signal \N__31189\ : std_logic;
signal \N__31184\ : std_logic;
signal \N__31181\ : std_logic;
signal \N__31180\ : std_logic;
signal \N__31179\ : std_logic;
signal \N__31178\ : std_logic;
signal \N__31177\ : std_logic;
signal \N__31176\ : std_logic;
signal \N__31175\ : std_logic;
signal \N__31174\ : std_logic;
signal \N__31173\ : std_logic;
signal \N__31172\ : std_logic;
signal \N__31171\ : std_logic;
signal \N__31170\ : std_logic;
signal \N__31169\ : std_logic;
signal \N__31168\ : std_logic;
signal \N__31167\ : std_logic;
signal \N__31166\ : std_logic;
signal \N__31165\ : std_logic;
signal \N__31164\ : std_logic;
signal \N__31161\ : std_logic;
signal \N__31158\ : std_logic;
signal \N__31151\ : std_logic;
signal \N__31148\ : std_logic;
signal \N__31139\ : std_logic;
signal \N__31130\ : std_logic;
signal \N__31129\ : std_logic;
signal \N__31120\ : std_logic;
signal \N__31119\ : std_logic;
signal \N__31118\ : std_logic;
signal \N__31117\ : std_logic;
signal \N__31116\ : std_logic;
signal \N__31115\ : std_logic;
signal \N__31114\ : std_logic;
signal \N__31113\ : std_logic;
signal \N__31112\ : std_logic;
signal \N__31111\ : std_logic;
signal \N__31110\ : std_logic;
signal \N__31105\ : std_logic;
signal \N__31096\ : std_logic;
signal \N__31093\ : std_logic;
signal \N__31090\ : std_logic;
signal \N__31077\ : std_logic;
signal \N__31068\ : std_logic;
signal \N__31061\ : std_logic;
signal \N__31056\ : std_logic;
signal \N__31049\ : std_logic;
signal \N__31046\ : std_logic;
signal \N__31043\ : std_logic;
signal \N__31042\ : std_logic;
signal \N__31041\ : std_logic;
signal \N__31038\ : std_logic;
signal \N__31037\ : std_logic;
signal \N__31034\ : std_logic;
signal \N__31031\ : std_logic;
signal \N__31028\ : std_logic;
signal \N__31025\ : std_logic;
signal \N__31022\ : std_logic;
signal \N__31019\ : std_logic;
signal \N__31014\ : std_logic;
signal \N__31011\ : std_logic;
signal \N__31010\ : std_logic;
signal \N__31007\ : std_logic;
signal \N__31002\ : std_logic;
signal \N__30999\ : std_logic;
signal \N__30992\ : std_logic;
signal \N__30991\ : std_logic;
signal \N__30990\ : std_logic;
signal \N__30989\ : std_logic;
signal \N__30988\ : std_logic;
signal \N__30987\ : std_logic;
signal \N__30984\ : std_logic;
signal \N__30983\ : std_logic;
signal \N__30982\ : std_logic;
signal \N__30981\ : std_logic;
signal \N__30980\ : std_logic;
signal \N__30979\ : std_logic;
signal \N__30978\ : std_logic;
signal \N__30977\ : std_logic;
signal \N__30972\ : std_logic;
signal \N__30971\ : std_logic;
signal \N__30968\ : std_logic;
signal \N__30965\ : std_logic;
signal \N__30962\ : std_logic;
signal \N__30961\ : std_logic;
signal \N__30958\ : std_logic;
signal \N__30957\ : std_logic;
signal \N__30956\ : std_logic;
signal \N__30953\ : std_logic;
signal \N__30950\ : std_logic;
signal \N__30947\ : std_logic;
signal \N__30946\ : std_logic;
signal \N__30945\ : std_logic;
signal \N__30942\ : std_logic;
signal \N__30941\ : std_logic;
signal \N__30938\ : std_logic;
signal \N__30935\ : std_logic;
signal \N__30932\ : std_logic;
signal \N__30931\ : std_logic;
signal \N__30928\ : std_logic;
signal \N__30925\ : std_logic;
signal \N__30922\ : std_logic;
signal \N__30915\ : std_logic;
signal \N__30912\ : std_logic;
signal \N__30911\ : std_logic;
signal \N__30910\ : std_logic;
signal \N__30907\ : std_logic;
signal \N__30904\ : std_logic;
signal \N__30901\ : std_logic;
signal \N__30894\ : std_logic;
signal \N__30889\ : std_logic;
signal \N__30882\ : std_logic;
signal \N__30879\ : std_logic;
signal \N__30876\ : std_logic;
signal \N__30875\ : std_logic;
signal \N__30874\ : std_logic;
signal \N__30869\ : std_logic;
signal \N__30862\ : std_logic;
signal \N__30861\ : std_logic;
signal \N__30860\ : std_logic;
signal \N__30857\ : std_logic;
signal \N__30854\ : std_logic;
signal \N__30849\ : std_logic;
signal \N__30846\ : std_logic;
signal \N__30843\ : std_logic;
signal \N__30840\ : std_logic;
signal \N__30837\ : std_logic;
signal \N__30834\ : std_logic;
signal \N__30831\ : std_logic;
signal \N__30828\ : std_logic;
signal \N__30825\ : std_logic;
signal \N__30820\ : std_logic;
signal \N__30811\ : std_logic;
signal \N__30806\ : std_logic;
signal \N__30799\ : std_logic;
signal \N__30792\ : std_logic;
signal \N__30787\ : std_logic;
signal \N__30780\ : std_logic;
signal \N__30777\ : std_logic;
signal \N__30770\ : std_logic;
signal \N__30769\ : std_logic;
signal \N__30768\ : std_logic;
signal \N__30765\ : std_logic;
signal \N__30762\ : std_logic;
signal \N__30761\ : std_logic;
signal \N__30758\ : std_logic;
signal \N__30755\ : std_logic;
signal \N__30752\ : std_logic;
signal \N__30749\ : std_logic;
signal \N__30746\ : std_logic;
signal \N__30743\ : std_logic;
signal \N__30738\ : std_logic;
signal \N__30733\ : std_logic;
signal \N__30728\ : std_logic;
signal \N__30725\ : std_logic;
signal \N__30724\ : std_logic;
signal \N__30723\ : std_logic;
signal \N__30720\ : std_logic;
signal \N__30717\ : std_logic;
signal \N__30714\ : std_logic;
signal \N__30709\ : std_logic;
signal \N__30704\ : std_logic;
signal \N__30701\ : std_logic;
signal \N__30698\ : std_logic;
signal \N__30695\ : std_logic;
signal \N__30692\ : std_logic;
signal \N__30691\ : std_logic;
signal \N__30690\ : std_logic;
signal \N__30687\ : std_logic;
signal \N__30684\ : std_logic;
signal \N__30681\ : std_logic;
signal \N__30674\ : std_logic;
signal \N__30671\ : std_logic;
signal \N__30670\ : std_logic;
signal \N__30669\ : std_logic;
signal \N__30664\ : std_logic;
signal \N__30661\ : std_logic;
signal \N__30658\ : std_logic;
signal \N__30657\ : std_logic;
signal \N__30654\ : std_logic;
signal \N__30651\ : std_logic;
signal \N__30648\ : std_logic;
signal \N__30645\ : std_logic;
signal \N__30638\ : std_logic;
signal \N__30635\ : std_logic;
signal \N__30632\ : std_logic;
signal \N__30629\ : std_logic;
signal \N__30628\ : std_logic;
signal \N__30627\ : std_logic;
signal \N__30626\ : std_logic;
signal \N__30625\ : std_logic;
signal \N__30624\ : std_logic;
signal \N__30623\ : std_logic;
signal \N__30622\ : std_logic;
signal \N__30615\ : std_logic;
signal \N__30614\ : std_logic;
signal \N__30613\ : std_logic;
signal \N__30612\ : std_logic;
signal \N__30611\ : std_logic;
signal \N__30610\ : std_logic;
signal \N__30609\ : std_logic;
signal \N__30608\ : std_logic;
signal \N__30607\ : std_logic;
signal \N__30606\ : std_logic;
signal \N__30601\ : std_logic;
signal \N__30594\ : std_logic;
signal \N__30591\ : std_logic;
signal \N__30584\ : std_logic;
signal \N__30577\ : std_logic;
signal \N__30570\ : std_logic;
signal \N__30557\ : std_logic;
signal \N__30556\ : std_logic;
signal \N__30555\ : std_logic;
signal \N__30554\ : std_logic;
signal \N__30553\ : std_logic;
signal \N__30552\ : std_logic;
signal \N__30549\ : std_logic;
signal \N__30546\ : std_logic;
signal \N__30543\ : std_logic;
signal \N__30540\ : std_logic;
signal \N__30537\ : std_logic;
signal \N__30534\ : std_logic;
signal \N__30531\ : std_logic;
signal \N__30528\ : std_logic;
signal \N__30525\ : std_logic;
signal \N__30522\ : std_logic;
signal \N__30517\ : std_logic;
signal \N__30512\ : std_logic;
signal \N__30503\ : std_logic;
signal \N__30500\ : std_logic;
signal \N__30497\ : std_logic;
signal \N__30494\ : std_logic;
signal \N__30493\ : std_logic;
signal \N__30492\ : std_logic;
signal \N__30491\ : std_logic;
signal \N__30488\ : std_logic;
signal \N__30485\ : std_logic;
signal \N__30480\ : std_logic;
signal \N__30473\ : std_logic;
signal \N__30472\ : std_logic;
signal \N__30471\ : std_logic;
signal \N__30468\ : std_logic;
signal \N__30467\ : std_logic;
signal \N__30466\ : std_logic;
signal \N__30463\ : std_logic;
signal \N__30460\ : std_logic;
signal \N__30457\ : std_logic;
signal \N__30452\ : std_logic;
signal \N__30449\ : std_logic;
signal \N__30446\ : std_logic;
signal \N__30443\ : std_logic;
signal \N__30434\ : std_logic;
signal \N__30433\ : std_logic;
signal \N__30430\ : std_logic;
signal \N__30427\ : std_logic;
signal \N__30426\ : std_logic;
signal \N__30423\ : std_logic;
signal \N__30422\ : std_logic;
signal \N__30421\ : std_logic;
signal \N__30420\ : std_logic;
signal \N__30419\ : std_logic;
signal \N__30418\ : std_logic;
signal \N__30417\ : std_logic;
signal \N__30416\ : std_logic;
signal \N__30413\ : std_logic;
signal \N__30412\ : std_logic;
signal \N__30411\ : std_logic;
signal \N__30408\ : std_logic;
signal \N__30405\ : std_logic;
signal \N__30402\ : std_logic;
signal \N__30397\ : std_logic;
signal \N__30390\ : std_logic;
signal \N__30387\ : std_logic;
signal \N__30384\ : std_logic;
signal \N__30383\ : std_logic;
signal \N__30380\ : std_logic;
signal \N__30379\ : std_logic;
signal \N__30378\ : std_logic;
signal \N__30377\ : std_logic;
signal \N__30376\ : std_logic;
signal \N__30375\ : std_logic;
signal \N__30372\ : std_logic;
signal \N__30371\ : std_logic;
signal \N__30368\ : std_logic;
signal \N__30361\ : std_logic;
signal \N__30358\ : std_logic;
signal \N__30355\ : std_logic;
signal \N__30352\ : std_logic;
signal \N__30343\ : std_logic;
signal \N__30338\ : std_logic;
signal \N__30335\ : std_logic;
signal \N__30330\ : std_logic;
signal \N__30321\ : std_logic;
signal \N__30308\ : std_logic;
signal \N__30305\ : std_logic;
signal \N__30304\ : std_logic;
signal \N__30303\ : std_logic;
signal \N__30302\ : std_logic;
signal \N__30299\ : std_logic;
signal \N__30294\ : std_logic;
signal \N__30291\ : std_logic;
signal \N__30286\ : std_logic;
signal \N__30281\ : std_logic;
signal \N__30278\ : std_logic;
signal \N__30277\ : std_logic;
signal \N__30274\ : std_logic;
signal \N__30271\ : std_logic;
signal \N__30268\ : std_logic;
signal \N__30265\ : std_logic;
signal \N__30260\ : std_logic;
signal \N__30257\ : std_logic;
signal \N__30254\ : std_logic;
signal \N__30251\ : std_logic;
signal \N__30248\ : std_logic;
signal \N__30245\ : std_logic;
signal \N__30244\ : std_logic;
signal \N__30243\ : std_logic;
signal \N__30240\ : std_logic;
signal \N__30237\ : std_logic;
signal \N__30234\ : std_logic;
signal \N__30233\ : std_logic;
signal \N__30232\ : std_logic;
signal \N__30227\ : std_logic;
signal \N__30224\ : std_logic;
signal \N__30221\ : std_logic;
signal \N__30218\ : std_logic;
signal \N__30217\ : std_logic;
signal \N__30214\ : std_logic;
signal \N__30211\ : std_logic;
signal \N__30208\ : std_logic;
signal \N__30205\ : std_logic;
signal \N__30202\ : std_logic;
signal \N__30191\ : std_logic;
signal \N__30188\ : std_logic;
signal \N__30185\ : std_logic;
signal \N__30182\ : std_logic;
signal \N__30179\ : std_logic;
signal \N__30176\ : std_logic;
signal \N__30175\ : std_logic;
signal \N__30172\ : std_logic;
signal \N__30171\ : std_logic;
signal \N__30168\ : std_logic;
signal \N__30165\ : std_logic;
signal \N__30162\ : std_logic;
signal \N__30159\ : std_logic;
signal \N__30158\ : std_logic;
signal \N__30153\ : std_logic;
signal \N__30150\ : std_logic;
signal \N__30147\ : std_logic;
signal \N__30144\ : std_logic;
signal \N__30137\ : std_logic;
signal \N__30136\ : std_logic;
signal \N__30133\ : std_logic;
signal \N__30132\ : std_logic;
signal \N__30129\ : std_logic;
signal \N__30126\ : std_logic;
signal \N__30123\ : std_logic;
signal \N__30120\ : std_logic;
signal \N__30115\ : std_logic;
signal \N__30110\ : std_logic;
signal \N__30109\ : std_logic;
signal \N__30106\ : std_logic;
signal \N__30103\ : std_logic;
signal \N__30100\ : std_logic;
signal \N__30095\ : std_logic;
signal \N__30092\ : std_logic;
signal \N__30089\ : std_logic;
signal \N__30086\ : std_logic;
signal \N__30083\ : std_logic;
signal \N__30080\ : std_logic;
signal \N__30077\ : std_logic;
signal \N__30074\ : std_logic;
signal \N__30071\ : std_logic;
signal \N__30068\ : std_logic;
signal \N__30065\ : std_logic;
signal \N__30062\ : std_logic;
signal \N__30059\ : std_logic;
signal \N__30056\ : std_logic;
signal \N__30053\ : std_logic;
signal \N__30050\ : std_logic;
signal \N__30047\ : std_logic;
signal \N__30044\ : std_logic;
signal \N__30041\ : std_logic;
signal \N__30038\ : std_logic;
signal \N__30035\ : std_logic;
signal \N__30034\ : std_logic;
signal \N__30031\ : std_logic;
signal \N__30028\ : std_logic;
signal \N__30025\ : std_logic;
signal \N__30020\ : std_logic;
signal \N__30017\ : std_logic;
signal \N__30014\ : std_logic;
signal \N__30011\ : std_logic;
signal \N__30008\ : std_logic;
signal \N__30005\ : std_logic;
signal \N__30004\ : std_logic;
signal \N__30003\ : std_logic;
signal \N__30000\ : std_logic;
signal \N__29997\ : std_logic;
signal \N__29994\ : std_logic;
signal \N__29989\ : std_logic;
signal \N__29988\ : std_logic;
signal \N__29987\ : std_logic;
signal \N__29984\ : std_logic;
signal \N__29981\ : std_logic;
signal \N__29978\ : std_logic;
signal \N__29975\ : std_logic;
signal \N__29966\ : std_logic;
signal \N__29965\ : std_logic;
signal \N__29964\ : std_logic;
signal \N__29961\ : std_logic;
signal \N__29956\ : std_logic;
signal \N__29953\ : std_logic;
signal \N__29950\ : std_logic;
signal \N__29949\ : std_logic;
signal \N__29948\ : std_logic;
signal \N__29945\ : std_logic;
signal \N__29942\ : std_logic;
signal \N__29939\ : std_logic;
signal \N__29936\ : std_logic;
signal \N__29927\ : std_logic;
signal \N__29926\ : std_logic;
signal \N__29925\ : std_logic;
signal \N__29922\ : std_logic;
signal \N__29919\ : std_logic;
signal \N__29916\ : std_logic;
signal \N__29913\ : std_logic;
signal \N__29910\ : std_logic;
signal \N__29909\ : std_logic;
signal \N__29906\ : std_logic;
signal \N__29903\ : std_logic;
signal \N__29900\ : std_logic;
signal \N__29899\ : std_logic;
signal \N__29896\ : std_logic;
signal \N__29891\ : std_logic;
signal \N__29888\ : std_logic;
signal \N__29885\ : std_logic;
signal \N__29882\ : std_logic;
signal \N__29873\ : std_logic;
signal \N__29870\ : std_logic;
signal \N__29867\ : std_logic;
signal \N__29864\ : std_logic;
signal \N__29863\ : std_logic;
signal \N__29860\ : std_logic;
signal \N__29857\ : std_logic;
signal \N__29852\ : std_logic;
signal \N__29849\ : std_logic;
signal \N__29846\ : std_logic;
signal \N__29843\ : std_logic;
signal \N__29840\ : std_logic;
signal \N__29839\ : std_logic;
signal \N__29838\ : std_logic;
signal \N__29837\ : std_logic;
signal \N__29834\ : std_logic;
signal \N__29831\ : std_logic;
signal \N__29828\ : std_logic;
signal \N__29825\ : std_logic;
signal \N__29822\ : std_logic;
signal \N__29819\ : std_logic;
signal \N__29814\ : std_logic;
signal \N__29811\ : std_logic;
signal \N__29806\ : std_logic;
signal \N__29801\ : std_logic;
signal \N__29798\ : std_logic;
signal \N__29795\ : std_logic;
signal \N__29792\ : std_logic;
signal \N__29789\ : std_logic;
signal \N__29786\ : std_logic;
signal \N__29783\ : std_logic;
signal \N__29780\ : std_logic;
signal \N__29777\ : std_logic;
signal \N__29774\ : std_logic;
signal \N__29771\ : std_logic;
signal \N__29768\ : std_logic;
signal \N__29765\ : std_logic;
signal \N__29762\ : std_logic;
signal \N__29759\ : std_logic;
signal \N__29756\ : std_logic;
signal \N__29753\ : std_logic;
signal \N__29750\ : std_logic;
signal \N__29747\ : std_logic;
signal \N__29744\ : std_logic;
signal \N__29741\ : std_logic;
signal \N__29738\ : std_logic;
signal \N__29737\ : std_logic;
signal \N__29736\ : std_logic;
signal \N__29733\ : std_logic;
signal \N__29730\ : std_logic;
signal \N__29727\ : std_logic;
signal \N__29726\ : std_logic;
signal \N__29725\ : std_logic;
signal \N__29718\ : std_logic;
signal \N__29715\ : std_logic;
signal \N__29712\ : std_logic;
signal \N__29709\ : std_logic;
signal \N__29702\ : std_logic;
signal \N__29701\ : std_logic;
signal \N__29698\ : std_logic;
signal \N__29695\ : std_logic;
signal \N__29692\ : std_logic;
signal \N__29691\ : std_logic;
signal \N__29688\ : std_logic;
signal \N__29685\ : std_logic;
signal \N__29682\ : std_logic;
signal \N__29675\ : std_logic;
signal \N__29674\ : std_logic;
signal \N__29671\ : std_logic;
signal \N__29668\ : std_logic;
signal \N__29665\ : std_logic;
signal \N__29664\ : std_logic;
signal \N__29661\ : std_logic;
signal \N__29658\ : std_logic;
signal \N__29655\ : std_logic;
signal \N__29648\ : std_logic;
signal \N__29645\ : std_logic;
signal \N__29642\ : std_logic;
signal \N__29639\ : std_logic;
signal \N__29636\ : std_logic;
signal \N__29635\ : std_logic;
signal \N__29634\ : std_logic;
signal \N__29633\ : std_logic;
signal \N__29630\ : std_logic;
signal \N__29627\ : std_logic;
signal \N__29622\ : std_logic;
signal \N__29619\ : std_logic;
signal \N__29616\ : std_logic;
signal \N__29615\ : std_logic;
signal \N__29612\ : std_logic;
signal \N__29609\ : std_logic;
signal \N__29606\ : std_logic;
signal \N__29603\ : std_logic;
signal \N__29600\ : std_logic;
signal \N__29591\ : std_logic;
signal \N__29590\ : std_logic;
signal \N__29589\ : std_logic;
signal \N__29586\ : std_logic;
signal \N__29583\ : std_logic;
signal \N__29580\ : std_logic;
signal \N__29577\ : std_logic;
signal \N__29574\ : std_logic;
signal \N__29571\ : std_logic;
signal \N__29566\ : std_logic;
signal \N__29561\ : std_logic;
signal \N__29560\ : std_logic;
signal \N__29559\ : std_logic;
signal \N__29556\ : std_logic;
signal \N__29553\ : std_logic;
signal \N__29552\ : std_logic;
signal \N__29551\ : std_logic;
signal \N__29548\ : std_logic;
signal \N__29545\ : std_logic;
signal \N__29542\ : std_logic;
signal \N__29539\ : std_logic;
signal \N__29536\ : std_logic;
signal \N__29533\ : std_logic;
signal \N__29530\ : std_logic;
signal \N__29525\ : std_logic;
signal \N__29522\ : std_logic;
signal \N__29513\ : std_logic;
signal \N__29512\ : std_logic;
signal \N__29509\ : std_logic;
signal \N__29506\ : std_logic;
signal \N__29505\ : std_logic;
signal \N__29502\ : std_logic;
signal \N__29499\ : std_logic;
signal \N__29496\ : std_logic;
signal \N__29493\ : std_logic;
signal \N__29486\ : std_logic;
signal \N__29485\ : std_logic;
signal \N__29484\ : std_logic;
signal \N__29481\ : std_logic;
signal \N__29478\ : std_logic;
signal \N__29475\ : std_logic;
signal \N__29474\ : std_logic;
signal \N__29469\ : std_logic;
signal \N__29466\ : std_logic;
signal \N__29465\ : std_logic;
signal \N__29462\ : std_logic;
signal \N__29457\ : std_logic;
signal \N__29454\ : std_logic;
signal \N__29451\ : std_logic;
signal \N__29444\ : std_logic;
signal \N__29443\ : std_logic;
signal \N__29442\ : std_logic;
signal \N__29439\ : std_logic;
signal \N__29436\ : std_logic;
signal \N__29433\ : std_logic;
signal \N__29426\ : std_logic;
signal \N__29425\ : std_logic;
signal \N__29424\ : std_logic;
signal \N__29421\ : std_logic;
signal \N__29418\ : std_logic;
signal \N__29415\ : std_logic;
signal \N__29412\ : std_logic;
signal \N__29409\ : std_logic;
signal \N__29406\ : std_logic;
signal \N__29401\ : std_logic;
signal \N__29396\ : std_logic;
signal \N__29395\ : std_logic;
signal \N__29392\ : std_logic;
signal \N__29391\ : std_logic;
signal \N__29390\ : std_logic;
signal \N__29387\ : std_logic;
signal \N__29386\ : std_logic;
signal \N__29383\ : std_logic;
signal \N__29380\ : std_logic;
signal \N__29375\ : std_logic;
signal \N__29372\ : std_logic;
signal \N__29369\ : std_logic;
signal \N__29366\ : std_logic;
signal \N__29363\ : std_logic;
signal \N__29360\ : std_logic;
signal \N__29351\ : std_logic;
signal \N__29350\ : std_logic;
signal \N__29349\ : std_logic;
signal \N__29346\ : std_logic;
signal \N__29343\ : std_logic;
signal \N__29340\ : std_logic;
signal \N__29337\ : std_logic;
signal \N__29334\ : std_logic;
signal \N__29331\ : std_logic;
signal \N__29326\ : std_logic;
signal \N__29321\ : std_logic;
signal \N__29320\ : std_logic;
signal \N__29319\ : std_logic;
signal \N__29316\ : std_logic;
signal \N__29313\ : std_logic;
signal \N__29310\ : std_logic;
signal \N__29307\ : std_logic;
signal \N__29304\ : std_logic;
signal \N__29301\ : std_logic;
signal \N__29298\ : std_logic;
signal \N__29291\ : std_logic;
signal \N__29290\ : std_logic;
signal \N__29287\ : std_logic;
signal \N__29286\ : std_logic;
signal \N__29283\ : std_logic;
signal \N__29280\ : std_logic;
signal \N__29277\ : std_logic;
signal \N__29274\ : std_logic;
signal \N__29271\ : std_logic;
signal \N__29268\ : std_logic;
signal \N__29265\ : std_logic;
signal \N__29258\ : std_logic;
signal \N__29257\ : std_logic;
signal \N__29256\ : std_logic;
signal \N__29253\ : std_logic;
signal \N__29250\ : std_logic;
signal \N__29247\ : std_logic;
signal \N__29246\ : std_logic;
signal \N__29245\ : std_logic;
signal \N__29240\ : std_logic;
signal \N__29237\ : std_logic;
signal \N__29234\ : std_logic;
signal \N__29231\ : std_logic;
signal \N__29228\ : std_logic;
signal \N__29225\ : std_logic;
signal \N__29220\ : std_logic;
signal \N__29213\ : std_logic;
signal \N__29212\ : std_logic;
signal \N__29209\ : std_logic;
signal \N__29208\ : std_logic;
signal \N__29205\ : std_logic;
signal \N__29202\ : std_logic;
signal \N__29199\ : std_logic;
signal \N__29196\ : std_logic;
signal \N__29193\ : std_logic;
signal \N__29190\ : std_logic;
signal \N__29187\ : std_logic;
signal \N__29180\ : std_logic;
signal \N__29177\ : std_logic;
signal \N__29174\ : std_logic;
signal \N__29171\ : std_logic;
signal \N__29168\ : std_logic;
signal \N__29165\ : std_logic;
signal \N__29162\ : std_logic;
signal \N__29159\ : std_logic;
signal \N__29158\ : std_logic;
signal \N__29157\ : std_logic;
signal \N__29154\ : std_logic;
signal \N__29153\ : std_logic;
signal \N__29150\ : std_logic;
signal \N__29147\ : std_logic;
signal \N__29144\ : std_logic;
signal \N__29141\ : std_logic;
signal \N__29138\ : std_logic;
signal \N__29135\ : std_logic;
signal \N__29130\ : std_logic;
signal \N__29127\ : std_logic;
signal \N__29120\ : std_logic;
signal \N__29117\ : std_logic;
signal \N__29114\ : std_logic;
signal \N__29111\ : std_logic;
signal \N__29108\ : std_logic;
signal \N__29105\ : std_logic;
signal \N__29102\ : std_logic;
signal \N__29101\ : std_logic;
signal \N__29098\ : std_logic;
signal \N__29097\ : std_logic;
signal \N__29094\ : std_logic;
signal \N__29091\ : std_logic;
signal \N__29090\ : std_logic;
signal \N__29087\ : std_logic;
signal \N__29084\ : std_logic;
signal \N__29081\ : std_logic;
signal \N__29078\ : std_logic;
signal \N__29073\ : std_logic;
signal \N__29066\ : std_logic;
signal \N__29065\ : std_logic;
signal \N__29062\ : std_logic;
signal \N__29061\ : std_logic;
signal \N__29060\ : std_logic;
signal \N__29057\ : std_logic;
signal \N__29054\ : std_logic;
signal \N__29049\ : std_logic;
signal \N__29046\ : std_logic;
signal \N__29045\ : std_logic;
signal \N__29042\ : std_logic;
signal \N__29039\ : std_logic;
signal \N__29036\ : std_logic;
signal \N__29033\ : std_logic;
signal \N__29024\ : std_logic;
signal \N__29023\ : std_logic;
signal \N__29022\ : std_logic;
signal \N__29019\ : std_logic;
signal \N__29016\ : std_logic;
signal \N__29013\ : std_logic;
signal \N__29010\ : std_logic;
signal \N__29007\ : std_logic;
signal \N__29004\ : std_logic;
signal \N__29001\ : std_logic;
signal \N__28994\ : std_logic;
signal \N__28991\ : std_logic;
signal \N__28990\ : std_logic;
signal \N__28987\ : std_logic;
signal \N__28984\ : std_logic;
signal \N__28983\ : std_logic;
signal \N__28982\ : std_logic;
signal \N__28977\ : std_logic;
signal \N__28972\ : std_logic;
signal \N__28971\ : std_logic;
signal \N__28968\ : std_logic;
signal \N__28965\ : std_logic;
signal \N__28962\ : std_logic;
signal \N__28959\ : std_logic;
signal \N__28952\ : std_logic;
signal \N__28951\ : std_logic;
signal \N__28948\ : std_logic;
signal \N__28945\ : std_logic;
signal \N__28944\ : std_logic;
signal \N__28941\ : std_logic;
signal \N__28938\ : std_logic;
signal \N__28935\ : std_logic;
signal \N__28932\ : std_logic;
signal \N__28929\ : std_logic;
signal \N__28926\ : std_logic;
signal \N__28923\ : std_logic;
signal \N__28916\ : std_logic;
signal \N__28915\ : std_logic;
signal \N__28912\ : std_logic;
signal \N__28911\ : std_logic;
signal \N__28908\ : std_logic;
signal \N__28905\ : std_logic;
signal \N__28902\ : std_logic;
signal \N__28899\ : std_logic;
signal \N__28896\ : std_logic;
signal \N__28893\ : std_logic;
signal \N__28890\ : std_logic;
signal \N__28883\ : std_logic;
signal \N__28882\ : std_logic;
signal \N__28881\ : std_logic;
signal \N__28878\ : std_logic;
signal \N__28875\ : std_logic;
signal \N__28872\ : std_logic;
signal \N__28869\ : std_logic;
signal \N__28866\ : std_logic;
signal \N__28863\ : std_logic;
signal \N__28860\ : std_logic;
signal \N__28853\ : std_logic;
signal \N__28852\ : std_logic;
signal \N__28849\ : std_logic;
signal \N__28846\ : std_logic;
signal \N__28841\ : std_logic;
signal \N__28840\ : std_logic;
signal \N__28839\ : std_logic;
signal \N__28836\ : std_logic;
signal \N__28833\ : std_logic;
signal \N__28830\ : std_logic;
signal \N__28823\ : std_logic;
signal \N__28820\ : std_logic;
signal \N__28817\ : std_logic;
signal \N__28814\ : std_logic;
signal \N__28813\ : std_logic;
signal \N__28810\ : std_logic;
signal \N__28807\ : std_logic;
signal \N__28802\ : std_logic;
signal \N__28799\ : std_logic;
signal \N__28796\ : std_logic;
signal \N__28795\ : std_logic;
signal \N__28792\ : std_logic;
signal \N__28789\ : std_logic;
signal \N__28784\ : std_logic;
signal \N__28783\ : std_logic;
signal \N__28780\ : std_logic;
signal \N__28779\ : std_logic;
signal \N__28776\ : std_logic;
signal \N__28773\ : std_logic;
signal \N__28770\ : std_logic;
signal \N__28767\ : std_logic;
signal \N__28764\ : std_logic;
signal \N__28761\ : std_logic;
signal \N__28760\ : std_logic;
signal \N__28757\ : std_logic;
signal \N__28752\ : std_logic;
signal \N__28751\ : std_logic;
signal \N__28748\ : std_logic;
signal \N__28745\ : std_logic;
signal \N__28742\ : std_logic;
signal \N__28739\ : std_logic;
signal \N__28736\ : std_logic;
signal \N__28727\ : std_logic;
signal \N__28726\ : std_logic;
signal \N__28723\ : std_logic;
signal \N__28720\ : std_logic;
signal \N__28717\ : std_logic;
signal \N__28712\ : std_logic;
signal \N__28709\ : std_logic;
signal \N__28708\ : std_logic;
signal \N__28707\ : std_logic;
signal \N__28704\ : std_logic;
signal \N__28699\ : std_logic;
signal \N__28694\ : std_logic;
signal \N__28693\ : std_logic;
signal \N__28692\ : std_logic;
signal \N__28689\ : std_logic;
signal \N__28684\ : std_logic;
signal \N__28679\ : std_logic;
signal \N__28676\ : std_logic;
signal \N__28675\ : std_logic;
signal \N__28672\ : std_logic;
signal \N__28671\ : std_logic;
signal \N__28668\ : std_logic;
signal \N__28663\ : std_logic;
signal \N__28658\ : std_logic;
signal \N__28655\ : std_logic;
signal \N__28654\ : std_logic;
signal \N__28653\ : std_logic;
signal \N__28652\ : std_logic;
signal \N__28647\ : std_logic;
signal \N__28642\ : std_logic;
signal \N__28637\ : std_logic;
signal \N__28634\ : std_logic;
signal \N__28633\ : std_logic;
signal \N__28632\ : std_logic;
signal \N__28629\ : std_logic;
signal \N__28624\ : std_logic;
signal \N__28619\ : std_logic;
signal \N__28616\ : std_logic;
signal \N__28615\ : std_logic;
signal \N__28614\ : std_logic;
signal \N__28611\ : std_logic;
signal \N__28610\ : std_logic;
signal \N__28607\ : std_logic;
signal \N__28604\ : std_logic;
signal \N__28601\ : std_logic;
signal \N__28598\ : std_logic;
signal \N__28589\ : std_logic;
signal \N__28588\ : std_logic;
signal \N__28585\ : std_logic;
signal \N__28584\ : std_logic;
signal \N__28581\ : std_logic;
signal \N__28578\ : std_logic;
signal \N__28575\ : std_logic;
signal \N__28574\ : std_logic;
signal \N__28571\ : std_logic;
signal \N__28566\ : std_logic;
signal \N__28563\ : std_logic;
signal \N__28558\ : std_logic;
signal \N__28553\ : std_logic;
signal \N__28550\ : std_logic;
signal \N__28547\ : std_logic;
signal \N__28546\ : std_logic;
signal \N__28543\ : std_logic;
signal \N__28540\ : std_logic;
signal \N__28537\ : std_logic;
signal \N__28534\ : std_logic;
signal \N__28529\ : std_logic;
signal \N__28526\ : std_logic;
signal \N__28525\ : std_logic;
signal \N__28522\ : std_logic;
signal \N__28521\ : std_logic;
signal \N__28518\ : std_logic;
signal \N__28515\ : std_logic;
signal \N__28514\ : std_logic;
signal \N__28511\ : std_logic;
signal \N__28508\ : std_logic;
signal \N__28505\ : std_logic;
signal \N__28502\ : std_logic;
signal \N__28497\ : std_logic;
signal \N__28490\ : std_logic;
signal \N__28487\ : std_logic;
signal \N__28484\ : std_logic;
signal \N__28481\ : std_logic;
signal \N__28480\ : std_logic;
signal \N__28477\ : std_logic;
signal \N__28474\ : std_logic;
signal \N__28469\ : std_logic;
signal \N__28466\ : std_logic;
signal \N__28463\ : std_logic;
signal \N__28460\ : std_logic;
signal \N__28457\ : std_logic;
signal \N__28454\ : std_logic;
signal \N__28453\ : std_logic;
signal \N__28452\ : std_logic;
signal \N__28449\ : std_logic;
signal \N__28446\ : std_logic;
signal \N__28441\ : std_logic;
signal \N__28436\ : std_logic;
signal \N__28433\ : std_logic;
signal \N__28430\ : std_logic;
signal \N__28427\ : std_logic;
signal \N__28426\ : std_logic;
signal \N__28425\ : std_logic;
signal \N__28422\ : std_logic;
signal \N__28419\ : std_logic;
signal \N__28418\ : std_logic;
signal \N__28409\ : std_logic;
signal \N__28406\ : std_logic;
signal \N__28405\ : std_logic;
signal \N__28402\ : std_logic;
signal \N__28399\ : std_logic;
signal \N__28396\ : std_logic;
signal \N__28393\ : std_logic;
signal \N__28390\ : std_logic;
signal \N__28385\ : std_logic;
signal \N__28384\ : std_logic;
signal \N__28381\ : std_logic;
signal \N__28378\ : std_logic;
signal \N__28375\ : std_logic;
signal \N__28372\ : std_logic;
signal \N__28369\ : std_logic;
signal \N__28364\ : std_logic;
signal \N__28361\ : std_logic;
signal \N__28358\ : std_logic;
signal \N__28355\ : std_logic;
signal \N__28352\ : std_logic;
signal \N__28349\ : std_logic;
signal \N__28346\ : std_logic;
signal \N__28343\ : std_logic;
signal \N__28340\ : std_logic;
signal \N__28339\ : std_logic;
signal \N__28338\ : std_logic;
signal \N__28337\ : std_logic;
signal \N__28334\ : std_logic;
signal \N__28333\ : std_logic;
signal \N__28332\ : std_logic;
signal \N__28331\ : std_logic;
signal \N__28328\ : std_logic;
signal \N__28325\ : std_logic;
signal \N__28322\ : std_logic;
signal \N__28319\ : std_logic;
signal \N__28314\ : std_logic;
signal \N__28313\ : std_logic;
signal \N__28310\ : std_logic;
signal \N__28307\ : std_logic;
signal \N__28304\ : std_logic;
signal \N__28301\ : std_logic;
signal \N__28298\ : std_logic;
signal \N__28297\ : std_logic;
signal \N__28294\ : std_logic;
signal \N__28293\ : std_logic;
signal \N__28290\ : std_logic;
signal \N__28287\ : std_logic;
signal \N__28282\ : std_logic;
signal \N__28277\ : std_logic;
signal \N__28274\ : std_logic;
signal \N__28271\ : std_logic;
signal \N__28268\ : std_logic;
signal \N__28253\ : std_logic;
signal \N__28252\ : std_logic;
signal \N__28249\ : std_logic;
signal \N__28246\ : std_logic;
signal \N__28243\ : std_logic;
signal \N__28240\ : std_logic;
signal \N__28239\ : std_logic;
signal \N__28238\ : std_logic;
signal \N__28235\ : std_logic;
signal \N__28234\ : std_logic;
signal \N__28233\ : std_logic;
signal \N__28230\ : std_logic;
signal \N__28225\ : std_logic;
signal \N__28222\ : std_logic;
signal \N__28217\ : std_logic;
signal \N__28208\ : std_logic;
signal \N__28207\ : std_logic;
signal \N__28206\ : std_logic;
signal \N__28205\ : std_logic;
signal \N__28204\ : std_logic;
signal \N__28203\ : std_logic;
signal \N__28202\ : std_logic;
signal \N__28201\ : std_logic;
signal \N__28198\ : std_logic;
signal \N__28197\ : std_logic;
signal \N__28192\ : std_logic;
signal \N__28189\ : std_logic;
signal \N__28186\ : std_logic;
signal \N__28185\ : std_logic;
signal \N__28184\ : std_logic;
signal \N__28183\ : std_logic;
signal \N__28178\ : std_logic;
signal \N__28175\ : std_logic;
signal \N__28174\ : std_logic;
signal \N__28173\ : std_logic;
signal \N__28170\ : std_logic;
signal \N__28167\ : std_logic;
signal \N__28164\ : std_logic;
signal \N__28161\ : std_logic;
signal \N__28158\ : std_logic;
signal \N__28151\ : std_logic;
signal \N__28148\ : std_logic;
signal \N__28145\ : std_logic;
signal \N__28142\ : std_logic;
signal \N__28139\ : std_logic;
signal \N__28138\ : std_logic;
signal \N__28137\ : std_logic;
signal \N__28136\ : std_logic;
signal \N__28133\ : std_logic;
signal \N__28130\ : std_logic;
signal \N__28127\ : std_logic;
signal \N__28116\ : std_logic;
signal \N__28113\ : std_logic;
signal \N__28110\ : std_logic;
signal \N__28107\ : std_logic;
signal \N__28102\ : std_logic;
signal \N__28099\ : std_logic;
signal \N__28096\ : std_logic;
signal \N__28091\ : std_logic;
signal \N__28076\ : std_logic;
signal \N__28073\ : std_logic;
signal \N__28070\ : std_logic;
signal \N__28067\ : std_logic;
signal \N__28066\ : std_logic;
signal \N__28065\ : std_logic;
signal \N__28064\ : std_logic;
signal \N__28061\ : std_logic;
signal \N__28058\ : std_logic;
signal \N__28053\ : std_logic;
signal \N__28050\ : std_logic;
signal \N__28047\ : std_logic;
signal \N__28046\ : std_logic;
signal \N__28045\ : std_logic;
signal \N__28040\ : std_logic;
signal \N__28037\ : std_logic;
signal \N__28032\ : std_logic;
signal \N__28025\ : std_logic;
signal \N__28022\ : std_logic;
signal \N__28019\ : std_logic;
signal \N__28016\ : std_logic;
signal \N__28013\ : std_logic;
signal \N__28010\ : std_logic;
signal \N__28007\ : std_logic;
signal \N__28004\ : std_logic;
signal \N__28003\ : std_logic;
signal \N__27998\ : std_logic;
signal \N__27997\ : std_logic;
signal \N__27994\ : std_logic;
signal \N__27993\ : std_logic;
signal \N__27990\ : std_logic;
signal \N__27987\ : std_logic;
signal \N__27984\ : std_logic;
signal \N__27983\ : std_logic;
signal \N__27980\ : std_logic;
signal \N__27975\ : std_logic;
signal \N__27972\ : std_logic;
signal \N__27967\ : std_logic;
signal \N__27962\ : std_logic;
signal \N__27961\ : std_logic;
signal \N__27960\ : std_logic;
signal \N__27959\ : std_logic;
signal \N__27954\ : std_logic;
signal \N__27951\ : std_logic;
signal \N__27950\ : std_logic;
signal \N__27947\ : std_logic;
signal \N__27944\ : std_logic;
signal \N__27941\ : std_logic;
signal \N__27938\ : std_logic;
signal \N__27935\ : std_logic;
signal \N__27932\ : std_logic;
signal \N__27925\ : std_logic;
signal \N__27920\ : std_logic;
signal \N__27919\ : std_logic;
signal \N__27918\ : std_logic;
signal \N__27917\ : std_logic;
signal \N__27914\ : std_logic;
signal \N__27911\ : std_logic;
signal \N__27910\ : std_logic;
signal \N__27909\ : std_logic;
signal \N__27902\ : std_logic;
signal \N__27899\ : std_logic;
signal \N__27896\ : std_logic;
signal \N__27893\ : std_logic;
signal \N__27890\ : std_logic;
signal \N__27887\ : std_logic;
signal \N__27886\ : std_logic;
signal \N__27883\ : std_logic;
signal \N__27880\ : std_logic;
signal \N__27877\ : std_logic;
signal \N__27874\ : std_logic;
signal \N__27871\ : std_logic;
signal \N__27866\ : std_logic;
signal \N__27859\ : std_logic;
signal \N__27856\ : std_logic;
signal \N__27853\ : std_logic;
signal \N__27850\ : std_logic;
signal \N__27845\ : std_logic;
signal \N__27844\ : std_logic;
signal \N__27841\ : std_logic;
signal \N__27840\ : std_logic;
signal \N__27839\ : std_logic;
signal \N__27838\ : std_logic;
signal \N__27837\ : std_logic;
signal \N__27834\ : std_logic;
signal \N__27833\ : std_logic;
signal \N__27830\ : std_logic;
signal \N__27827\ : std_logic;
signal \N__27822\ : std_logic;
signal \N__27819\ : std_logic;
signal \N__27816\ : std_logic;
signal \N__27813\ : std_logic;
signal \N__27808\ : std_logic;
signal \N__27805\ : std_logic;
signal \N__27802\ : std_logic;
signal \N__27799\ : std_logic;
signal \N__27796\ : std_logic;
signal \N__27793\ : std_logic;
signal \N__27788\ : std_logic;
signal \N__27787\ : std_logic;
signal \N__27782\ : std_logic;
signal \N__27779\ : std_logic;
signal \N__27776\ : std_logic;
signal \N__27773\ : std_logic;
signal \N__27768\ : std_logic;
signal \N__27763\ : std_logic;
signal \N__27760\ : std_logic;
signal \N__27757\ : std_logic;
signal \N__27754\ : std_logic;
signal \N__27751\ : std_logic;
signal \N__27746\ : std_logic;
signal \N__27745\ : std_logic;
signal \N__27742\ : std_logic;
signal \N__27739\ : std_logic;
signal \N__27736\ : std_logic;
signal \N__27733\ : std_logic;
signal \N__27728\ : std_logic;
signal \N__27727\ : std_logic;
signal \N__27724\ : std_logic;
signal \N__27721\ : std_logic;
signal \N__27718\ : std_logic;
signal \N__27715\ : std_logic;
signal \N__27710\ : std_logic;
signal \N__27709\ : std_logic;
signal \N__27706\ : std_logic;
signal \N__27703\ : std_logic;
signal \N__27700\ : std_logic;
signal \N__27697\ : std_logic;
signal \N__27692\ : std_logic;
signal \N__27691\ : std_logic;
signal \N__27688\ : std_logic;
signal \N__27685\ : std_logic;
signal \N__27682\ : std_logic;
signal \N__27679\ : std_logic;
signal \N__27676\ : std_logic;
signal \N__27671\ : std_logic;
signal \N__27670\ : std_logic;
signal \N__27667\ : std_logic;
signal \N__27664\ : std_logic;
signal \N__27661\ : std_logic;
signal \N__27658\ : std_logic;
signal \N__27655\ : std_logic;
signal \N__27650\ : std_logic;
signal \N__27649\ : std_logic;
signal \N__27646\ : std_logic;
signal \N__27643\ : std_logic;
signal \N__27640\ : std_logic;
signal \N__27637\ : std_logic;
signal \N__27632\ : std_logic;
signal \N__27631\ : std_logic;
signal \N__27628\ : std_logic;
signal \N__27625\ : std_logic;
signal \N__27622\ : std_logic;
signal \N__27619\ : std_logic;
signal \N__27616\ : std_logic;
signal \N__27611\ : std_logic;
signal \N__27610\ : std_logic;
signal \N__27607\ : std_logic;
signal \N__27604\ : std_logic;
signal \N__27601\ : std_logic;
signal \N__27598\ : std_logic;
signal \N__27595\ : std_logic;
signal \N__27590\ : std_logic;
signal \N__27587\ : std_logic;
signal \N__27586\ : std_logic;
signal \N__27585\ : std_logic;
signal \N__27582\ : std_logic;
signal \N__27579\ : std_logic;
signal \N__27576\ : std_logic;
signal \N__27575\ : std_logic;
signal \N__27572\ : std_logic;
signal \N__27569\ : std_logic;
signal \N__27566\ : std_logic;
signal \N__27563\ : std_logic;
signal \N__27562\ : std_logic;
signal \N__27559\ : std_logic;
signal \N__27552\ : std_logic;
signal \N__27549\ : std_logic;
signal \N__27542\ : std_logic;
signal \N__27539\ : std_logic;
signal \N__27536\ : std_logic;
signal \N__27533\ : std_logic;
signal \N__27530\ : std_logic;
signal \N__27527\ : std_logic;
signal \N__27524\ : std_logic;
signal \N__27521\ : std_logic;
signal \N__27520\ : std_logic;
signal \N__27517\ : std_logic;
signal \N__27514\ : std_logic;
signal \N__27511\ : std_logic;
signal \N__27506\ : std_logic;
signal \N__27505\ : std_logic;
signal \N__27502\ : std_logic;
signal \N__27499\ : std_logic;
signal \N__27496\ : std_logic;
signal \N__27493\ : std_logic;
signal \N__27488\ : std_logic;
signal \N__27487\ : std_logic;
signal \N__27486\ : std_logic;
signal \N__27483\ : std_logic;
signal \N__27480\ : std_logic;
signal \N__27479\ : std_logic;
signal \N__27476\ : std_logic;
signal \N__27471\ : std_logic;
signal \N__27468\ : std_logic;
signal \N__27465\ : std_logic;
signal \N__27460\ : std_logic;
signal \N__27455\ : std_logic;
signal \N__27452\ : std_logic;
signal \N__27449\ : std_logic;
signal \N__27448\ : std_logic;
signal \N__27445\ : std_logic;
signal \N__27442\ : std_logic;
signal \N__27441\ : std_logic;
signal \N__27438\ : std_logic;
signal \N__27435\ : std_logic;
signal \N__27434\ : std_logic;
signal \N__27431\ : std_logic;
signal \N__27430\ : std_logic;
signal \N__27425\ : std_logic;
signal \N__27422\ : std_logic;
signal \N__27419\ : std_logic;
signal \N__27416\ : std_logic;
signal \N__27413\ : std_logic;
signal \N__27410\ : std_logic;
signal \N__27405\ : std_logic;
signal \N__27398\ : std_logic;
signal \N__27395\ : std_logic;
signal \N__27394\ : std_logic;
signal \N__27393\ : std_logic;
signal \N__27390\ : std_logic;
signal \N__27387\ : std_logic;
signal \N__27384\ : std_logic;
signal \N__27383\ : std_logic;
signal \N__27380\ : std_logic;
signal \N__27377\ : std_logic;
signal \N__27374\ : std_logic;
signal \N__27371\ : std_logic;
signal \N__27370\ : std_logic;
signal \N__27365\ : std_logic;
signal \N__27360\ : std_logic;
signal \N__27357\ : std_logic;
signal \N__27350\ : std_logic;
signal \N__27349\ : std_logic;
signal \N__27348\ : std_logic;
signal \N__27345\ : std_logic;
signal \N__27342\ : std_logic;
signal \N__27339\ : std_logic;
signal \N__27336\ : std_logic;
signal \N__27333\ : std_logic;
signal \N__27330\ : std_logic;
signal \N__27327\ : std_logic;
signal \N__27324\ : std_logic;
signal \N__27321\ : std_logic;
signal \N__27320\ : std_logic;
signal \N__27319\ : std_logic;
signal \N__27312\ : std_logic;
signal \N__27309\ : std_logic;
signal \N__27306\ : std_logic;
signal \N__27299\ : std_logic;
signal \N__27296\ : std_logic;
signal \N__27293\ : std_logic;
signal \N__27290\ : std_logic;
signal \N__27287\ : std_logic;
signal \N__27284\ : std_logic;
signal \N__27283\ : std_logic;
signal \N__27280\ : std_logic;
signal \N__27277\ : std_logic;
signal \N__27276\ : std_logic;
signal \N__27271\ : std_logic;
signal \N__27270\ : std_logic;
signal \N__27267\ : std_logic;
signal \N__27264\ : std_logic;
signal \N__27261\ : std_logic;
signal \N__27254\ : std_logic;
signal \N__27251\ : std_logic;
signal \N__27250\ : std_logic;
signal \N__27249\ : std_logic;
signal \N__27248\ : std_logic;
signal \N__27245\ : std_logic;
signal \N__27242\ : std_logic;
signal \N__27239\ : std_logic;
signal \N__27236\ : std_logic;
signal \N__27233\ : std_logic;
signal \N__27228\ : std_logic;
signal \N__27225\ : std_logic;
signal \N__27222\ : std_logic;
signal \N__27217\ : std_logic;
signal \N__27214\ : std_logic;
signal \N__27211\ : std_logic;
signal \N__27206\ : std_logic;
signal \N__27205\ : std_logic;
signal \N__27204\ : std_logic;
signal \N__27203\ : std_logic;
signal \N__27200\ : std_logic;
signal \N__27197\ : std_logic;
signal \N__27196\ : std_logic;
signal \N__27193\ : std_logic;
signal \N__27192\ : std_logic;
signal \N__27191\ : std_logic;
signal \N__27190\ : std_logic;
signal \N__27189\ : std_logic;
signal \N__27188\ : std_logic;
signal \N__27183\ : std_logic;
signal \N__27182\ : std_logic;
signal \N__27179\ : std_logic;
signal \N__27174\ : std_logic;
signal \N__27171\ : std_logic;
signal \N__27168\ : std_logic;
signal \N__27163\ : std_logic;
signal \N__27162\ : std_logic;
signal \N__27159\ : std_logic;
signal \N__27156\ : std_logic;
signal \N__27153\ : std_logic;
signal \N__27150\ : std_logic;
signal \N__27147\ : std_logic;
signal \N__27146\ : std_logic;
signal \N__27143\ : std_logic;
signal \N__27138\ : std_logic;
signal \N__27133\ : std_logic;
signal \N__27130\ : std_logic;
signal \N__27127\ : std_logic;
signal \N__27122\ : std_logic;
signal \N__27119\ : std_logic;
signal \N__27104\ : std_logic;
signal \N__27101\ : std_logic;
signal \N__27098\ : std_logic;
signal \N__27097\ : std_logic;
signal \N__27094\ : std_logic;
signal \N__27091\ : std_logic;
signal \N__27086\ : std_logic;
signal \N__27083\ : std_logic;
signal \N__27080\ : std_logic;
signal \N__27077\ : std_logic;
signal \N__27074\ : std_logic;
signal \N__27073\ : std_logic;
signal \N__27070\ : std_logic;
signal \N__27067\ : std_logic;
signal \N__27062\ : std_logic;
signal \N__27059\ : std_logic;
signal \N__27058\ : std_logic;
signal \N__27055\ : std_logic;
signal \N__27052\ : std_logic;
signal \N__27049\ : std_logic;
signal \N__27046\ : std_logic;
signal \N__27043\ : std_logic;
signal \N__27040\ : std_logic;
signal \N__27035\ : std_logic;
signal \N__27032\ : std_logic;
signal \N__27029\ : std_logic;
signal \N__27026\ : std_logic;
signal \N__27023\ : std_logic;
signal \N__27022\ : std_logic;
signal \N__27019\ : std_logic;
signal \N__27018\ : std_logic;
signal \N__27015\ : std_logic;
signal \N__27012\ : std_logic;
signal \N__27009\ : std_logic;
signal \N__27006\ : std_logic;
signal \N__26999\ : std_logic;
signal \N__26998\ : std_logic;
signal \N__26995\ : std_logic;
signal \N__26992\ : std_logic;
signal \N__26987\ : std_logic;
signal \N__26986\ : std_logic;
signal \N__26983\ : std_logic;
signal \N__26982\ : std_logic;
signal \N__26979\ : std_logic;
signal \N__26976\ : std_logic;
signal \N__26971\ : std_logic;
signal \N__26966\ : std_logic;
signal \N__26965\ : std_logic;
signal \N__26962\ : std_logic;
signal \N__26959\ : std_logic;
signal \N__26954\ : std_logic;
signal \N__26951\ : std_logic;
signal \N__26950\ : std_logic;
signal \N__26947\ : std_logic;
signal \N__26944\ : std_logic;
signal \N__26941\ : std_logic;
signal \N__26938\ : std_logic;
signal \N__26935\ : std_logic;
signal \N__26934\ : std_logic;
signal \N__26929\ : std_logic;
signal \N__26926\ : std_logic;
signal \N__26921\ : std_logic;
signal \N__26918\ : std_logic;
signal \N__26915\ : std_logic;
signal \N__26912\ : std_logic;
signal \N__26909\ : std_logic;
signal \N__26906\ : std_logic;
signal \N__26903\ : std_logic;
signal \N__26902\ : std_logic;
signal \N__26901\ : std_logic;
signal \N__26900\ : std_logic;
signal \N__26899\ : std_logic;
signal \N__26898\ : std_logic;
signal \N__26897\ : std_logic;
signal \N__26894\ : std_logic;
signal \N__26891\ : std_logic;
signal \N__26886\ : std_logic;
signal \N__26885\ : std_logic;
signal \N__26884\ : std_logic;
signal \N__26883\ : std_logic;
signal \N__26882\ : std_logic;
signal \N__26881\ : std_logic;
signal \N__26878\ : std_logic;
signal \N__26875\ : std_logic;
signal \N__26874\ : std_logic;
signal \N__26871\ : std_logic;
signal \N__26866\ : std_logic;
signal \N__26863\ : std_logic;
signal \N__26856\ : std_logic;
signal \N__26851\ : std_logic;
signal \N__26848\ : std_logic;
signal \N__26845\ : std_logic;
signal \N__26842\ : std_logic;
signal \N__26837\ : std_logic;
signal \N__26828\ : std_logic;
signal \N__26819\ : std_logic;
signal \N__26816\ : std_logic;
signal \N__26813\ : std_logic;
signal \N__26810\ : std_logic;
signal \N__26807\ : std_logic;
signal \N__26804\ : std_logic;
signal \N__26801\ : std_logic;
signal \N__26800\ : std_logic;
signal \N__26797\ : std_logic;
signal \N__26796\ : std_logic;
signal \N__26793\ : std_logic;
signal \N__26790\ : std_logic;
signal \N__26785\ : std_logic;
signal \N__26780\ : std_logic;
signal \N__26777\ : std_logic;
signal \N__26774\ : std_logic;
signal \N__26773\ : std_logic;
signal \N__26770\ : std_logic;
signal \N__26767\ : std_logic;
signal \N__26762\ : std_logic;
signal \N__26761\ : std_logic;
signal \N__26758\ : std_logic;
signal \N__26755\ : std_logic;
signal \N__26752\ : std_logic;
signal \N__26749\ : std_logic;
signal \N__26744\ : std_logic;
signal \N__26741\ : std_logic;
signal \N__26738\ : std_logic;
signal \N__26737\ : std_logic;
signal \N__26734\ : std_logic;
signal \N__26731\ : std_logic;
signal \N__26728\ : std_logic;
signal \N__26725\ : std_logic;
signal \N__26720\ : std_logic;
signal \N__26717\ : std_logic;
signal \N__26716\ : std_logic;
signal \N__26713\ : std_logic;
signal \N__26712\ : std_logic;
signal \N__26709\ : std_logic;
signal \N__26706\ : std_logic;
signal \N__26703\ : std_logic;
signal \N__26700\ : std_logic;
signal \N__26697\ : std_logic;
signal \N__26690\ : std_logic;
signal \N__26689\ : std_logic;
signal \N__26686\ : std_logic;
signal \N__26683\ : std_logic;
signal \N__26678\ : std_logic;
signal \N__26675\ : std_logic;
signal \N__26674\ : std_logic;
signal \N__26671\ : std_logic;
signal \N__26668\ : std_logic;
signal \N__26665\ : std_logic;
signal \N__26660\ : std_logic;
signal \N__26657\ : std_logic;
signal \N__26654\ : std_logic;
signal \N__26651\ : std_logic;
signal \N__26648\ : std_logic;
signal \N__26647\ : std_logic;
signal \N__26644\ : std_logic;
signal \N__26641\ : std_logic;
signal \N__26638\ : std_logic;
signal \N__26635\ : std_logic;
signal \N__26630\ : std_logic;
signal \N__26627\ : std_logic;
signal \N__26624\ : std_logic;
signal \N__26621\ : std_logic;
signal \N__26618\ : std_logic;
signal \N__26617\ : std_logic;
signal \N__26614\ : std_logic;
signal \N__26611\ : std_logic;
signal \N__26608\ : std_logic;
signal \N__26603\ : std_logic;
signal \N__26600\ : std_logic;
signal \N__26597\ : std_logic;
signal \N__26594\ : std_logic;
signal \N__26591\ : std_logic;
signal \N__26590\ : std_logic;
signal \N__26587\ : std_logic;
signal \N__26584\ : std_logic;
signal \N__26579\ : std_logic;
signal \N__26576\ : std_logic;
signal \N__26573\ : std_logic;
signal \N__26570\ : std_logic;
signal \N__26569\ : std_logic;
signal \N__26566\ : std_logic;
signal \N__26563\ : std_logic;
signal \N__26558\ : std_logic;
signal \N__26555\ : std_logic;
signal \N__26552\ : std_logic;
signal \N__26551\ : std_logic;
signal \N__26548\ : std_logic;
signal \N__26545\ : std_logic;
signal \N__26540\ : std_logic;
signal \N__26537\ : std_logic;
signal \N__26534\ : std_logic;
signal \N__26531\ : std_logic;
signal \N__26528\ : std_logic;
signal \N__26527\ : std_logic;
signal \N__26526\ : std_logic;
signal \N__26525\ : std_logic;
signal \N__26524\ : std_logic;
signal \N__26523\ : std_logic;
signal \N__26522\ : std_logic;
signal \N__26521\ : std_logic;
signal \N__26520\ : std_logic;
signal \N__26519\ : std_logic;
signal \N__26518\ : std_logic;
signal \N__26503\ : std_logic;
signal \N__26500\ : std_logic;
signal \N__26493\ : std_logic;
signal \N__26490\ : std_logic;
signal \N__26485\ : std_logic;
signal \N__26482\ : std_logic;
signal \N__26479\ : std_logic;
signal \N__26476\ : std_logic;
signal \N__26473\ : std_logic;
signal \N__26470\ : std_logic;
signal \N__26467\ : std_logic;
signal \N__26462\ : std_logic;
signal \N__26459\ : std_logic;
signal \N__26458\ : std_logic;
signal \N__26455\ : std_logic;
signal \N__26452\ : std_logic;
signal \N__26451\ : std_logic;
signal \N__26450\ : std_logic;
signal \N__26449\ : std_logic;
signal \N__26446\ : std_logic;
signal \N__26443\ : std_logic;
signal \N__26442\ : std_logic;
signal \N__26441\ : std_logic;
signal \N__26436\ : std_logic;
signal \N__26433\ : std_logic;
signal \N__26430\ : std_logic;
signal \N__26427\ : std_logic;
signal \N__26422\ : std_logic;
signal \N__26417\ : std_logic;
signal \N__26408\ : std_logic;
signal \N__26405\ : std_logic;
signal \N__26402\ : std_logic;
signal \N__26399\ : std_logic;
signal \N__26396\ : std_logic;
signal \N__26393\ : std_logic;
signal \N__26390\ : std_logic;
signal \N__26387\ : std_logic;
signal \N__26384\ : std_logic;
signal \N__26381\ : std_logic;
signal \N__26378\ : std_logic;
signal \N__26375\ : std_logic;
signal \N__26372\ : std_logic;
signal \N__26369\ : std_logic;
signal \N__26366\ : std_logic;
signal \N__26363\ : std_logic;
signal \N__26360\ : std_logic;
signal \N__26357\ : std_logic;
signal \N__26354\ : std_logic;
signal \N__26351\ : std_logic;
signal \N__26348\ : std_logic;
signal \N__26345\ : std_logic;
signal \N__26342\ : std_logic;
signal \N__26339\ : std_logic;
signal \N__26336\ : std_logic;
signal \N__26333\ : std_logic;
signal \N__26330\ : std_logic;
signal \N__26327\ : std_logic;
signal \N__26324\ : std_logic;
signal \N__26321\ : std_logic;
signal \N__26318\ : std_logic;
signal \N__26315\ : std_logic;
signal \N__26312\ : std_logic;
signal \N__26309\ : std_logic;
signal \N__26306\ : std_logic;
signal \N__26303\ : std_logic;
signal \N__26300\ : std_logic;
signal \N__26297\ : std_logic;
signal \N__26294\ : std_logic;
signal \N__26291\ : std_logic;
signal \N__26288\ : std_logic;
signal \N__26285\ : std_logic;
signal \N__26282\ : std_logic;
signal \N__26279\ : std_logic;
signal \N__26276\ : std_logic;
signal \N__26273\ : std_logic;
signal \N__26270\ : std_logic;
signal \N__26267\ : std_logic;
signal \N__26264\ : std_logic;
signal \N__26261\ : std_logic;
signal \N__26260\ : std_logic;
signal \N__26257\ : std_logic;
signal \N__26254\ : std_logic;
signal \N__26251\ : std_logic;
signal \N__26248\ : std_logic;
signal \N__26245\ : std_logic;
signal \N__26242\ : std_logic;
signal \N__26239\ : std_logic;
signal \N__26236\ : std_logic;
signal \N__26233\ : std_logic;
signal \N__26230\ : std_logic;
signal \N__26225\ : std_logic;
signal \N__26222\ : std_logic;
signal \N__26221\ : std_logic;
signal \N__26218\ : std_logic;
signal \N__26215\ : std_logic;
signal \N__26210\ : std_logic;
signal \N__26207\ : std_logic;
signal \N__26206\ : std_logic;
signal \N__26205\ : std_logic;
signal \N__26202\ : std_logic;
signal \N__26199\ : std_logic;
signal \N__26198\ : std_logic;
signal \N__26197\ : std_logic;
signal \N__26194\ : std_logic;
signal \N__26191\ : std_logic;
signal \N__26190\ : std_logic;
signal \N__26187\ : std_logic;
signal \N__26184\ : std_logic;
signal \N__26181\ : std_logic;
signal \N__26180\ : std_logic;
signal \N__26177\ : std_logic;
signal \N__26174\ : std_logic;
signal \N__26171\ : std_logic;
signal \N__26168\ : std_logic;
signal \N__26163\ : std_logic;
signal \N__26160\ : std_logic;
signal \N__26153\ : std_logic;
signal \N__26150\ : std_logic;
signal \N__26145\ : std_logic;
signal \N__26144\ : std_logic;
signal \N__26141\ : std_logic;
signal \N__26136\ : std_logic;
signal \N__26133\ : std_logic;
signal \N__26130\ : std_logic;
signal \N__26127\ : std_logic;
signal \N__26124\ : std_logic;
signal \N__26121\ : std_logic;
signal \N__26116\ : std_logic;
signal \N__26111\ : std_logic;
signal \N__26108\ : std_logic;
signal \N__26105\ : std_logic;
signal \N__26102\ : std_logic;
signal \N__26099\ : std_logic;
signal \N__26096\ : std_logic;
signal \N__26093\ : std_logic;
signal \N__26090\ : std_logic;
signal \N__26087\ : std_logic;
signal \N__26084\ : std_logic;
signal \N__26081\ : std_logic;
signal \N__26078\ : std_logic;
signal \N__26075\ : std_logic;
signal \N__26074\ : std_logic;
signal \N__26071\ : std_logic;
signal \N__26068\ : std_logic;
signal \N__26067\ : std_logic;
signal \N__26062\ : std_logic;
signal \N__26061\ : std_logic;
signal \N__26060\ : std_logic;
signal \N__26057\ : std_logic;
signal \N__26054\ : std_logic;
signal \N__26051\ : std_logic;
signal \N__26048\ : std_logic;
signal \N__26045\ : std_logic;
signal \N__26042\ : std_logic;
signal \N__26033\ : std_logic;
signal \N__26032\ : std_logic;
signal \N__26031\ : std_logic;
signal \N__26028\ : std_logic;
signal \N__26025\ : std_logic;
signal \N__26022\ : std_logic;
signal \N__26021\ : std_logic;
signal \N__26018\ : std_logic;
signal \N__26015\ : std_logic;
signal \N__26014\ : std_logic;
signal \N__26011\ : std_logic;
signal \N__26008\ : std_logic;
signal \N__26005\ : std_logic;
signal \N__26004\ : std_logic;
signal \N__26001\ : std_logic;
signal \N__25998\ : std_logic;
signal \N__25995\ : std_logic;
signal \N__25992\ : std_logic;
signal \N__25989\ : std_logic;
signal \N__25986\ : std_logic;
signal \N__25981\ : std_logic;
signal \N__25978\ : std_logic;
signal \N__25975\ : std_logic;
signal \N__25970\ : std_logic;
signal \N__25963\ : std_logic;
signal \N__25958\ : std_logic;
signal \N__25957\ : std_logic;
signal \N__25956\ : std_logic;
signal \N__25955\ : std_logic;
signal \N__25954\ : std_logic;
signal \N__25953\ : std_logic;
signal \N__25952\ : std_logic;
signal \N__25951\ : std_logic;
signal \N__25942\ : std_logic;
signal \N__25939\ : std_logic;
signal \N__25936\ : std_logic;
signal \N__25935\ : std_logic;
signal \N__25934\ : std_logic;
signal \N__25933\ : std_logic;
signal \N__25930\ : std_logic;
signal \N__25927\ : std_logic;
signal \N__25922\ : std_logic;
signal \N__25919\ : std_logic;
signal \N__25916\ : std_logic;
signal \N__25913\ : std_logic;
signal \N__25912\ : std_logic;
signal \N__25911\ : std_logic;
signal \N__25910\ : std_logic;
signal \N__25909\ : std_logic;
signal \N__25906\ : std_logic;
signal \N__25903\ : std_logic;
signal \N__25900\ : std_logic;
signal \N__25899\ : std_logic;
signal \N__25896\ : std_logic;
signal \N__25893\ : std_logic;
signal \N__25890\ : std_logic;
signal \N__25887\ : std_logic;
signal \N__25876\ : std_logic;
signal \N__25873\ : std_logic;
signal \N__25870\ : std_logic;
signal \N__25867\ : std_logic;
signal \N__25864\ : std_logic;
signal \N__25861\ : std_logic;
signal \N__25858\ : std_logic;
signal \N__25853\ : std_logic;
signal \N__25850\ : std_logic;
signal \N__25847\ : std_logic;
signal \N__25844\ : std_logic;
signal \N__25829\ : std_logic;
signal \N__25828\ : std_logic;
signal \N__25827\ : std_logic;
signal \N__25824\ : std_logic;
signal \N__25821\ : std_logic;
signal \N__25818\ : std_logic;
signal \N__25817\ : std_logic;
signal \N__25816\ : std_logic;
signal \N__25815\ : std_logic;
signal \N__25814\ : std_logic;
signal \N__25807\ : std_logic;
signal \N__25804\ : std_logic;
signal \N__25799\ : std_logic;
signal \N__25796\ : std_logic;
signal \N__25793\ : std_logic;
signal \N__25784\ : std_logic;
signal \N__25781\ : std_logic;
signal \N__25778\ : std_logic;
signal \N__25775\ : std_logic;
signal \N__25774\ : std_logic;
signal \N__25771\ : std_logic;
signal \N__25768\ : std_logic;
signal \N__25763\ : std_logic;
signal \N__25760\ : std_logic;
signal \N__25757\ : std_logic;
signal \N__25754\ : std_logic;
signal \N__25751\ : std_logic;
signal \N__25748\ : std_logic;
signal \N__25745\ : std_logic;
signal \N__25742\ : std_logic;
signal \N__25739\ : std_logic;
signal \N__25738\ : std_logic;
signal \N__25735\ : std_logic;
signal \N__25732\ : std_logic;
signal \N__25731\ : std_logic;
signal \N__25728\ : std_logic;
signal \N__25725\ : std_logic;
signal \N__25724\ : std_logic;
signal \N__25723\ : std_logic;
signal \N__25722\ : std_logic;
signal \N__25721\ : std_logic;
signal \N__25718\ : std_logic;
signal \N__25713\ : std_logic;
signal \N__25708\ : std_logic;
signal \N__25701\ : std_logic;
signal \N__25698\ : std_logic;
signal \N__25691\ : std_logic;
signal \N__25688\ : std_logic;
signal \N__25687\ : std_logic;
signal \N__25686\ : std_logic;
signal \N__25685\ : std_logic;
signal \N__25682\ : std_logic;
signal \N__25679\ : std_logic;
signal \N__25676\ : std_logic;
signal \N__25673\ : std_logic;
signal \N__25672\ : std_logic;
signal \N__25667\ : std_logic;
signal \N__25664\ : std_logic;
signal \N__25661\ : std_logic;
signal \N__25658\ : std_logic;
signal \N__25655\ : std_logic;
signal \N__25650\ : std_logic;
signal \N__25647\ : std_logic;
signal \N__25640\ : std_logic;
signal \N__25639\ : std_logic;
signal \N__25636\ : std_logic;
signal \N__25635\ : std_logic;
signal \N__25634\ : std_logic;
signal \N__25633\ : std_logic;
signal \N__25632\ : std_logic;
signal \N__25629\ : std_logic;
signal \N__25628\ : std_logic;
signal \N__25625\ : std_logic;
signal \N__25624\ : std_logic;
signal \N__25617\ : std_logic;
signal \N__25614\ : std_logic;
signal \N__25609\ : std_logic;
signal \N__25606\ : std_logic;
signal \N__25603\ : std_logic;
signal \N__25598\ : std_logic;
signal \N__25595\ : std_logic;
signal \N__25590\ : std_logic;
signal \N__25587\ : std_logic;
signal \N__25584\ : std_logic;
signal \N__25577\ : std_logic;
signal \N__25574\ : std_logic;
signal \N__25571\ : std_logic;
signal \N__25568\ : std_logic;
signal \N__25565\ : std_logic;
signal \N__25562\ : std_logic;
signal \N__25559\ : std_logic;
signal \N__25556\ : std_logic;
signal \N__25553\ : std_logic;
signal \N__25550\ : std_logic;
signal \N__25547\ : std_logic;
signal \N__25544\ : std_logic;
signal \N__25541\ : std_logic;
signal \N__25538\ : std_logic;
signal \N__25537\ : std_logic;
signal \N__25532\ : std_logic;
signal \N__25531\ : std_logic;
signal \N__25530\ : std_logic;
signal \N__25529\ : std_logic;
signal \N__25528\ : std_logic;
signal \N__25525\ : std_logic;
signal \N__25524\ : std_logic;
signal \N__25521\ : std_logic;
signal \N__25516\ : std_logic;
signal \N__25513\ : std_logic;
signal \N__25510\ : std_logic;
signal \N__25505\ : std_logic;
signal \N__25502\ : std_logic;
signal \N__25495\ : std_logic;
signal \N__25492\ : std_logic;
signal \N__25489\ : std_logic;
signal \N__25484\ : std_logic;
signal \N__25483\ : std_logic;
signal \N__25480\ : std_logic;
signal \N__25477\ : std_logic;
signal \N__25474\ : std_logic;
signal \N__25471\ : std_logic;
signal \N__25470\ : std_logic;
signal \N__25469\ : std_logic;
signal \N__25464\ : std_logic;
signal \N__25459\ : std_logic;
signal \N__25458\ : std_logic;
signal \N__25457\ : std_logic;
signal \N__25454\ : std_logic;
signal \N__25451\ : std_logic;
signal \N__25446\ : std_logic;
signal \N__25439\ : std_logic;
signal \N__25438\ : std_logic;
signal \N__25437\ : std_logic;
signal \N__25434\ : std_logic;
signal \N__25431\ : std_logic;
signal \N__25428\ : std_logic;
signal \N__25423\ : std_logic;
signal \N__25420\ : std_logic;
signal \N__25419\ : std_logic;
signal \N__25418\ : std_logic;
signal \N__25417\ : std_logic;
signal \N__25416\ : std_logic;
signal \N__25413\ : std_logic;
signal \N__25410\ : std_logic;
signal \N__25407\ : std_logic;
signal \N__25400\ : std_logic;
signal \N__25397\ : std_logic;
signal \N__25388\ : std_logic;
signal \N__25385\ : std_logic;
signal \N__25382\ : std_logic;
signal \N__25379\ : std_logic;
signal \N__25376\ : std_logic;
signal \N__25373\ : std_logic;
signal \N__25370\ : std_logic;
signal \N__25367\ : std_logic;
signal \N__25366\ : std_logic;
signal \N__25365\ : std_logic;
signal \N__25364\ : std_logic;
signal \N__25363\ : std_logic;
signal \N__25360\ : std_logic;
signal \N__25359\ : std_logic;
signal \N__25358\ : std_logic;
signal \N__25355\ : std_logic;
signal \N__25350\ : std_logic;
signal \N__25349\ : std_logic;
signal \N__25348\ : std_logic;
signal \N__25347\ : std_logic;
signal \N__25344\ : std_logic;
signal \N__25341\ : std_logic;
signal \N__25340\ : std_logic;
signal \N__25339\ : std_logic;
signal \N__25336\ : std_logic;
signal \N__25333\ : std_logic;
signal \N__25330\ : std_logic;
signal \N__25327\ : std_logic;
signal \N__25324\ : std_logic;
signal \N__25321\ : std_logic;
signal \N__25316\ : std_logic;
signal \N__25313\ : std_logic;
signal \N__25308\ : std_logic;
signal \N__25301\ : std_logic;
signal \N__25286\ : std_logic;
signal \N__25283\ : std_logic;
signal \N__25280\ : std_logic;
signal \N__25277\ : std_logic;
signal \N__25274\ : std_logic;
signal \N__25271\ : std_logic;
signal \N__25268\ : std_logic;
signal \N__25267\ : std_logic;
signal \N__25264\ : std_logic;
signal \N__25261\ : std_logic;
signal \N__25260\ : std_logic;
signal \N__25259\ : std_logic;
signal \N__25258\ : std_logic;
signal \N__25257\ : std_logic;
signal \N__25256\ : std_logic;
signal \N__25255\ : std_logic;
signal \N__25254\ : std_logic;
signal \N__25253\ : std_logic;
signal \N__25250\ : std_logic;
signal \N__25249\ : std_logic;
signal \N__25248\ : std_logic;
signal \N__25245\ : std_logic;
signal \N__25242\ : std_logic;
signal \N__25237\ : std_logic;
signal \N__25234\ : std_logic;
signal \N__25231\ : std_logic;
signal \N__25228\ : std_logic;
signal \N__25225\ : std_logic;
signal \N__25222\ : std_logic;
signal \N__25219\ : std_logic;
signal \N__25214\ : std_logic;
signal \N__25207\ : std_logic;
signal \N__25202\ : std_logic;
signal \N__25187\ : std_logic;
signal \N__25184\ : std_logic;
signal \N__25181\ : std_logic;
signal \N__25178\ : std_logic;
signal \N__25175\ : std_logic;
signal \N__25172\ : std_logic;
signal \N__25169\ : std_logic;
signal \N__25166\ : std_logic;
signal \N__25163\ : std_logic;
signal \N__25160\ : std_logic;
signal \N__25157\ : std_logic;
signal \N__25154\ : std_logic;
signal \N__25151\ : std_logic;
signal \N__25148\ : std_logic;
signal \N__25145\ : std_logic;
signal \N__25142\ : std_logic;
signal \N__25141\ : std_logic;
signal \N__25138\ : std_logic;
signal \N__25135\ : std_logic;
signal \N__25132\ : std_logic;
signal \N__25129\ : std_logic;
signal \N__25126\ : std_logic;
signal \N__25123\ : std_logic;
signal \N__25120\ : std_logic;
signal \N__25117\ : std_logic;
signal \N__25112\ : std_logic;
signal \N__25109\ : std_logic;
signal \N__25106\ : std_logic;
signal \N__25105\ : std_logic;
signal \N__25102\ : std_logic;
signal \N__25099\ : std_logic;
signal \N__25096\ : std_logic;
signal \N__25093\ : std_logic;
signal \N__25088\ : std_logic;
signal \N__25085\ : std_logic;
signal \N__25082\ : std_logic;
signal \N__25079\ : std_logic;
signal \N__25076\ : std_logic;
signal \N__25073\ : std_logic;
signal \N__25070\ : std_logic;
signal \N__25067\ : std_logic;
signal \N__25064\ : std_logic;
signal \N__25061\ : std_logic;
signal \N__25058\ : std_logic;
signal \N__25057\ : std_logic;
signal \N__25054\ : std_logic;
signal \N__25051\ : std_logic;
signal \N__25048\ : std_logic;
signal \N__25045\ : std_logic;
signal \N__25042\ : std_logic;
signal \N__25039\ : std_logic;
signal \N__25034\ : std_logic;
signal \N__25031\ : std_logic;
signal \N__25028\ : std_logic;
signal \N__25025\ : std_logic;
signal \N__25022\ : std_logic;
signal \N__25019\ : std_logic;
signal \N__25016\ : std_logic;
signal \N__25013\ : std_logic;
signal \N__25010\ : std_logic;
signal \N__25009\ : std_logic;
signal \N__25006\ : std_logic;
signal \N__25003\ : std_logic;
signal \N__25000\ : std_logic;
signal \N__24995\ : std_logic;
signal \N__24992\ : std_logic;
signal \N__24989\ : std_logic;
signal \N__24986\ : std_logic;
signal \N__24983\ : std_logic;
signal \N__24980\ : std_logic;
signal \N__24977\ : std_logic;
signal \N__24976\ : std_logic;
signal \N__24973\ : std_logic;
signal \N__24970\ : std_logic;
signal \N__24967\ : std_logic;
signal \N__24964\ : std_logic;
signal \N__24961\ : std_logic;
signal \N__24958\ : std_logic;
signal \N__24955\ : std_logic;
signal \N__24952\ : std_logic;
signal \N__24947\ : std_logic;
signal \N__24944\ : std_logic;
signal \N__24943\ : std_logic;
signal \N__24940\ : std_logic;
signal \N__24937\ : std_logic;
signal \N__24932\ : std_logic;
signal \N__24929\ : std_logic;
signal \N__24926\ : std_logic;
signal \N__24923\ : std_logic;
signal \N__24920\ : std_logic;
signal \N__24917\ : std_logic;
signal \N__24914\ : std_logic;
signal \N__24911\ : std_logic;
signal \N__24908\ : std_logic;
signal \N__24907\ : std_logic;
signal \N__24904\ : std_logic;
signal \N__24901\ : std_logic;
signal \N__24898\ : std_logic;
signal \N__24893\ : std_logic;
signal \N__24890\ : std_logic;
signal \N__24887\ : std_logic;
signal \N__24884\ : std_logic;
signal \N__24881\ : std_logic;
signal \N__24880\ : std_logic;
signal \N__24877\ : std_logic;
signal \N__24874\ : std_logic;
signal \N__24871\ : std_logic;
signal \N__24866\ : std_logic;
signal \N__24863\ : std_logic;
signal \N__24860\ : std_logic;
signal \N__24857\ : std_logic;
signal \N__24854\ : std_logic;
signal \N__24851\ : std_logic;
signal \N__24848\ : std_logic;
signal \N__24845\ : std_logic;
signal \N__24842\ : std_logic;
signal \N__24839\ : std_logic;
signal \N__24836\ : std_logic;
signal \N__24835\ : std_logic;
signal \N__24832\ : std_logic;
signal \N__24829\ : std_logic;
signal \N__24826\ : std_logic;
signal \N__24823\ : std_logic;
signal \N__24820\ : std_logic;
signal \N__24815\ : std_logic;
signal \N__24812\ : std_logic;
signal \N__24809\ : std_logic;
signal \N__24806\ : std_logic;
signal \N__24803\ : std_logic;
signal \N__24800\ : std_logic;
signal \N__24797\ : std_logic;
signal \N__24794\ : std_logic;
signal \N__24791\ : std_logic;
signal \N__24790\ : std_logic;
signal \N__24787\ : std_logic;
signal \N__24784\ : std_logic;
signal \N__24779\ : std_logic;
signal \N__24776\ : std_logic;
signal \N__24773\ : std_logic;
signal \N__24770\ : std_logic;
signal \N__24767\ : std_logic;
signal \N__24764\ : std_logic;
signal \N__24763\ : std_logic;
signal \N__24760\ : std_logic;
signal \N__24757\ : std_logic;
signal \N__24754\ : std_logic;
signal \N__24751\ : std_logic;
signal \N__24746\ : std_logic;
signal \N__24743\ : std_logic;
signal \N__24740\ : std_logic;
signal \N__24737\ : std_logic;
signal \N__24734\ : std_logic;
signal \N__24731\ : std_logic;
signal \N__24728\ : std_logic;
signal \N__24727\ : std_logic;
signal \N__24724\ : std_logic;
signal \N__24721\ : std_logic;
signal \N__24718\ : std_logic;
signal \N__24715\ : std_logic;
signal \N__24710\ : std_logic;
signal \N__24707\ : std_logic;
signal \N__24704\ : std_logic;
signal \N__24701\ : std_logic;
signal \N__24698\ : std_logic;
signal \N__24695\ : std_logic;
signal \N__24692\ : std_logic;
signal \N__24689\ : std_logic;
signal \N__24686\ : std_logic;
signal \N__24683\ : std_logic;
signal \N__24680\ : std_logic;
signal \N__24677\ : std_logic;
signal \N__24674\ : std_logic;
signal \N__24671\ : std_logic;
signal \N__24668\ : std_logic;
signal \N__24665\ : std_logic;
signal \N__24662\ : std_logic;
signal \N__24661\ : std_logic;
signal \N__24660\ : std_logic;
signal \N__24659\ : std_logic;
signal \N__24658\ : std_logic;
signal \N__24653\ : std_logic;
signal \N__24650\ : std_logic;
signal \N__24647\ : std_logic;
signal \N__24644\ : std_logic;
signal \N__24639\ : std_logic;
signal \N__24634\ : std_logic;
signal \N__24629\ : std_logic;
signal \N__24626\ : std_logic;
signal \N__24623\ : std_logic;
signal \N__24620\ : std_logic;
signal \N__24617\ : std_logic;
signal \N__24614\ : std_logic;
signal \N__24611\ : std_logic;
signal \N__24608\ : std_logic;
signal \N__24605\ : std_logic;
signal \N__24602\ : std_logic;
signal \N__24599\ : std_logic;
signal \N__24596\ : std_logic;
signal \N__24593\ : std_logic;
signal \N__24592\ : std_logic;
signal \N__24591\ : std_logic;
signal \N__24590\ : std_logic;
signal \N__24587\ : std_logic;
signal \N__24584\ : std_logic;
signal \N__24581\ : std_logic;
signal \N__24578\ : std_logic;
signal \N__24575\ : std_logic;
signal \N__24570\ : std_logic;
signal \N__24567\ : std_logic;
signal \N__24560\ : std_logic;
signal \N__24559\ : std_logic;
signal \N__24558\ : std_logic;
signal \N__24551\ : std_logic;
signal \N__24550\ : std_logic;
signal \N__24549\ : std_logic;
signal \N__24548\ : std_logic;
signal \N__24545\ : std_logic;
signal \N__24540\ : std_logic;
signal \N__24537\ : std_logic;
signal \N__24530\ : std_logic;
signal \N__24527\ : std_logic;
signal \N__24524\ : std_logic;
signal \N__24523\ : std_logic;
signal \N__24522\ : std_logic;
signal \N__24521\ : std_logic;
signal \N__24516\ : std_logic;
signal \N__24515\ : std_logic;
signal \N__24514\ : std_logic;
signal \N__24513\ : std_logic;
signal \N__24508\ : std_logic;
signal \N__24505\ : std_logic;
signal \N__24500\ : std_logic;
signal \N__24497\ : std_logic;
signal \N__24488\ : std_logic;
signal \N__24487\ : std_logic;
signal \N__24484\ : std_logic;
signal \N__24481\ : std_logic;
signal \N__24478\ : std_logic;
signal \N__24477\ : std_logic;
signal \N__24476\ : std_logic;
signal \N__24475\ : std_logic;
signal \N__24470\ : std_logic;
signal \N__24467\ : std_logic;
signal \N__24466\ : std_logic;
signal \N__24463\ : std_logic;
signal \N__24460\ : std_logic;
signal \N__24457\ : std_logic;
signal \N__24452\ : std_logic;
signal \N__24449\ : std_logic;
signal \N__24446\ : std_logic;
signal \N__24437\ : std_logic;
signal \N__24434\ : std_logic;
signal \N__24431\ : std_logic;
signal \N__24428\ : std_logic;
signal \N__24425\ : std_logic;
signal \N__24422\ : std_logic;
signal \N__24421\ : std_logic;
signal \N__24418\ : std_logic;
signal \N__24415\ : std_logic;
signal \N__24412\ : std_logic;
signal \N__24409\ : std_logic;
signal \N__24404\ : std_logic;
signal \N__24401\ : std_logic;
signal \N__24398\ : std_logic;
signal \N__24395\ : std_logic;
signal \N__24392\ : std_logic;
signal \N__24389\ : std_logic;
signal \N__24388\ : std_logic;
signal \N__24385\ : std_logic;
signal \N__24382\ : std_logic;
signal \N__24379\ : std_logic;
signal \N__24376\ : std_logic;
signal \N__24371\ : std_logic;
signal \N__24368\ : std_logic;
signal \N__24365\ : std_logic;
signal \N__24362\ : std_logic;
signal \N__24359\ : std_logic;
signal \N__24356\ : std_logic;
signal \N__24353\ : std_logic;
signal \N__24350\ : std_logic;
signal \N__24347\ : std_logic;
signal \N__24344\ : std_logic;
signal \N__24343\ : std_logic;
signal \N__24340\ : std_logic;
signal \N__24335\ : std_logic;
signal \N__24332\ : std_logic;
signal \N__24329\ : std_logic;
signal \N__24326\ : std_logic;
signal \N__24323\ : std_logic;
signal \N__24320\ : std_logic;
signal \N__24317\ : std_logic;
signal \N__24314\ : std_logic;
signal \N__24311\ : std_logic;
signal \N__24308\ : std_logic;
signal \N__24305\ : std_logic;
signal \N__24302\ : std_logic;
signal \N__24299\ : std_logic;
signal \N__24296\ : std_logic;
signal \N__24293\ : std_logic;
signal \N__24290\ : std_logic;
signal \N__24287\ : std_logic;
signal \N__24284\ : std_logic;
signal \N__24281\ : std_logic;
signal \N__24280\ : std_logic;
signal \N__24277\ : std_logic;
signal \N__24276\ : std_logic;
signal \N__24275\ : std_logic;
signal \N__24274\ : std_logic;
signal \N__24273\ : std_logic;
signal \N__24270\ : std_logic;
signal \N__24267\ : std_logic;
signal \N__24258\ : std_logic;
signal \N__24257\ : std_logic;
signal \N__24256\ : std_logic;
signal \N__24255\ : std_logic;
signal \N__24254\ : std_logic;
signal \N__24251\ : std_logic;
signal \N__24246\ : std_logic;
signal \N__24237\ : std_logic;
signal \N__24230\ : std_logic;
signal \N__24227\ : std_logic;
signal \N__24226\ : std_logic;
signal \N__24223\ : std_logic;
signal \N__24220\ : std_logic;
signal \N__24217\ : std_logic;
signal \N__24214\ : std_logic;
signal \N__24209\ : std_logic;
signal \N__24206\ : std_logic;
signal \N__24205\ : std_logic;
signal \N__24202\ : std_logic;
signal \N__24199\ : std_logic;
signal \N__24196\ : std_logic;
signal \N__24193\ : std_logic;
signal \N__24188\ : std_logic;
signal \N__24185\ : std_logic;
signal \N__24182\ : std_logic;
signal \N__24181\ : std_logic;
signal \N__24180\ : std_logic;
signal \N__24179\ : std_logic;
signal \N__24176\ : std_logic;
signal \N__24173\ : std_logic;
signal \N__24170\ : std_logic;
signal \N__24167\ : std_logic;
signal \N__24162\ : std_logic;
signal \N__24159\ : std_logic;
signal \N__24156\ : std_logic;
signal \N__24153\ : std_logic;
signal \N__24150\ : std_logic;
signal \N__24147\ : std_logic;
signal \N__24144\ : std_logic;
signal \N__24137\ : std_logic;
signal \N__24134\ : std_logic;
signal \N__24131\ : std_logic;
signal \N__24128\ : std_logic;
signal \N__24125\ : std_logic;
signal \N__24122\ : std_logic;
signal \N__24119\ : std_logic;
signal \N__24116\ : std_logic;
signal \N__24113\ : std_logic;
signal \N__24110\ : std_logic;
signal \N__24107\ : std_logic;
signal \N__24104\ : std_logic;
signal \N__24101\ : std_logic;
signal \N__24098\ : std_logic;
signal \N__24095\ : std_logic;
signal \N__24092\ : std_logic;
signal \N__24089\ : std_logic;
signal \N__24088\ : std_logic;
signal \N__24085\ : std_logic;
signal \N__24082\ : std_logic;
signal \N__24079\ : std_logic;
signal \N__24076\ : std_logic;
signal \N__24073\ : std_logic;
signal \N__24070\ : std_logic;
signal \N__24067\ : std_logic;
signal \N__24064\ : std_logic;
signal \N__24059\ : std_logic;
signal \N__24056\ : std_logic;
signal \N__24053\ : std_logic;
signal \N__24050\ : std_logic;
signal \N__24047\ : std_logic;
signal \N__24044\ : std_logic;
signal \N__24041\ : std_logic;
signal \N__24038\ : std_logic;
signal \N__24035\ : std_logic;
signal \N__24032\ : std_logic;
signal \N__24029\ : std_logic;
signal \N__24026\ : std_logic;
signal \N__24023\ : std_logic;
signal \N__24020\ : std_logic;
signal \N__24017\ : std_logic;
signal \N__24014\ : std_logic;
signal \N__24011\ : std_logic;
signal \N__24008\ : std_logic;
signal \N__24005\ : std_logic;
signal \N__24002\ : std_logic;
signal \N__23999\ : std_logic;
signal \N__23996\ : std_logic;
signal \N__23993\ : std_logic;
signal \N__23990\ : std_logic;
signal \N__23987\ : std_logic;
signal \N__23984\ : std_logic;
signal \N__23981\ : std_logic;
signal \N__23978\ : std_logic;
signal \N__23977\ : std_logic;
signal \N__23976\ : std_logic;
signal \N__23973\ : std_logic;
signal \N__23970\ : std_logic;
signal \N__23969\ : std_logic;
signal \N__23968\ : std_logic;
signal \N__23967\ : std_logic;
signal \N__23966\ : std_logic;
signal \N__23963\ : std_logic;
signal \N__23960\ : std_logic;
signal \N__23951\ : std_logic;
signal \N__23950\ : std_logic;
signal \N__23949\ : std_logic;
signal \N__23948\ : std_logic;
signal \N__23945\ : std_logic;
signal \N__23942\ : std_logic;
signal \N__23939\ : std_logic;
signal \N__23936\ : std_logic;
signal \N__23929\ : std_logic;
signal \N__23926\ : std_logic;
signal \N__23921\ : std_logic;
signal \N__23916\ : std_logic;
signal \N__23915\ : std_logic;
signal \N__23914\ : std_logic;
signal \N__23913\ : std_logic;
signal \N__23912\ : std_logic;
signal \N__23909\ : std_logic;
signal \N__23904\ : std_logic;
signal \N__23899\ : std_logic;
signal \N__23894\ : std_logic;
signal \N__23885\ : std_logic;
signal \N__23882\ : std_logic;
signal \N__23879\ : std_logic;
signal \N__23876\ : std_logic;
signal \N__23875\ : std_logic;
signal \N__23874\ : std_logic;
signal \N__23873\ : std_logic;
signal \N__23872\ : std_logic;
signal \N__23871\ : std_logic;
signal \N__23870\ : std_logic;
signal \N__23869\ : std_logic;
signal \N__23868\ : std_logic;
signal \N__23867\ : std_logic;
signal \N__23866\ : std_logic;
signal \N__23865\ : std_logic;
signal \N__23862\ : std_logic;
signal \N__23847\ : std_logic;
signal \N__23838\ : std_logic;
signal \N__23835\ : std_logic;
signal \N__23828\ : std_logic;
signal \N__23825\ : std_logic;
signal \N__23822\ : std_logic;
signal \N__23819\ : std_logic;
signal \N__23818\ : std_logic;
signal \N__23815\ : std_logic;
signal \N__23812\ : std_logic;
signal \N__23809\ : std_logic;
signal \N__23804\ : std_logic;
signal \N__23801\ : std_logic;
signal \N__23800\ : std_logic;
signal \N__23799\ : std_logic;
signal \N__23796\ : std_logic;
signal \N__23793\ : std_logic;
signal \N__23790\ : std_logic;
signal \N__23785\ : std_logic;
signal \N__23782\ : std_logic;
signal \N__23779\ : std_logic;
signal \N__23774\ : std_logic;
signal \N__23771\ : std_logic;
signal \N__23768\ : std_logic;
signal \N__23765\ : std_logic;
signal \N__23764\ : std_logic;
signal \N__23763\ : std_logic;
signal \N__23756\ : std_logic;
signal \N__23753\ : std_logic;
signal \N__23750\ : std_logic;
signal \N__23749\ : std_logic;
signal \N__23748\ : std_logic;
signal \N__23745\ : std_logic;
signal \N__23742\ : std_logic;
signal \N__23739\ : std_logic;
signal \N__23736\ : std_logic;
signal \N__23733\ : std_logic;
signal \N__23726\ : std_logic;
signal \N__23723\ : std_logic;
signal \N__23720\ : std_logic;
signal \N__23719\ : std_logic;
signal \N__23718\ : std_logic;
signal \N__23715\ : std_logic;
signal \N__23710\ : std_logic;
signal \N__23705\ : std_logic;
signal \N__23704\ : std_logic;
signal \N__23701\ : std_logic;
signal \N__23698\ : std_logic;
signal \N__23695\ : std_logic;
signal \N__23692\ : std_logic;
signal \N__23687\ : std_logic;
signal \N__23684\ : std_logic;
signal \N__23681\ : std_logic;
signal \N__23678\ : std_logic;
signal \N__23675\ : std_logic;
signal \N__23674\ : std_logic;
signal \N__23671\ : std_logic;
signal \N__23668\ : std_logic;
signal \N__23665\ : std_logic;
signal \N__23662\ : std_logic;
signal \N__23659\ : std_logic;
signal \N__23654\ : std_logic;
signal \N__23653\ : std_logic;
signal \N__23650\ : std_logic;
signal \N__23647\ : std_logic;
signal \N__23644\ : std_logic;
signal \N__23641\ : std_logic;
signal \N__23638\ : std_logic;
signal \N__23635\ : std_logic;
signal \N__23632\ : std_logic;
signal \N__23629\ : std_logic;
signal \N__23626\ : std_logic;
signal \N__23621\ : std_logic;
signal \N__23618\ : std_logic;
signal \N__23615\ : std_logic;
signal \N__23612\ : std_logic;
signal \N__23609\ : std_logic;
signal \N__23606\ : std_logic;
signal \N__23603\ : std_logic;
signal \N__23600\ : std_logic;
signal \N__23597\ : std_logic;
signal \N__23594\ : std_logic;
signal \N__23591\ : std_logic;
signal \N__23588\ : std_logic;
signal \N__23585\ : std_logic;
signal \N__23582\ : std_logic;
signal \N__23579\ : std_logic;
signal \N__23576\ : std_logic;
signal \N__23573\ : std_logic;
signal \N__23570\ : std_logic;
signal \N__23567\ : std_logic;
signal \N__23564\ : std_logic;
signal \N__23561\ : std_logic;
signal \N__23558\ : std_logic;
signal \N__23555\ : std_logic;
signal \N__23552\ : std_logic;
signal \N__23549\ : std_logic;
signal \N__23546\ : std_logic;
signal \N__23543\ : std_logic;
signal \N__23540\ : std_logic;
signal \N__23537\ : std_logic;
signal \N__23534\ : std_logic;
signal \N__23531\ : std_logic;
signal \N__23528\ : std_logic;
signal \N__23525\ : std_logic;
signal \N__23522\ : std_logic;
signal \N__23519\ : std_logic;
signal \N__23516\ : std_logic;
signal \N__23513\ : std_logic;
signal \N__23512\ : std_logic;
signal \N__23509\ : std_logic;
signal \N__23506\ : std_logic;
signal \N__23501\ : std_logic;
signal \N__23498\ : std_logic;
signal \N__23497\ : std_logic;
signal \N__23496\ : std_logic;
signal \N__23493\ : std_logic;
signal \N__23488\ : std_logic;
signal \N__23483\ : std_logic;
signal \N__23480\ : std_logic;
signal \N__23477\ : std_logic;
signal \N__23474\ : std_logic;
signal \N__23471\ : std_logic;
signal \N__23468\ : std_logic;
signal \N__23465\ : std_logic;
signal \N__23462\ : std_logic;
signal \N__23459\ : std_logic;
signal \N__23458\ : std_logic;
signal \N__23455\ : std_logic;
signal \N__23452\ : std_logic;
signal \N__23451\ : std_logic;
signal \N__23450\ : std_logic;
signal \N__23447\ : std_logic;
signal \N__23440\ : std_logic;
signal \N__23435\ : std_logic;
signal \N__23432\ : std_logic;
signal \N__23431\ : std_logic;
signal \N__23430\ : std_logic;
signal \N__23427\ : std_logic;
signal \N__23424\ : std_logic;
signal \N__23423\ : std_logic;
signal \N__23420\ : std_logic;
signal \N__23417\ : std_logic;
signal \N__23410\ : std_logic;
signal \N__23405\ : std_logic;
signal \N__23404\ : std_logic;
signal \N__23401\ : std_logic;
signal \N__23398\ : std_logic;
signal \N__23395\ : std_logic;
signal \N__23392\ : std_logic;
signal \N__23389\ : std_logic;
signal \N__23386\ : std_logic;
signal \N__23383\ : std_logic;
signal \N__23380\ : std_logic;
signal \N__23377\ : std_logic;
signal \N__23372\ : std_logic;
signal \N__23371\ : std_logic;
signal \N__23368\ : std_logic;
signal \N__23365\ : std_logic;
signal \N__23362\ : std_logic;
signal \N__23359\ : std_logic;
signal \N__23356\ : std_logic;
signal \N__23353\ : std_logic;
signal \N__23350\ : std_logic;
signal \N__23347\ : std_logic;
signal \N__23344\ : std_logic;
signal \N__23341\ : std_logic;
signal \N__23336\ : std_logic;
signal \N__23333\ : std_logic;
signal \N__23332\ : std_logic;
signal \N__23329\ : std_logic;
signal \N__23326\ : std_logic;
signal \N__23323\ : std_logic;
signal \N__23320\ : std_logic;
signal \N__23317\ : std_logic;
signal \N__23314\ : std_logic;
signal \N__23311\ : std_logic;
signal \N__23308\ : std_logic;
signal \N__23305\ : std_logic;
signal \N__23300\ : std_logic;
signal \N__23299\ : std_logic;
signal \N__23298\ : std_logic;
signal \N__23297\ : std_logic;
signal \N__23296\ : std_logic;
signal \N__23293\ : std_logic;
signal \N__23288\ : std_logic;
signal \N__23285\ : std_logic;
signal \N__23282\ : std_logic;
signal \N__23273\ : std_logic;
signal \N__23272\ : std_logic;
signal \N__23269\ : std_logic;
signal \N__23268\ : std_logic;
signal \N__23265\ : std_logic;
signal \N__23262\ : std_logic;
signal \N__23259\ : std_logic;
signal \N__23256\ : std_logic;
signal \N__23249\ : std_logic;
signal \N__23248\ : std_logic;
signal \N__23245\ : std_logic;
signal \N__23242\ : std_logic;
signal \N__23239\ : std_logic;
signal \N__23234\ : std_logic;
signal \N__23233\ : std_logic;
signal \N__23230\ : std_logic;
signal \N__23227\ : std_logic;
signal \N__23224\ : std_logic;
signal \N__23219\ : std_logic;
signal \N__23216\ : std_logic;
signal \N__23215\ : std_logic;
signal \N__23212\ : std_logic;
signal \N__23209\ : std_logic;
signal \N__23206\ : std_logic;
signal \N__23201\ : std_logic;
signal \N__23200\ : std_logic;
signal \N__23197\ : std_logic;
signal \N__23194\ : std_logic;
signal \N__23189\ : std_logic;
signal \N__23186\ : std_logic;
signal \N__23185\ : std_logic;
signal \N__23182\ : std_logic;
signal \N__23179\ : std_logic;
signal \N__23176\ : std_logic;
signal \N__23171\ : std_logic;
signal \N__23170\ : std_logic;
signal \N__23167\ : std_logic;
signal \N__23164\ : std_logic;
signal \N__23159\ : std_logic;
signal \N__23156\ : std_logic;
signal \N__23153\ : std_logic;
signal \N__23152\ : std_logic;
signal \N__23149\ : std_logic;
signal \N__23146\ : std_logic;
signal \N__23141\ : std_logic;
signal \N__23138\ : std_logic;
signal \N__23135\ : std_logic;
signal \N__23132\ : std_logic;
signal \N__23131\ : std_logic;
signal \N__23128\ : std_logic;
signal \N__23125\ : std_logic;
signal \N__23120\ : std_logic;
signal \N__23117\ : std_logic;
signal \N__23116\ : std_logic;
signal \N__23113\ : std_logic;
signal \N__23110\ : std_logic;
signal \N__23107\ : std_logic;
signal \N__23104\ : std_logic;
signal \N__23099\ : std_logic;
signal \N__23096\ : std_logic;
signal \N__23093\ : std_logic;
signal \N__23092\ : std_logic;
signal \N__23089\ : std_logic;
signal \N__23086\ : std_logic;
signal \N__23081\ : std_logic;
signal \N__23078\ : std_logic;
signal \N__23075\ : std_logic;
signal \N__23074\ : std_logic;
signal \N__23071\ : std_logic;
signal \N__23068\ : std_logic;
signal \N__23065\ : std_logic;
signal \N__23060\ : std_logic;
signal \N__23057\ : std_logic;
signal \N__23056\ : std_logic;
signal \N__23055\ : std_logic;
signal \N__23052\ : std_logic;
signal \N__23047\ : std_logic;
signal \N__23042\ : std_logic;
signal \N__23039\ : std_logic;
signal \N__23036\ : std_logic;
signal \N__23033\ : std_logic;
signal \N__23030\ : std_logic;
signal \N__23027\ : std_logic;
signal \N__23024\ : std_logic;
signal \N__23021\ : std_logic;
signal \N__23018\ : std_logic;
signal \N__23017\ : std_logic;
signal \N__23016\ : std_logic;
signal \N__23015\ : std_logic;
signal \N__23014\ : std_logic;
signal \N__23011\ : std_logic;
signal \N__23006\ : std_logic;
signal \N__23005\ : std_logic;
signal \N__23004\ : std_logic;
signal \N__23001\ : std_logic;
signal \N__23000\ : std_logic;
signal \N__22997\ : std_logic;
signal \N__22996\ : std_logic;
signal \N__22995\ : std_logic;
signal \N__22994\ : std_logic;
signal \N__22993\ : std_logic;
signal \N__22992\ : std_logic;
signal \N__22989\ : std_logic;
signal \N__22986\ : std_logic;
signal \N__22979\ : std_logic;
signal \N__22972\ : std_logic;
signal \N__22969\ : std_logic;
signal \N__22968\ : std_logic;
signal \N__22963\ : std_logic;
signal \N__22960\ : std_logic;
signal \N__22951\ : std_logic;
signal \N__22946\ : std_logic;
signal \N__22937\ : std_logic;
signal \N__22936\ : std_logic;
signal \N__22933\ : std_logic;
signal \N__22930\ : std_logic;
signal \N__22925\ : std_logic;
signal \N__22924\ : std_logic;
signal \N__22923\ : std_logic;
signal \N__22920\ : std_logic;
signal \N__22917\ : std_logic;
signal \N__22916\ : std_logic;
signal \N__22915\ : std_logic;
signal \N__22912\ : std_logic;
signal \N__22909\ : std_logic;
signal \N__22908\ : std_logic;
signal \N__22907\ : std_logic;
signal \N__22904\ : std_logic;
signal \N__22897\ : std_logic;
signal \N__22894\ : std_logic;
signal \N__22893\ : std_logic;
signal \N__22890\ : std_logic;
signal \N__22887\ : std_logic;
signal \N__22884\ : std_logic;
signal \N__22881\ : std_logic;
signal \N__22878\ : std_logic;
signal \N__22875\ : std_logic;
signal \N__22872\ : std_logic;
signal \N__22869\ : std_logic;
signal \N__22864\ : std_logic;
signal \N__22863\ : std_logic;
signal \N__22862\ : std_logic;
signal \N__22859\ : std_logic;
signal \N__22856\ : std_logic;
signal \N__22853\ : std_logic;
signal \N__22848\ : std_logic;
signal \N__22843\ : std_logic;
signal \N__22832\ : std_logic;
signal \N__22831\ : std_logic;
signal \N__22830\ : std_logic;
signal \N__22829\ : std_logic;
signal \N__22828\ : std_logic;
signal \N__22827\ : std_logic;
signal \N__22826\ : std_logic;
signal \N__22823\ : std_logic;
signal \N__22820\ : std_logic;
signal \N__22817\ : std_logic;
signal \N__22816\ : std_logic;
signal \N__22813\ : std_logic;
signal \N__22812\ : std_logic;
signal \N__22809\ : std_logic;
signal \N__22804\ : std_logic;
signal \N__22801\ : std_logic;
signal \N__22796\ : std_logic;
signal \N__22793\ : std_logic;
signal \N__22790\ : std_logic;
signal \N__22787\ : std_logic;
signal \N__22786\ : std_logic;
signal \N__22785\ : std_logic;
signal \N__22782\ : std_logic;
signal \N__22777\ : std_logic;
signal \N__22770\ : std_logic;
signal \N__22767\ : std_logic;
signal \N__22762\ : std_logic;
signal \N__22759\ : std_logic;
signal \N__22756\ : std_logic;
signal \N__22753\ : std_logic;
signal \N__22748\ : std_logic;
signal \N__22739\ : std_logic;
signal \N__22738\ : std_logic;
signal \N__22737\ : std_logic;
signal \N__22734\ : std_logic;
signal \N__22733\ : std_logic;
signal \N__22728\ : std_logic;
signal \N__22725\ : std_logic;
signal \N__22724\ : std_logic;
signal \N__22721\ : std_logic;
signal \N__22720\ : std_logic;
signal \N__22717\ : std_logic;
signal \N__22714\ : std_logic;
signal \N__22713\ : std_logic;
signal \N__22710\ : std_logic;
signal \N__22707\ : std_logic;
signal \N__22704\ : std_logic;
signal \N__22701\ : std_logic;
signal \N__22698\ : std_logic;
signal \N__22695\ : std_logic;
signal \N__22690\ : std_logic;
signal \N__22685\ : std_logic;
signal \N__22676\ : std_logic;
signal \N__22673\ : std_logic;
signal \N__22670\ : std_logic;
signal \N__22667\ : std_logic;
signal \N__22664\ : std_logic;
signal \N__22661\ : std_logic;
signal \N__22658\ : std_logic;
signal \N__22655\ : std_logic;
signal \N__22652\ : std_logic;
signal \N__22649\ : std_logic;
signal \N__22646\ : std_logic;
signal \N__22643\ : std_logic;
signal \N__22642\ : std_logic;
signal \N__22639\ : std_logic;
signal \N__22638\ : std_logic;
signal \N__22635\ : std_logic;
signal \N__22634\ : std_logic;
signal \N__22631\ : std_logic;
signal \N__22628\ : std_logic;
signal \N__22627\ : std_logic;
signal \N__22626\ : std_logic;
signal \N__22625\ : std_logic;
signal \N__22624\ : std_logic;
signal \N__22621\ : std_logic;
signal \N__22620\ : std_logic;
signal \N__22619\ : std_logic;
signal \N__22616\ : std_logic;
signal \N__22611\ : std_logic;
signal \N__22608\ : std_logic;
signal \N__22601\ : std_logic;
signal \N__22598\ : std_logic;
signal \N__22593\ : std_logic;
signal \N__22590\ : std_logic;
signal \N__22583\ : std_logic;
signal \N__22580\ : std_logic;
signal \N__22577\ : std_logic;
signal \N__22574\ : std_logic;
signal \N__22573\ : std_logic;
signal \N__22570\ : std_logic;
signal \N__22567\ : std_logic;
signal \N__22564\ : std_logic;
signal \N__22561\ : std_logic;
signal \N__22558\ : std_logic;
signal \N__22555\ : std_logic;
signal \N__22544\ : std_logic;
signal \N__22541\ : std_logic;
signal \N__22538\ : std_logic;
signal \N__22535\ : std_logic;
signal \N__22532\ : std_logic;
signal \N__22531\ : std_logic;
signal \N__22528\ : std_logic;
signal \N__22527\ : std_logic;
signal \N__22526\ : std_logic;
signal \N__22525\ : std_logic;
signal \N__22524\ : std_logic;
signal \N__22523\ : std_logic;
signal \N__22520\ : std_logic;
signal \N__22515\ : std_logic;
signal \N__22512\ : std_logic;
signal \N__22511\ : std_logic;
signal \N__22508\ : std_logic;
signal \N__22505\ : std_logic;
signal \N__22502\ : std_logic;
signal \N__22501\ : std_logic;
signal \N__22500\ : std_logic;
signal \N__22499\ : std_logic;
signal \N__22494\ : std_logic;
signal \N__22491\ : std_logic;
signal \N__22488\ : std_logic;
signal \N__22481\ : std_logic;
signal \N__22476\ : std_logic;
signal \N__22473\ : std_logic;
signal \N__22460\ : std_logic;
signal \N__22457\ : std_logic;
signal \N__22454\ : std_logic;
signal \N__22451\ : std_logic;
signal \N__22448\ : std_logic;
signal \N__22445\ : std_logic;
signal \N__22444\ : std_logic;
signal \N__22443\ : std_logic;
signal \N__22440\ : std_logic;
signal \N__22439\ : std_logic;
signal \N__22438\ : std_logic;
signal \N__22435\ : std_logic;
signal \N__22432\ : std_logic;
signal \N__22431\ : std_logic;
signal \N__22430\ : std_logic;
signal \N__22429\ : std_logic;
signal \N__22426\ : std_logic;
signal \N__22421\ : std_logic;
signal \N__22420\ : std_logic;
signal \N__22415\ : std_logic;
signal \N__22410\ : std_logic;
signal \N__22407\ : std_logic;
signal \N__22406\ : std_logic;
signal \N__22405\ : std_logic;
signal \N__22404\ : std_logic;
signal \N__22399\ : std_logic;
signal \N__22396\ : std_logic;
signal \N__22389\ : std_logic;
signal \N__22386\ : std_logic;
signal \N__22381\ : std_logic;
signal \N__22370\ : std_logic;
signal \N__22367\ : std_logic;
signal \N__22364\ : std_logic;
signal \N__22361\ : std_logic;
signal \N__22358\ : std_logic;
signal \N__22355\ : std_logic;
signal \N__22352\ : std_logic;
signal \N__22349\ : std_logic;
signal \N__22346\ : std_logic;
signal \N__22343\ : std_logic;
signal \N__22340\ : std_logic;
signal \N__22337\ : std_logic;
signal \N__22334\ : std_logic;
signal \N__22331\ : std_logic;
signal \N__22328\ : std_logic;
signal \N__22325\ : std_logic;
signal \N__22322\ : std_logic;
signal \N__22319\ : std_logic;
signal \N__22316\ : std_logic;
signal \N__22313\ : std_logic;
signal \N__22310\ : std_logic;
signal \N__22307\ : std_logic;
signal \N__22304\ : std_logic;
signal \N__22301\ : std_logic;
signal \N__22298\ : std_logic;
signal \N__22295\ : std_logic;
signal \N__22292\ : std_logic;
signal \N__22289\ : std_logic;
signal \N__22286\ : std_logic;
signal \N__22283\ : std_logic;
signal \N__22280\ : std_logic;
signal \N__22277\ : std_logic;
signal \N__22274\ : std_logic;
signal \N__22271\ : std_logic;
signal \N__22270\ : std_logic;
signal \N__22267\ : std_logic;
signal \N__22266\ : std_logic;
signal \N__22259\ : std_logic;
signal \N__22256\ : std_logic;
signal \N__22253\ : std_logic;
signal \N__22250\ : std_logic;
signal \N__22249\ : std_logic;
signal \N__22248\ : std_logic;
signal \N__22245\ : std_logic;
signal \N__22238\ : std_logic;
signal \N__22237\ : std_logic;
signal \N__22234\ : std_logic;
signal \N__22231\ : std_logic;
signal \N__22228\ : std_logic;
signal \N__22225\ : std_logic;
signal \N__22222\ : std_logic;
signal \N__22217\ : std_logic;
signal \N__22214\ : std_logic;
signal \N__22211\ : std_logic;
signal \N__22208\ : std_logic;
signal \N__22205\ : std_logic;
signal \N__22202\ : std_logic;
signal \N__22199\ : std_logic;
signal \N__22196\ : std_logic;
signal \N__22195\ : std_logic;
signal \N__22192\ : std_logic;
signal \N__22189\ : std_logic;
signal \N__22188\ : std_logic;
signal \N__22187\ : std_logic;
signal \N__22186\ : std_logic;
signal \N__22183\ : std_logic;
signal \N__22180\ : std_logic;
signal \N__22177\ : std_logic;
signal \N__22174\ : std_logic;
signal \N__22171\ : std_logic;
signal \N__22170\ : std_logic;
signal \N__22169\ : std_logic;
signal \N__22166\ : std_logic;
signal \N__22163\ : std_logic;
signal \N__22160\ : std_logic;
signal \N__22157\ : std_logic;
signal \N__22154\ : std_logic;
signal \N__22151\ : std_logic;
signal \N__22150\ : std_logic;
signal \N__22149\ : std_logic;
signal \N__22146\ : std_logic;
signal \N__22139\ : std_logic;
signal \N__22136\ : std_logic;
signal \N__22131\ : std_logic;
signal \N__22128\ : std_logic;
signal \N__22125\ : std_logic;
signal \N__22122\ : std_logic;
signal \N__22109\ : std_logic;
signal \N__22108\ : std_logic;
signal \N__22107\ : std_logic;
signal \N__22106\ : std_logic;
signal \N__22097\ : std_logic;
signal \N__22096\ : std_logic;
signal \N__22095\ : std_logic;
signal \N__22092\ : std_logic;
signal \N__22089\ : std_logic;
signal \N__22088\ : std_logic;
signal \N__22087\ : std_logic;
signal \N__22086\ : std_logic;
signal \N__22085\ : std_logic;
signal \N__22082\ : std_logic;
signal \N__22077\ : std_logic;
signal \N__22070\ : std_logic;
signal \N__22067\ : std_logic;
signal \N__22058\ : std_logic;
signal \N__22057\ : std_logic;
signal \N__22056\ : std_logic;
signal \N__22053\ : std_logic;
signal \N__22050\ : std_logic;
signal \N__22047\ : std_logic;
signal \N__22046\ : std_logic;
signal \N__22043\ : std_logic;
signal \N__22040\ : std_logic;
signal \N__22037\ : std_logic;
signal \N__22034\ : std_logic;
signal \N__22033\ : std_logic;
signal \N__22030\ : std_logic;
signal \N__22027\ : std_logic;
signal \N__22022\ : std_logic;
signal \N__22019\ : std_logic;
signal \N__22016\ : std_logic;
signal \N__22011\ : std_logic;
signal \N__22008\ : std_logic;
signal \N__22001\ : std_logic;
signal \N__21998\ : std_logic;
signal \N__21995\ : std_logic;
signal \N__21992\ : std_logic;
signal \N__21989\ : std_logic;
signal \N__21986\ : std_logic;
signal \N__21983\ : std_logic;
signal \N__21980\ : std_logic;
signal \N__21977\ : std_logic;
signal \N__21974\ : std_logic;
signal \N__21971\ : std_logic;
signal \N__21968\ : std_logic;
signal \N__21965\ : std_logic;
signal \N__21962\ : std_logic;
signal \N__21959\ : std_logic;
signal \N__21956\ : std_logic;
signal \N__21953\ : std_logic;
signal \N__21950\ : std_logic;
signal \N__21947\ : std_logic;
signal \N__21944\ : std_logic;
signal \N__21941\ : std_logic;
signal \N__21938\ : std_logic;
signal \N__21935\ : std_logic;
signal \N__21932\ : std_logic;
signal \N__21931\ : std_logic;
signal \N__21928\ : std_logic;
signal \N__21925\ : std_logic;
signal \N__21920\ : std_logic;
signal \N__21917\ : std_logic;
signal \N__21914\ : std_logic;
signal \N__21911\ : std_logic;
signal \N__21908\ : std_logic;
signal \N__21905\ : std_logic;
signal \N__21902\ : std_logic;
signal \N__21899\ : std_logic;
signal \N__21896\ : std_logic;
signal \N__21893\ : std_logic;
signal \N__21892\ : std_logic;
signal \N__21891\ : std_logic;
signal \N__21890\ : std_logic;
signal \N__21889\ : std_logic;
signal \N__21888\ : std_logic;
signal \N__21883\ : std_logic;
signal \N__21882\ : std_logic;
signal \N__21879\ : std_logic;
signal \N__21878\ : std_logic;
signal \N__21871\ : std_logic;
signal \N__21868\ : std_logic;
signal \N__21865\ : std_logic;
signal \N__21864\ : std_logic;
signal \N__21863\ : std_logic;
signal \N__21860\ : std_logic;
signal \N__21857\ : std_logic;
signal \N__21854\ : std_logic;
signal \N__21851\ : std_logic;
signal \N__21848\ : std_logic;
signal \N__21845\ : std_logic;
signal \N__21842\ : std_logic;
signal \N__21827\ : std_logic;
signal \N__21824\ : std_logic;
signal \N__21821\ : std_logic;
signal \N__21818\ : std_logic;
signal \N__21815\ : std_logic;
signal \N__21812\ : std_logic;
signal \N__21809\ : std_logic;
signal \N__21806\ : std_logic;
signal \N__21803\ : std_logic;
signal \N__21800\ : std_logic;
signal \N__21797\ : std_logic;
signal \N__21794\ : std_logic;
signal \N__21791\ : std_logic;
signal \N__21788\ : std_logic;
signal \N__21785\ : std_logic;
signal \N__21782\ : std_logic;
signal \N__21779\ : std_logic;
signal \N__21776\ : std_logic;
signal \N__21773\ : std_logic;
signal \N__21770\ : std_logic;
signal \N__21767\ : std_logic;
signal \N__21764\ : std_logic;
signal \N__21761\ : std_logic;
signal \N__21758\ : std_logic;
signal \N__21755\ : std_logic;
signal \N__21752\ : std_logic;
signal \N__21749\ : std_logic;
signal \N__21746\ : std_logic;
signal \N__21743\ : std_logic;
signal \N__21740\ : std_logic;
signal \N__21737\ : std_logic;
signal \N__21734\ : std_logic;
signal \N__21731\ : std_logic;
signal \N__21728\ : std_logic;
signal \N__21725\ : std_logic;
signal \N__21722\ : std_logic;
signal \N__21719\ : std_logic;
signal \N__21718\ : std_logic;
signal \N__21717\ : std_logic;
signal \N__21714\ : std_logic;
signal \N__21711\ : std_logic;
signal \N__21710\ : std_logic;
signal \N__21709\ : std_logic;
signal \N__21708\ : std_logic;
signal \N__21707\ : std_logic;
signal \N__21706\ : std_logic;
signal \N__21705\ : std_logic;
signal \N__21704\ : std_logic;
signal \N__21701\ : std_logic;
signal \N__21698\ : std_logic;
signal \N__21695\ : std_logic;
signal \N__21692\ : std_logic;
signal \N__21687\ : std_logic;
signal \N__21678\ : std_logic;
signal \N__21665\ : std_logic;
signal \N__21664\ : std_logic;
signal \N__21663\ : std_logic;
signal \N__21662\ : std_logic;
signal \N__21655\ : std_logic;
signal \N__21654\ : std_logic;
signal \N__21651\ : std_logic;
signal \N__21648\ : std_logic;
signal \N__21645\ : std_logic;
signal \N__21642\ : std_logic;
signal \N__21637\ : std_logic;
signal \N__21636\ : std_logic;
signal \N__21635\ : std_logic;
signal \N__21634\ : std_logic;
signal \N__21633\ : std_logic;
signal \N__21632\ : std_logic;
signal \N__21631\ : std_logic;
signal \N__21628\ : std_logic;
signal \N__21625\ : std_logic;
signal \N__21622\ : std_logic;
signal \N__21619\ : std_logic;
signal \N__21610\ : std_logic;
signal \N__21599\ : std_logic;
signal \N__21596\ : std_logic;
signal \N__21595\ : std_logic;
signal \N__21592\ : std_logic;
signal \N__21589\ : std_logic;
signal \N__21586\ : std_logic;
signal \N__21583\ : std_logic;
signal \N__21580\ : std_logic;
signal \N__21577\ : std_logic;
signal \N__21574\ : std_logic;
signal \N__21571\ : std_logic;
signal \N__21568\ : std_logic;
signal \N__21565\ : std_logic;
signal \N__21562\ : std_logic;
signal \N__21559\ : std_logic;
signal \N__21556\ : std_logic;
signal \N__21553\ : std_logic;
signal \N__21550\ : std_logic;
signal \N__21547\ : std_logic;
signal \N__21544\ : std_logic;
signal \N__21541\ : std_logic;
signal \N__21538\ : std_logic;
signal \N__21535\ : std_logic;
signal \N__21532\ : std_logic;
signal \N__21529\ : std_logic;
signal \N__21526\ : std_logic;
signal \N__21523\ : std_logic;
signal \N__21520\ : std_logic;
signal \N__21517\ : std_logic;
signal \N__21514\ : std_logic;
signal \N__21511\ : std_logic;
signal \N__21506\ : std_logic;
signal \N__21503\ : std_logic;
signal \N__21500\ : std_logic;
signal \N__21497\ : std_logic;
signal \N__21494\ : std_logic;
signal \N__21491\ : std_logic;
signal \N__21488\ : std_logic;
signal \N__21485\ : std_logic;
signal \N__21482\ : std_logic;
signal \N__21479\ : std_logic;
signal \N__21476\ : std_logic;
signal \N__21473\ : std_logic;
signal \N__21470\ : std_logic;
signal \N__21469\ : std_logic;
signal \N__21468\ : std_logic;
signal \N__21467\ : std_logic;
signal \N__21464\ : std_logic;
signal \N__21461\ : std_logic;
signal \N__21458\ : std_logic;
signal \N__21457\ : std_logic;
signal \N__21456\ : std_logic;
signal \N__21455\ : std_logic;
signal \N__21454\ : std_logic;
signal \N__21453\ : std_logic;
signal \N__21450\ : std_logic;
signal \N__21449\ : std_logic;
signal \N__21448\ : std_logic;
signal \N__21447\ : std_logic;
signal \N__21440\ : std_logic;
signal \N__21437\ : std_logic;
signal \N__21434\ : std_logic;
signal \N__21431\ : std_logic;
signal \N__21428\ : std_logic;
signal \N__21427\ : std_logic;
signal \N__21426\ : std_logic;
signal \N__21423\ : std_logic;
signal \N__21420\ : std_logic;
signal \N__21417\ : std_logic;
signal \N__21414\ : std_logic;
signal \N__21411\ : std_logic;
signal \N__21410\ : std_logic;
signal \N__21403\ : std_logic;
signal \N__21398\ : std_logic;
signal \N__21395\ : std_logic;
signal \N__21392\ : std_logic;
signal \N__21391\ : std_logic;
signal \N__21388\ : std_logic;
signal \N__21381\ : std_logic;
signal \N__21378\ : std_logic;
signal \N__21375\ : std_logic;
signal \N__21368\ : std_logic;
signal \N__21365\ : std_logic;
signal \N__21362\ : std_logic;
signal \N__21359\ : std_logic;
signal \N__21352\ : std_logic;
signal \N__21349\ : std_logic;
signal \N__21344\ : std_logic;
signal \N__21341\ : std_logic;
signal \N__21338\ : std_logic;
signal \N__21335\ : std_logic;
signal \N__21332\ : std_logic;
signal \N__21327\ : std_logic;
signal \N__21324\ : std_logic;
signal \N__21319\ : std_logic;
signal \N__21314\ : std_logic;
signal \N__21313\ : std_logic;
signal \N__21312\ : std_logic;
signal \N__21309\ : std_logic;
signal \N__21304\ : std_logic;
signal \N__21303\ : std_logic;
signal \N__21302\ : std_logic;
signal \N__21299\ : std_logic;
signal \N__21296\ : std_logic;
signal \N__21293\ : std_logic;
signal \N__21290\ : std_logic;
signal \N__21287\ : std_logic;
signal \N__21284\ : std_logic;
signal \N__21281\ : std_logic;
signal \N__21278\ : std_logic;
signal \N__21269\ : std_logic;
signal \N__21266\ : std_logic;
signal \N__21265\ : std_logic;
signal \N__21262\ : std_logic;
signal \N__21259\ : std_logic;
signal \N__21258\ : std_logic;
signal \N__21255\ : std_logic;
signal \N__21254\ : std_logic;
signal \N__21253\ : std_logic;
signal \N__21252\ : std_logic;
signal \N__21251\ : std_logic;
signal \N__21250\ : std_logic;
signal \N__21249\ : std_logic;
signal \N__21244\ : std_logic;
signal \N__21241\ : std_logic;
signal \N__21236\ : std_logic;
signal \N__21229\ : std_logic;
signal \N__21226\ : std_logic;
signal \N__21223\ : std_logic;
signal \N__21218\ : std_logic;
signal \N__21209\ : std_logic;
signal \N__21206\ : std_logic;
signal \N__21203\ : std_logic;
signal \N__21200\ : std_logic;
signal \N__21197\ : std_logic;
signal \N__21194\ : std_logic;
signal \N__21191\ : std_logic;
signal \N__21190\ : std_logic;
signal \N__21185\ : std_logic;
signal \N__21182\ : std_logic;
signal \N__21181\ : std_logic;
signal \N__21178\ : std_logic;
signal \N__21175\ : std_logic;
signal \N__21170\ : std_logic;
signal \N__21167\ : std_logic;
signal \N__21166\ : std_logic;
signal \N__21165\ : std_logic;
signal \N__21160\ : std_logic;
signal \N__21157\ : std_logic;
signal \N__21154\ : std_logic;
signal \N__21151\ : std_logic;
signal \N__21150\ : std_logic;
signal \N__21147\ : std_logic;
signal \N__21146\ : std_logic;
signal \N__21145\ : std_logic;
signal \N__21142\ : std_logic;
signal \N__21139\ : std_logic;
signal \N__21136\ : std_logic;
signal \N__21131\ : std_logic;
signal \N__21122\ : std_logic;
signal \N__21119\ : std_logic;
signal \N__21116\ : std_logic;
signal \N__21113\ : std_logic;
signal \N__21112\ : std_logic;
signal \N__21111\ : std_logic;
signal \N__21110\ : std_logic;
signal \N__21109\ : std_logic;
signal \N__21108\ : std_logic;
signal \N__21105\ : std_logic;
signal \N__21102\ : std_logic;
signal \N__21097\ : std_logic;
signal \N__21092\ : std_logic;
signal \N__21083\ : std_logic;
signal \N__21082\ : std_logic;
signal \N__21079\ : std_logic;
signal \N__21078\ : std_logic;
signal \N__21077\ : std_logic;
signal \N__21076\ : std_logic;
signal \N__21073\ : std_logic;
signal \N__21068\ : std_logic;
signal \N__21067\ : std_logic;
signal \N__21064\ : std_logic;
signal \N__21061\ : std_logic;
signal \N__21058\ : std_logic;
signal \N__21055\ : std_logic;
signal \N__21052\ : std_logic;
signal \N__21049\ : std_logic;
signal \N__21046\ : std_logic;
signal \N__21043\ : std_logic;
signal \N__21040\ : std_logic;
signal \N__21035\ : std_logic;
signal \N__21026\ : std_logic;
signal \N__21023\ : std_logic;
signal \N__21022\ : std_logic;
signal \N__21019\ : std_logic;
signal \N__21018\ : std_logic;
signal \N__21011\ : std_logic;
signal \N__21008\ : std_logic;
signal \N__21005\ : std_logic;
signal \N__21002\ : std_logic;
signal \N__20999\ : std_logic;
signal \N__20996\ : std_logic;
signal \N__20993\ : std_logic;
signal \N__20990\ : std_logic;
signal \N__20987\ : std_logic;
signal \N__20986\ : std_logic;
signal \N__20983\ : std_logic;
signal \N__20980\ : std_logic;
signal \N__20975\ : std_logic;
signal \N__20972\ : std_logic;
signal \N__20969\ : std_logic;
signal \N__20968\ : std_logic;
signal \N__20965\ : std_logic;
signal \N__20964\ : std_logic;
signal \N__20961\ : std_logic;
signal \N__20958\ : std_logic;
signal \N__20955\ : std_logic;
signal \N__20948\ : std_logic;
signal \N__20947\ : std_logic;
signal \N__20946\ : std_logic;
signal \N__20943\ : std_logic;
signal \N__20942\ : std_logic;
signal \N__20939\ : std_logic;
signal \N__20936\ : std_logic;
signal \N__20933\ : std_logic;
signal \N__20930\ : std_logic;
signal \N__20927\ : std_logic;
signal \N__20918\ : std_logic;
signal \N__20915\ : std_logic;
signal \N__20912\ : std_logic;
signal \N__20909\ : std_logic;
signal \N__20906\ : std_logic;
signal \N__20903\ : std_logic;
signal \N__20902\ : std_logic;
signal \N__20899\ : std_logic;
signal \N__20896\ : std_logic;
signal \N__20891\ : std_logic;
signal \N__20888\ : std_logic;
signal \N__20885\ : std_logic;
signal \N__20882\ : std_logic;
signal \N__20879\ : std_logic;
signal \N__20876\ : std_logic;
signal \N__20873\ : std_logic;
signal \N__20870\ : std_logic;
signal \N__20867\ : std_logic;
signal \N__20864\ : std_logic;
signal \N__20861\ : std_logic;
signal \N__20858\ : std_logic;
signal \N__20855\ : std_logic;
signal \N__20852\ : std_logic;
signal \N__20849\ : std_logic;
signal \N__20846\ : std_logic;
signal \N__20843\ : std_logic;
signal \N__20840\ : std_logic;
signal \N__20837\ : std_logic;
signal \N__20834\ : std_logic;
signal \N__20831\ : std_logic;
signal \N__20828\ : std_logic;
signal \N__20825\ : std_logic;
signal \N__20822\ : std_logic;
signal \N__20819\ : std_logic;
signal \N__20816\ : std_logic;
signal \N__20813\ : std_logic;
signal \N__20810\ : std_logic;
signal \N__20807\ : std_logic;
signal \N__20804\ : std_logic;
signal \N__20801\ : std_logic;
signal \N__20798\ : std_logic;
signal \N__20795\ : std_logic;
signal \N__20792\ : std_logic;
signal \N__20789\ : std_logic;
signal \N__20786\ : std_logic;
signal \N__20783\ : std_logic;
signal \N__20780\ : std_logic;
signal \N__20779\ : std_logic;
signal \N__20776\ : std_logic;
signal \N__20773\ : std_logic;
signal \N__20770\ : std_logic;
signal \N__20767\ : std_logic;
signal \N__20764\ : std_logic;
signal \N__20761\ : std_logic;
signal \N__20756\ : std_logic;
signal \N__20753\ : std_logic;
signal \N__20750\ : std_logic;
signal \N__20747\ : std_logic;
signal \N__20744\ : std_logic;
signal \N__20741\ : std_logic;
signal \N__20738\ : std_logic;
signal \N__20735\ : std_logic;
signal \N__20734\ : std_logic;
signal \N__20731\ : std_logic;
signal \N__20728\ : std_logic;
signal \N__20723\ : std_logic;
signal \N__20720\ : std_logic;
signal \N__20717\ : std_logic;
signal \N__20714\ : std_logic;
signal \N__20711\ : std_logic;
signal \N__20708\ : std_logic;
signal \N__20705\ : std_logic;
signal \N__20702\ : std_logic;
signal \N__20701\ : std_logic;
signal \N__20698\ : std_logic;
signal \N__20695\ : std_logic;
signal \N__20690\ : std_logic;
signal \N__20689\ : std_logic;
signal \N__20686\ : std_logic;
signal \N__20685\ : std_logic;
signal \N__20684\ : std_logic;
signal \N__20683\ : std_logic;
signal \N__20682\ : std_logic;
signal \N__20681\ : std_logic;
signal \N__20680\ : std_logic;
signal \N__20679\ : std_logic;
signal \N__20672\ : std_logic;
signal \N__20659\ : std_logic;
signal \N__20656\ : std_logic;
signal \N__20653\ : std_logic;
signal \N__20648\ : std_logic;
signal \N__20647\ : std_logic;
signal \N__20646\ : std_logic;
signal \N__20645\ : std_logic;
signal \N__20644\ : std_logic;
signal \N__20643\ : std_logic;
signal \N__20642\ : std_logic;
signal \N__20641\ : std_logic;
signal \N__20640\ : std_logic;
signal \N__20639\ : std_logic;
signal \N__20638\ : std_logic;
signal \N__20627\ : std_logic;
signal \N__20614\ : std_logic;
signal \N__20611\ : std_logic;
signal \N__20606\ : std_logic;
signal \N__20603\ : std_logic;
signal \N__20602\ : std_logic;
signal \N__20599\ : std_logic;
signal \N__20596\ : std_logic;
signal \N__20591\ : std_logic;
signal \N__20588\ : std_logic;
signal \N__20585\ : std_logic;
signal \N__20582\ : std_logic;
signal \N__20579\ : std_logic;
signal \N__20576\ : std_logic;
signal \N__20573\ : std_logic;
signal \N__20570\ : std_logic;
signal \N__20567\ : std_logic;
signal \N__20564\ : std_logic;
signal \N__20561\ : std_logic;
signal \N__20558\ : std_logic;
signal \N__20555\ : std_logic;
signal \N__20552\ : std_logic;
signal \N__20549\ : std_logic;
signal \N__20546\ : std_logic;
signal \N__20543\ : std_logic;
signal \N__20540\ : std_logic;
signal \N__20537\ : std_logic;
signal \N__20534\ : std_logic;
signal \N__20533\ : std_logic;
signal \N__20530\ : std_logic;
signal \N__20527\ : std_logic;
signal \N__20524\ : std_logic;
signal \N__20521\ : std_logic;
signal \N__20518\ : std_logic;
signal \N__20515\ : std_logic;
signal \N__20512\ : std_logic;
signal \N__20509\ : std_logic;
signal \N__20506\ : std_logic;
signal \N__20503\ : std_logic;
signal \N__20500\ : std_logic;
signal \N__20497\ : std_logic;
signal \N__20494\ : std_logic;
signal \N__20491\ : std_logic;
signal \N__20488\ : std_logic;
signal \N__20485\ : std_logic;
signal \N__20482\ : std_logic;
signal \N__20479\ : std_logic;
signal \N__20476\ : std_logic;
signal \N__20473\ : std_logic;
signal \N__20470\ : std_logic;
signal \N__20467\ : std_logic;
signal \N__20464\ : std_logic;
signal \N__20461\ : std_logic;
signal \N__20458\ : std_logic;
signal \N__20455\ : std_logic;
signal \N__20452\ : std_logic;
signal \N__20449\ : std_logic;
signal \N__20444\ : std_logic;
signal \N__20441\ : std_logic;
signal \N__20438\ : std_logic;
signal \N__20435\ : std_logic;
signal \N__20432\ : std_logic;
signal \N__20429\ : std_logic;
signal \N__20426\ : std_logic;
signal \N__20425\ : std_logic;
signal \N__20422\ : std_logic;
signal \N__20419\ : std_logic;
signal \N__20416\ : std_logic;
signal \N__20413\ : std_logic;
signal \N__20410\ : std_logic;
signal \N__20407\ : std_logic;
signal \N__20404\ : std_logic;
signal \N__20401\ : std_logic;
signal \N__20396\ : std_logic;
signal \N__20393\ : std_logic;
signal \N__20390\ : std_logic;
signal \N__20387\ : std_logic;
signal \N__20384\ : std_logic;
signal \N__20381\ : std_logic;
signal \N__20378\ : std_logic;
signal \N__20375\ : std_logic;
signal \N__20372\ : std_logic;
signal \N__20369\ : std_logic;
signal \N__20366\ : std_logic;
signal \N__20363\ : std_logic;
signal \N__20360\ : std_logic;
signal \N__20357\ : std_logic;
signal \N__20354\ : std_logic;
signal \N__20351\ : std_logic;
signal \N__20350\ : std_logic;
signal \N__20349\ : std_logic;
signal \N__20346\ : std_logic;
signal \N__20341\ : std_logic;
signal \N__20338\ : std_logic;
signal \N__20337\ : std_logic;
signal \N__20334\ : std_logic;
signal \N__20331\ : std_logic;
signal \N__20328\ : std_logic;
signal \N__20321\ : std_logic;
signal \N__20320\ : std_logic;
signal \N__20317\ : std_logic;
signal \N__20314\ : std_logic;
signal \N__20311\ : std_logic;
signal \N__20310\ : std_logic;
signal \N__20307\ : std_logic;
signal \N__20304\ : std_logic;
signal \N__20301\ : std_logic;
signal \N__20298\ : std_logic;
signal \N__20293\ : std_logic;
signal \N__20288\ : std_logic;
signal \N__20285\ : std_logic;
signal \N__20282\ : std_logic;
signal \N__20279\ : std_logic;
signal \N__20276\ : std_logic;
signal \N__20273\ : std_logic;
signal \N__20270\ : std_logic;
signal \N__20269\ : std_logic;
signal \N__20266\ : std_logic;
signal \N__20261\ : std_logic;
signal \N__20260\ : std_logic;
signal \N__20257\ : std_logic;
signal \N__20254\ : std_logic;
signal \N__20249\ : std_logic;
signal \N__20248\ : std_logic;
signal \N__20245\ : std_logic;
signal \N__20242\ : std_logic;
signal \N__20241\ : std_logic;
signal \N__20236\ : std_logic;
signal \N__20233\ : std_logic;
signal \N__20228\ : std_logic;
signal \N__20225\ : std_logic;
signal \N__20222\ : std_logic;
signal \N__20219\ : std_logic;
signal \N__20216\ : std_logic;
signal \N__20213\ : std_logic;
signal \N__20212\ : std_logic;
signal \N__20211\ : std_logic;
signal \N__20210\ : std_logic;
signal \N__20205\ : std_logic;
signal \N__20200\ : std_logic;
signal \N__20195\ : std_logic;
signal \N__20192\ : std_logic;
signal \N__20189\ : std_logic;
signal \N__20186\ : std_logic;
signal \N__20183\ : std_logic;
signal \N__20180\ : std_logic;
signal \N__20177\ : std_logic;
signal \N__20174\ : std_logic;
signal \N__20171\ : std_logic;
signal \N__20168\ : std_logic;
signal \N__20165\ : std_logic;
signal \N__20162\ : std_logic;
signal \N__20159\ : std_logic;
signal \N__20156\ : std_logic;
signal \N__20153\ : std_logic;
signal \N__20150\ : std_logic;
signal \N__20149\ : std_logic;
signal \N__20146\ : std_logic;
signal \N__20143\ : std_logic;
signal \N__20140\ : std_logic;
signal \N__20137\ : std_logic;
signal \N__20134\ : std_logic;
signal \N__20131\ : std_logic;
signal \N__20128\ : std_logic;
signal \N__20125\ : std_logic;
signal \N__20122\ : std_logic;
signal \N__20119\ : std_logic;
signal \N__20116\ : std_logic;
signal \N__20113\ : std_logic;
signal \N__20110\ : std_logic;
signal \N__20107\ : std_logic;
signal \N__20104\ : std_logic;
signal \N__20101\ : std_logic;
signal \N__20098\ : std_logic;
signal \N__20095\ : std_logic;
signal \N__20092\ : std_logic;
signal \N__20089\ : std_logic;
signal \N__20086\ : std_logic;
signal \N__20083\ : std_logic;
signal \N__20080\ : std_logic;
signal \N__20077\ : std_logic;
signal \N__20074\ : std_logic;
signal \N__20071\ : std_logic;
signal \N__20068\ : std_logic;
signal \N__20065\ : std_logic;
signal \N__20062\ : std_logic;
signal \N__20059\ : std_logic;
signal \N__20056\ : std_logic;
signal \N__20053\ : std_logic;
signal \N__20048\ : std_logic;
signal \N__20045\ : std_logic;
signal \N__20042\ : std_logic;
signal \N__20039\ : std_logic;
signal \N__20036\ : std_logic;
signal \N__20033\ : std_logic;
signal \N__20030\ : std_logic;
signal \N__20027\ : std_logic;
signal \N__20024\ : std_logic;
signal \N__20021\ : std_logic;
signal \N__20018\ : std_logic;
signal \N__20017\ : std_logic;
signal \N__20014\ : std_logic;
signal \N__20011\ : std_logic;
signal \N__20008\ : std_logic;
signal \N__20005\ : std_logic;
signal \N__20002\ : std_logic;
signal \N__19999\ : std_logic;
signal \N__19996\ : std_logic;
signal \N__19993\ : std_logic;
signal \N__19990\ : std_logic;
signal \N__19987\ : std_logic;
signal \N__19984\ : std_logic;
signal \N__19981\ : std_logic;
signal \N__19978\ : std_logic;
signal \N__19975\ : std_logic;
signal \N__19972\ : std_logic;
signal \N__19969\ : std_logic;
signal \N__19966\ : std_logic;
signal \N__19963\ : std_logic;
signal \N__19960\ : std_logic;
signal \N__19957\ : std_logic;
signal \N__19954\ : std_logic;
signal \N__19951\ : std_logic;
signal \N__19948\ : std_logic;
signal \N__19945\ : std_logic;
signal \N__19942\ : std_logic;
signal \N__19939\ : std_logic;
signal \N__19936\ : std_logic;
signal \N__19933\ : std_logic;
signal \N__19928\ : std_logic;
signal \N__19925\ : std_logic;
signal \N__19922\ : std_logic;
signal \N__19919\ : std_logic;
signal \N__19916\ : std_logic;
signal \N__19913\ : std_logic;
signal \N__19910\ : std_logic;
signal \N__19907\ : std_logic;
signal \N__19904\ : std_logic;
signal \N__19901\ : std_logic;
signal \N__19900\ : std_logic;
signal \N__19897\ : std_logic;
signal \N__19894\ : std_logic;
signal \N__19891\ : std_logic;
signal \N__19888\ : std_logic;
signal \N__19885\ : std_logic;
signal \N__19882\ : std_logic;
signal \N__19879\ : std_logic;
signal \N__19876\ : std_logic;
signal \N__19873\ : std_logic;
signal \N__19870\ : std_logic;
signal \N__19867\ : std_logic;
signal \N__19864\ : std_logic;
signal \N__19861\ : std_logic;
signal \N__19858\ : std_logic;
signal \N__19855\ : std_logic;
signal \N__19852\ : std_logic;
signal \N__19849\ : std_logic;
signal \N__19846\ : std_logic;
signal \N__19843\ : std_logic;
signal \N__19840\ : std_logic;
signal \N__19837\ : std_logic;
signal \N__19834\ : std_logic;
signal \N__19831\ : std_logic;
signal \N__19828\ : std_logic;
signal \N__19825\ : std_logic;
signal \N__19822\ : std_logic;
signal \N__19819\ : std_logic;
signal \N__19816\ : std_logic;
signal \N__19811\ : std_logic;
signal \N__19808\ : std_logic;
signal \N__19805\ : std_logic;
signal \N__19802\ : std_logic;
signal \N__19799\ : std_logic;
signal \N__19796\ : std_logic;
signal \N__19793\ : std_logic;
signal \N__19790\ : std_logic;
signal \N__19787\ : std_logic;
signal \N__19784\ : std_logic;
signal \N__19781\ : std_logic;
signal \N__19778\ : std_logic;
signal \N__19775\ : std_logic;
signal \N__19772\ : std_logic;
signal \N__19769\ : std_logic;
signal \N__19766\ : std_logic;
signal \N__19763\ : std_logic;
signal \N__19760\ : std_logic;
signal \N__19757\ : std_logic;
signal \N__19754\ : std_logic;
signal \N__19751\ : std_logic;
signal \N__19748\ : std_logic;
signal \N__19745\ : std_logic;
signal \N__19742\ : std_logic;
signal \N__19739\ : std_logic;
signal \N__19736\ : std_logic;
signal \N__19733\ : std_logic;
signal \N__19730\ : std_logic;
signal \N__19729\ : std_logic;
signal \N__19728\ : std_logic;
signal \N__19725\ : std_logic;
signal \N__19720\ : std_logic;
signal \N__19715\ : std_logic;
signal \N__19712\ : std_logic;
signal \N__19709\ : std_logic;
signal \N__19706\ : std_logic;
signal \N__19703\ : std_logic;
signal \N__19700\ : std_logic;
signal \N__19697\ : std_logic;
signal \N__19694\ : std_logic;
signal \N__19693\ : std_logic;
signal \N__19692\ : std_logic;
signal \N__19691\ : std_logic;
signal \N__19688\ : std_logic;
signal \N__19685\ : std_logic;
signal \N__19682\ : std_logic;
signal \N__19679\ : std_logic;
signal \N__19676\ : std_logic;
signal \N__19671\ : std_logic;
signal \N__19664\ : std_logic;
signal \N__19661\ : std_logic;
signal \N__19658\ : std_logic;
signal \N__19655\ : std_logic;
signal \N__19652\ : std_logic;
signal \N__19651\ : std_logic;
signal \N__19648\ : std_logic;
signal \N__19645\ : std_logic;
signal \N__19642\ : std_logic;
signal \N__19639\ : std_logic;
signal \N__19636\ : std_logic;
signal \N__19633\ : std_logic;
signal \N__19630\ : std_logic;
signal \N__19627\ : std_logic;
signal \N__19624\ : std_logic;
signal \N__19621\ : std_logic;
signal \N__19618\ : std_logic;
signal \N__19615\ : std_logic;
signal \N__19612\ : std_logic;
signal \N__19609\ : std_logic;
signal \N__19606\ : std_logic;
signal \N__19603\ : std_logic;
signal \N__19600\ : std_logic;
signal \N__19597\ : std_logic;
signal \N__19594\ : std_logic;
signal \N__19591\ : std_logic;
signal \N__19588\ : std_logic;
signal \N__19585\ : std_logic;
signal \N__19582\ : std_logic;
signal \N__19579\ : std_logic;
signal \N__19576\ : std_logic;
signal \N__19573\ : std_logic;
signal \N__19570\ : std_logic;
signal \N__19565\ : std_logic;
signal \N__19562\ : std_logic;
signal \N__19559\ : std_logic;
signal \N__19556\ : std_logic;
signal \N__19553\ : std_logic;
signal \N__19550\ : std_logic;
signal \N__19547\ : std_logic;
signal \N__19544\ : std_logic;
signal \N__19541\ : std_logic;
signal \N__19538\ : std_logic;
signal \N__19535\ : std_logic;
signal \N__19532\ : std_logic;
signal \N__19529\ : std_logic;
signal \N__19526\ : std_logic;
signal \N__19525\ : std_logic;
signal \N__19522\ : std_logic;
signal \N__19519\ : std_logic;
signal \N__19516\ : std_logic;
signal \N__19511\ : std_logic;
signal \N__19508\ : std_logic;
signal \N__19505\ : std_logic;
signal \N__19502\ : std_logic;
signal \N__19499\ : std_logic;
signal \N__19496\ : std_logic;
signal \N__19493\ : std_logic;
signal \N__19490\ : std_logic;
signal \N__19487\ : std_logic;
signal \N__19484\ : std_logic;
signal \N__19481\ : std_logic;
signal \N__19478\ : std_logic;
signal \N__19475\ : std_logic;
signal \N__19472\ : std_logic;
signal \N__19471\ : std_logic;
signal \N__19468\ : std_logic;
signal \N__19465\ : std_logic;
signal \N__19462\ : std_logic;
signal \N__19459\ : std_logic;
signal \N__19456\ : std_logic;
signal \N__19453\ : std_logic;
signal \N__19450\ : std_logic;
signal \N__19447\ : std_logic;
signal \N__19444\ : std_logic;
signal \N__19441\ : std_logic;
signal \N__19438\ : std_logic;
signal \N__19435\ : std_logic;
signal \N__19432\ : std_logic;
signal \N__19429\ : std_logic;
signal \N__19426\ : std_logic;
signal \N__19423\ : std_logic;
signal \N__19420\ : std_logic;
signal \N__19417\ : std_logic;
signal \N__19414\ : std_logic;
signal \N__19411\ : std_logic;
signal \N__19408\ : std_logic;
signal \N__19405\ : std_logic;
signal \N__19402\ : std_logic;
signal \N__19399\ : std_logic;
signal \N__19394\ : std_logic;
signal \N__19391\ : std_logic;
signal \N__19388\ : std_logic;
signal \N__19385\ : std_logic;
signal \N__19382\ : std_logic;
signal \N__19379\ : std_logic;
signal \N__19376\ : std_logic;
signal \N__19373\ : std_logic;
signal \N__19370\ : std_logic;
signal \N__19367\ : std_logic;
signal \N__19364\ : std_logic;
signal \N__19361\ : std_logic;
signal \N__19358\ : std_logic;
signal \N__19355\ : std_logic;
signal \N__19352\ : std_logic;
signal \N__19349\ : std_logic;
signal \N__19346\ : std_logic;
signal \N__19343\ : std_logic;
signal \N__19340\ : std_logic;
signal \N__19337\ : std_logic;
signal \N__19334\ : std_logic;
signal \N__19331\ : std_logic;
signal \N__19328\ : std_logic;
signal \N__19325\ : std_logic;
signal \N__19322\ : std_logic;
signal \N__19319\ : std_logic;
signal \N__19316\ : std_logic;
signal \N__19313\ : std_logic;
signal \N__19310\ : std_logic;
signal \N__19307\ : std_logic;
signal \N__19304\ : std_logic;
signal \N__19301\ : std_logic;
signal \N__19298\ : std_logic;
signal \N__19295\ : std_logic;
signal \N__19292\ : std_logic;
signal \N__19289\ : std_logic;
signal \N__19286\ : std_logic;
signal \N__19283\ : std_logic;
signal \N__19282\ : std_logic;
signal \N__19279\ : std_logic;
signal \N__19276\ : std_logic;
signal \N__19275\ : std_logic;
signal \N__19270\ : std_logic;
signal \N__19267\ : std_logic;
signal \N__19264\ : std_logic;
signal \N__19261\ : std_logic;
signal \N__19256\ : std_logic;
signal \N__19253\ : std_logic;
signal \N__19250\ : std_logic;
signal \N__19249\ : std_logic;
signal \N__19248\ : std_logic;
signal \N__19247\ : std_logic;
signal \N__19246\ : std_logic;
signal \N__19245\ : std_logic;
signal \N__19244\ : std_logic;
signal \N__19243\ : std_logic;
signal \N__19242\ : std_logic;
signal \N__19241\ : std_logic;
signal \N__19236\ : std_logic;
signal \N__19229\ : std_logic;
signal \N__19218\ : std_logic;
signal \N__19211\ : std_logic;
signal \N__19210\ : std_logic;
signal \N__19207\ : std_logic;
signal \N__19204\ : std_logic;
signal \N__19201\ : std_logic;
signal \N__19200\ : std_logic;
signal \N__19195\ : std_logic;
signal \N__19192\ : std_logic;
signal \N__19189\ : std_logic;
signal \N__19186\ : std_logic;
signal \N__19181\ : std_logic;
signal \N__19180\ : std_logic;
signal \N__19179\ : std_logic;
signal \N__19178\ : std_logic;
signal \N__19175\ : std_logic;
signal \N__19172\ : std_logic;
signal \N__19169\ : std_logic;
signal \N__19168\ : std_logic;
signal \N__19167\ : std_logic;
signal \N__19166\ : std_logic;
signal \N__19165\ : std_logic;
signal \N__19164\ : std_logic;
signal \N__19159\ : std_logic;
signal \N__19156\ : std_logic;
signal \N__19151\ : std_logic;
signal \N__19142\ : std_logic;
signal \N__19139\ : std_logic;
signal \N__19130\ : std_logic;
signal \N__19127\ : std_logic;
signal \N__19124\ : std_logic;
signal \N__19123\ : std_logic;
signal \N__19120\ : std_logic;
signal \N__19117\ : std_logic;
signal \N__19112\ : std_logic;
signal \N__19111\ : std_logic;
signal \N__19108\ : std_logic;
signal \N__19105\ : std_logic;
signal \N__19104\ : std_logic;
signal \N__19101\ : std_logic;
signal \N__19098\ : std_logic;
signal \N__19095\ : std_logic;
signal \N__19092\ : std_logic;
signal \N__19089\ : std_logic;
signal \N__19086\ : std_logic;
signal \N__19079\ : std_logic;
signal \N__19076\ : std_logic;
signal \N__19073\ : std_logic;
signal \N__19070\ : std_logic;
signal \N__19067\ : std_logic;
signal \N__19064\ : std_logic;
signal \N__19061\ : std_logic;
signal \N__19060\ : std_logic;
signal \N__19059\ : std_logic;
signal \N__19056\ : std_logic;
signal \N__19053\ : std_logic;
signal \N__19050\ : std_logic;
signal \N__19043\ : std_logic;
signal \N__19040\ : std_logic;
signal \N__19037\ : std_logic;
signal \N__19036\ : std_logic;
signal \N__19035\ : std_logic;
signal \N__19032\ : std_logic;
signal \N__19029\ : std_logic;
signal \N__19026\ : std_logic;
signal \N__19019\ : std_logic;
signal \N__19016\ : std_logic;
signal \N__19013\ : std_logic;
signal \N__19010\ : std_logic;
signal \N__19007\ : std_logic;
signal \N__19004\ : std_logic;
signal \N__19001\ : std_logic;
signal \N__18998\ : std_logic;
signal \N__18997\ : std_logic;
signal \N__18994\ : std_logic;
signal \N__18991\ : std_logic;
signal \N__18986\ : std_logic;
signal \N__18983\ : std_logic;
signal \N__18980\ : std_logic;
signal \N__18979\ : std_logic;
signal \N__18976\ : std_logic;
signal \N__18973\ : std_logic;
signal \N__18968\ : std_logic;
signal \N__18967\ : std_logic;
signal \N__18966\ : std_logic;
signal \N__18961\ : std_logic;
signal \N__18958\ : std_logic;
signal \N__18953\ : std_logic;
signal \N__18950\ : std_logic;
signal \N__18949\ : std_logic;
signal \N__18948\ : std_logic;
signal \N__18943\ : std_logic;
signal \N__18940\ : std_logic;
signal \N__18935\ : std_logic;
signal \N__18932\ : std_logic;
signal \N__18929\ : std_logic;
signal \N__18926\ : std_logic;
signal \N__18923\ : std_logic;
signal \N__18920\ : std_logic;
signal \N__18917\ : std_logic;
signal \N__18914\ : std_logic;
signal \N__18911\ : std_logic;
signal \N__18908\ : std_logic;
signal \N__18905\ : std_logic;
signal \N__18902\ : std_logic;
signal \N__18899\ : std_logic;
signal \N__18896\ : std_logic;
signal \N__18893\ : std_logic;
signal \N__18890\ : std_logic;
signal \N__18887\ : std_logic;
signal \N__18884\ : std_logic;
signal \N__18881\ : std_logic;
signal \N__18878\ : std_logic;
signal \N__18875\ : std_logic;
signal \N__18874\ : std_logic;
signal \N__18871\ : std_logic;
signal \N__18868\ : std_logic;
signal \N__18865\ : std_logic;
signal \N__18862\ : std_logic;
signal \N__18859\ : std_logic;
signal \N__18856\ : std_logic;
signal \N__18853\ : std_logic;
signal \N__18850\ : std_logic;
signal \N__18845\ : std_logic;
signal \N__18842\ : std_logic;
signal \N__18841\ : std_logic;
signal \N__18838\ : std_logic;
signal \N__18835\ : std_logic;
signal \N__18834\ : std_logic;
signal \N__18831\ : std_logic;
signal \N__18828\ : std_logic;
signal \N__18825\ : std_logic;
signal \N__18820\ : std_logic;
signal \N__18817\ : std_logic;
signal \N__18812\ : std_logic;
signal \N__18809\ : std_logic;
signal \N__18808\ : std_logic;
signal \N__18805\ : std_logic;
signal \N__18802\ : std_logic;
signal \N__18797\ : std_logic;
signal \N__18796\ : std_logic;
signal \N__18793\ : std_logic;
signal \N__18790\ : std_logic;
signal \N__18785\ : std_logic;
signal \N__18784\ : std_logic;
signal \N__18781\ : std_logic;
signal \N__18780\ : std_logic;
signal \N__18777\ : std_logic;
signal \N__18774\ : std_logic;
signal \N__18771\ : std_logic;
signal \N__18768\ : std_logic;
signal \N__18765\ : std_logic;
signal \N__18762\ : std_logic;
signal \N__18759\ : std_logic;
signal \N__18754\ : std_logic;
signal \N__18749\ : std_logic;
signal \N__18746\ : std_logic;
signal \N__18743\ : std_logic;
signal \N__18740\ : std_logic;
signal \N__18737\ : std_logic;
signal \N__18734\ : std_logic;
signal \N__18731\ : std_logic;
signal \N__18728\ : std_logic;
signal \N__18725\ : std_logic;
signal \N__18724\ : std_logic;
signal \N__18721\ : std_logic;
signal \N__18718\ : std_logic;
signal \N__18715\ : std_logic;
signal \N__18712\ : std_logic;
signal \N__18709\ : std_logic;
signal \N__18706\ : std_logic;
signal \N__18703\ : std_logic;
signal \N__18700\ : std_logic;
signal \N__18697\ : std_logic;
signal \N__18694\ : std_logic;
signal \N__18691\ : std_logic;
signal \N__18688\ : std_logic;
signal \N__18685\ : std_logic;
signal \N__18682\ : std_logic;
signal \N__18679\ : std_logic;
signal \N__18676\ : std_logic;
signal \N__18673\ : std_logic;
signal \N__18670\ : std_logic;
signal \N__18667\ : std_logic;
signal \N__18664\ : std_logic;
signal \N__18661\ : std_logic;
signal \N__18658\ : std_logic;
signal \N__18655\ : std_logic;
signal \N__18652\ : std_logic;
signal \N__18649\ : std_logic;
signal \N__18646\ : std_logic;
signal \N__18643\ : std_logic;
signal \N__18640\ : std_logic;
signal \N__18635\ : std_logic;
signal \N__18632\ : std_logic;
signal \N__18629\ : std_logic;
signal \N__18626\ : std_logic;
signal \N__18623\ : std_logic;
signal \N__18620\ : std_logic;
signal \N__18617\ : std_logic;
signal \N__18614\ : std_logic;
signal \N__18611\ : std_logic;
signal \N__18608\ : std_logic;
signal \N__18605\ : std_logic;
signal \N__18602\ : std_logic;
signal \N__18599\ : std_logic;
signal \N__18596\ : std_logic;
signal \N__18593\ : std_logic;
signal \N__18590\ : std_logic;
signal \N__18587\ : std_logic;
signal \N__18584\ : std_logic;
signal \N__18581\ : std_logic;
signal \N__18578\ : std_logic;
signal \N__18575\ : std_logic;
signal \N__18572\ : std_logic;
signal \N__18569\ : std_logic;
signal \N__18566\ : std_logic;
signal \N__18563\ : std_logic;
signal \N__18560\ : std_logic;
signal \N__18557\ : std_logic;
signal \N__18554\ : std_logic;
signal \N__18551\ : std_logic;
signal \N__18548\ : std_logic;
signal \N__18545\ : std_logic;
signal \N__18542\ : std_logic;
signal \N__18539\ : std_logic;
signal \N__18536\ : std_logic;
signal \N__18533\ : std_logic;
signal \N__18530\ : std_logic;
signal \N__18527\ : std_logic;
signal \N__18524\ : std_logic;
signal \N__18521\ : std_logic;
signal \N__18518\ : std_logic;
signal \N__18515\ : std_logic;
signal \N__18512\ : std_logic;
signal \N__18509\ : std_logic;
signal \N__18506\ : std_logic;
signal \N__18503\ : std_logic;
signal \N__18500\ : std_logic;
signal \N__18497\ : std_logic;
signal \N__18494\ : std_logic;
signal \N__18491\ : std_logic;
signal \N__18488\ : std_logic;
signal \N__18485\ : std_logic;
signal \N__18482\ : std_logic;
signal \N__18479\ : std_logic;
signal \N__18476\ : std_logic;
signal \N__18473\ : std_logic;
signal \N__18470\ : std_logic;
signal \N__18469\ : std_logic;
signal \N__18466\ : std_logic;
signal \N__18463\ : std_logic;
signal \N__18460\ : std_logic;
signal \N__18457\ : std_logic;
signal \N__18454\ : std_logic;
signal \N__18451\ : std_logic;
signal \N__18448\ : std_logic;
signal \N__18445\ : std_logic;
signal \N__18442\ : std_logic;
signal \N__18439\ : std_logic;
signal \N__18436\ : std_logic;
signal \N__18433\ : std_logic;
signal \N__18430\ : std_logic;
signal \N__18427\ : std_logic;
signal \N__18424\ : std_logic;
signal \N__18421\ : std_logic;
signal \N__18418\ : std_logic;
signal \N__18415\ : std_logic;
signal \N__18412\ : std_logic;
signal \N__18409\ : std_logic;
signal \N__18406\ : std_logic;
signal \N__18403\ : std_logic;
signal \N__18400\ : std_logic;
signal \N__18397\ : std_logic;
signal \N__18394\ : std_logic;
signal \N__18391\ : std_logic;
signal \N__18388\ : std_logic;
signal \N__18385\ : std_logic;
signal \N__18382\ : std_logic;
signal \N__18377\ : std_logic;
signal \N__18374\ : std_logic;
signal \N__18371\ : std_logic;
signal \N__18368\ : std_logic;
signal \N__18365\ : std_logic;
signal \N__18362\ : std_logic;
signal \N__18361\ : std_logic;
signal \N__18358\ : std_logic;
signal \N__18355\ : std_logic;
signal \N__18352\ : std_logic;
signal \N__18351\ : std_logic;
signal \N__18348\ : std_logic;
signal \N__18345\ : std_logic;
signal \N__18342\ : std_logic;
signal \N__18335\ : std_logic;
signal \N__18332\ : std_logic;
signal \N__18329\ : std_logic;
signal \N__18326\ : std_logic;
signal \N__18325\ : std_logic;
signal \N__18324\ : std_logic;
signal \N__18323\ : std_logic;
signal \N__18322\ : std_logic;
signal \N__18319\ : std_logic;
signal \N__18318\ : std_logic;
signal \N__18315\ : std_logic;
signal \N__18314\ : std_logic;
signal \N__18313\ : std_logic;
signal \N__18310\ : std_logic;
signal \N__18307\ : std_logic;
signal \N__18306\ : std_logic;
signal \N__18303\ : std_logic;
signal \N__18300\ : std_logic;
signal \N__18295\ : std_logic;
signal \N__18288\ : std_logic;
signal \N__18285\ : std_logic;
signal \N__18280\ : std_logic;
signal \N__18269\ : std_logic;
signal \N__18266\ : std_logic;
signal \N__18263\ : std_logic;
signal \N__18262\ : std_logic;
signal \N__18261\ : std_logic;
signal \N__18260\ : std_logic;
signal \N__18259\ : std_logic;
signal \N__18258\ : std_logic;
signal \N__18257\ : std_logic;
signal \N__18256\ : std_logic;
signal \N__18255\ : std_logic;
signal \N__18254\ : std_logic;
signal \N__18253\ : std_logic;
signal \N__18250\ : std_logic;
signal \N__18247\ : std_logic;
signal \N__18242\ : std_logic;
signal \N__18227\ : std_logic;
signal \N__18218\ : std_logic;
signal \N__18215\ : std_logic;
signal \N__18212\ : std_logic;
signal \N__18209\ : std_logic;
signal \N__18208\ : std_logic;
signal \N__18205\ : std_logic;
signal \N__18204\ : std_logic;
signal \N__18203\ : std_logic;
signal \N__18200\ : std_logic;
signal \N__18197\ : std_logic;
signal \N__18194\ : std_logic;
signal \N__18191\ : std_logic;
signal \N__18188\ : std_logic;
signal \N__18183\ : std_logic;
signal \N__18180\ : std_logic;
signal \N__18177\ : std_logic;
signal \N__18174\ : std_logic;
signal \N__18167\ : std_logic;
signal \N__18166\ : std_logic;
signal \N__18161\ : std_logic;
signal \N__18158\ : std_logic;
signal \N__18155\ : std_logic;
signal \N__18152\ : std_logic;
signal \N__18149\ : std_logic;
signal \N__18146\ : std_logic;
signal \N__18143\ : std_logic;
signal \N__18140\ : std_logic;
signal \N__18139\ : std_logic;
signal \N__18134\ : std_logic;
signal \N__18131\ : std_logic;
signal \N__18128\ : std_logic;
signal \N__18125\ : std_logic;
signal \N__18122\ : std_logic;
signal \N__18119\ : std_logic;
signal \N__18116\ : std_logic;
signal \N__18113\ : std_logic;
signal \N__18112\ : std_logic;
signal \N__18109\ : std_logic;
signal \N__18106\ : std_logic;
signal \N__18103\ : std_logic;
signal \N__18100\ : std_logic;
signal \N__18097\ : std_logic;
signal \N__18094\ : std_logic;
signal \N__18089\ : std_logic;
signal \N__18086\ : std_logic;
signal \N__18083\ : std_logic;
signal \N__18080\ : std_logic;
signal \N__18077\ : std_logic;
signal \N__18074\ : std_logic;
signal \N__18071\ : std_logic;
signal \N__18068\ : std_logic;
signal \N__18065\ : std_logic;
signal \N__18062\ : std_logic;
signal \N__18059\ : std_logic;
signal \N__18056\ : std_logic;
signal \N__18053\ : std_logic;
signal \N__18050\ : std_logic;
signal \N__18047\ : std_logic;
signal \N__18044\ : std_logic;
signal \N__18041\ : std_logic;
signal \N__18038\ : std_logic;
signal \N__18035\ : std_logic;
signal \N__18032\ : std_logic;
signal \N__18029\ : std_logic;
signal \N__18026\ : std_logic;
signal \N__18023\ : std_logic;
signal \N__18020\ : std_logic;
signal \N__18017\ : std_logic;
signal \N__18014\ : std_logic;
signal \N__18013\ : std_logic;
signal \N__18010\ : std_logic;
signal \N__18007\ : std_logic;
signal \N__18002\ : std_logic;
signal \N__17999\ : std_logic;
signal \N__17998\ : std_logic;
signal \N__17995\ : std_logic;
signal \N__17992\ : std_logic;
signal \N__17987\ : std_logic;
signal \N__17986\ : std_logic;
signal \N__17983\ : std_logic;
signal \N__17980\ : std_logic;
signal \N__17977\ : std_logic;
signal \N__17974\ : std_logic;
signal \N__17971\ : std_logic;
signal \N__17966\ : std_logic;
signal \N__17963\ : std_logic;
signal \N__17960\ : std_logic;
signal \N__17957\ : std_logic;
signal \N__17954\ : std_logic;
signal \N__17951\ : std_logic;
signal \N__17948\ : std_logic;
signal \N__17945\ : std_logic;
signal \N__17942\ : std_logic;
signal \N__17939\ : std_logic;
signal \N__17936\ : std_logic;
signal \N__17933\ : std_logic;
signal \N__17930\ : std_logic;
signal \N__17927\ : std_logic;
signal \N__17924\ : std_logic;
signal \N__17921\ : std_logic;
signal \N__17920\ : std_logic;
signal \N__17917\ : std_logic;
signal \N__17914\ : std_logic;
signal \N__17911\ : std_logic;
signal \N__17906\ : std_logic;
signal \N__17903\ : std_logic;
signal \N__17900\ : std_logic;
signal \N__17897\ : std_logic;
signal \N__17894\ : std_logic;
signal \N__17891\ : std_logic;
signal \N__17888\ : std_logic;
signal \N__17885\ : std_logic;
signal \N__17882\ : std_logic;
signal \N__17879\ : std_logic;
signal \N__17876\ : std_logic;
signal \N__17873\ : std_logic;
signal \N__17870\ : std_logic;
signal \N__17867\ : std_logic;
signal \N__17864\ : std_logic;
signal \N__17861\ : std_logic;
signal \N__17858\ : std_logic;
signal \N__17857\ : std_logic;
signal \N__17854\ : std_logic;
signal \N__17851\ : std_logic;
signal \N__17848\ : std_logic;
signal \N__17843\ : std_logic;
signal \N__17840\ : std_logic;
signal \N__17837\ : std_logic;
signal \N__17834\ : std_logic;
signal \N__17831\ : std_logic;
signal \N__17828\ : std_logic;
signal \N__17825\ : std_logic;
signal \N__17822\ : std_logic;
signal \N__17821\ : std_logic;
signal \N__17818\ : std_logic;
signal \N__17815\ : std_logic;
signal \N__17812\ : std_logic;
signal \N__17809\ : std_logic;
signal \N__17806\ : std_logic;
signal \N__17803\ : std_logic;
signal \N__17798\ : std_logic;
signal \N__17795\ : std_logic;
signal \N__17792\ : std_logic;
signal \N__17789\ : std_logic;
signal \N__17786\ : std_logic;
signal \N__17783\ : std_logic;
signal \N__17782\ : std_logic;
signal \N__17779\ : std_logic;
signal \N__17776\ : std_logic;
signal \N__17773\ : std_logic;
signal \N__17770\ : std_logic;
signal \N__17765\ : std_logic;
signal \N__17764\ : std_logic;
signal \N__17761\ : std_logic;
signal \N__17758\ : std_logic;
signal \N__17755\ : std_logic;
signal \N__17752\ : std_logic;
signal \N__17749\ : std_logic;
signal \N__17746\ : std_logic;
signal \N__17743\ : std_logic;
signal \N__17738\ : std_logic;
signal \N__17735\ : std_logic;
signal \N__17732\ : std_logic;
signal \N__17731\ : std_logic;
signal \N__17730\ : std_logic;
signal \N__17729\ : std_logic;
signal \N__17728\ : std_logic;
signal \N__17727\ : std_logic;
signal \N__17724\ : std_logic;
signal \N__17723\ : std_logic;
signal \N__17722\ : std_logic;
signal \N__17715\ : std_logic;
signal \N__17714\ : std_logic;
signal \N__17713\ : std_logic;
signal \N__17710\ : std_logic;
signal \N__17709\ : std_logic;
signal \N__17706\ : std_logic;
signal \N__17705\ : std_logic;
signal \N__17702\ : std_logic;
signal \N__17699\ : std_logic;
signal \N__17696\ : std_logic;
signal \N__17695\ : std_logic;
signal \N__17692\ : std_logic;
signal \N__17689\ : std_logic;
signal \N__17686\ : std_logic;
signal \N__17685\ : std_logic;
signal \N__17682\ : std_logic;
signal \N__17677\ : std_logic;
signal \N__17674\ : std_logic;
signal \N__17671\ : std_logic;
signal \N__17668\ : std_logic;
signal \N__17665\ : std_logic;
signal \N__17662\ : std_logic;
signal \N__17659\ : std_logic;
signal \N__17656\ : std_logic;
signal \N__17653\ : std_logic;
signal \N__17650\ : std_logic;
signal \N__17645\ : std_logic;
signal \N__17636\ : std_logic;
signal \N__17621\ : std_logic;
signal \N__17620\ : std_logic;
signal \N__17617\ : std_logic;
signal \N__17614\ : std_logic;
signal \N__17613\ : std_logic;
signal \N__17612\ : std_logic;
signal \N__17611\ : std_logic;
signal \N__17610\ : std_logic;
signal \N__17605\ : std_logic;
signal \N__17602\ : std_logic;
signal \N__17599\ : std_logic;
signal \N__17598\ : std_logic;
signal \N__17595\ : std_logic;
signal \N__17594\ : std_logic;
signal \N__17593\ : std_logic;
signal \N__17592\ : std_logic;
signal \N__17589\ : std_logic;
signal \N__17584\ : std_logic;
signal \N__17581\ : std_logic;
signal \N__17578\ : std_logic;
signal \N__17575\ : std_logic;
signal \N__17572\ : std_logic;
signal \N__17569\ : std_logic;
signal \N__17566\ : std_logic;
signal \N__17565\ : std_logic;
signal \N__17562\ : std_logic;
signal \N__17559\ : std_logic;
signal \N__17552\ : std_logic;
signal \N__17549\ : std_logic;
signal \N__17544\ : std_logic;
signal \N__17541\ : std_logic;
signal \N__17538\ : std_logic;
signal \N__17525\ : std_logic;
signal \N__17524\ : std_logic;
signal \N__17521\ : std_logic;
signal \N__17518\ : std_logic;
signal \N__17513\ : std_logic;
signal \N__17510\ : std_logic;
signal \N__17509\ : std_logic;
signal \N__17506\ : std_logic;
signal \N__17503\ : std_logic;
signal \N__17502\ : std_logic;
signal \N__17501\ : std_logic;
signal \N__17500\ : std_logic;
signal \N__17497\ : std_logic;
signal \N__17494\ : std_logic;
signal \N__17491\ : std_logic;
signal \N__17490\ : std_logic;
signal \N__17485\ : std_logic;
signal \N__17484\ : std_logic;
signal \N__17483\ : std_logic;
signal \N__17476\ : std_logic;
signal \N__17473\ : std_logic;
signal \N__17470\ : std_logic;
signal \N__17467\ : std_logic;
signal \N__17464\ : std_logic;
signal \N__17461\ : std_logic;
signal \N__17456\ : std_logic;
signal \N__17447\ : std_logic;
signal \N__17446\ : std_logic;
signal \N__17445\ : std_logic;
signal \N__17444\ : std_logic;
signal \N__17441\ : std_logic;
signal \N__17438\ : std_logic;
signal \N__17437\ : std_logic;
signal \N__17436\ : std_logic;
signal \N__17433\ : std_logic;
signal \N__17432\ : std_logic;
signal \N__17431\ : std_logic;
signal \N__17428\ : std_logic;
signal \N__17423\ : std_logic;
signal \N__17420\ : std_logic;
signal \N__17417\ : std_logic;
signal \N__17414\ : std_logic;
signal \N__17411\ : std_logic;
signal \N__17408\ : std_logic;
signal \N__17405\ : std_logic;
signal \N__17402\ : std_logic;
signal \N__17397\ : std_logic;
signal \N__17394\ : std_logic;
signal \N__17381\ : std_logic;
signal \N__17380\ : std_logic;
signal \N__17377\ : std_logic;
signal \N__17376\ : std_logic;
signal \N__17373\ : std_logic;
signal \N__17370\ : std_logic;
signal \N__17365\ : std_logic;
signal \N__17360\ : std_logic;
signal \N__17357\ : std_logic;
signal \N__17354\ : std_logic;
signal \N__17351\ : std_logic;
signal \N__17348\ : std_logic;
signal \N__17345\ : std_logic;
signal \N__17342\ : std_logic;
signal \N__17339\ : std_logic;
signal \N__17336\ : std_logic;
signal \N__17333\ : std_logic;
signal \N__17330\ : std_logic;
signal \N__17327\ : std_logic;
signal \N__17324\ : std_logic;
signal \N__17321\ : std_logic;
signal \N__17318\ : std_logic;
signal \N__17315\ : std_logic;
signal \N__17314\ : std_logic;
signal \N__17311\ : std_logic;
signal \N__17308\ : std_logic;
signal \N__17303\ : std_logic;
signal \N__17302\ : std_logic;
signal \N__17301\ : std_logic;
signal \N__17300\ : std_logic;
signal \N__17299\ : std_logic;
signal \N__17294\ : std_logic;
signal \N__17291\ : std_logic;
signal \N__17290\ : std_logic;
signal \N__17289\ : std_logic;
signal \N__17286\ : std_logic;
signal \N__17285\ : std_logic;
signal \N__17282\ : std_logic;
signal \N__17279\ : std_logic;
signal \N__17276\ : std_logic;
signal \N__17273\ : std_logic;
signal \N__17270\ : std_logic;
signal \N__17267\ : std_logic;
signal \N__17264\ : std_logic;
signal \N__17261\ : std_logic;
signal \N__17254\ : std_logic;
signal \N__17247\ : std_logic;
signal \N__17242\ : std_logic;
signal \N__17239\ : std_logic;
signal \N__17234\ : std_logic;
signal \N__17231\ : std_logic;
signal \N__17228\ : std_logic;
signal \N__17225\ : std_logic;
signal \N__17222\ : std_logic;
signal \N__17221\ : std_logic;
signal \N__17218\ : std_logic;
signal \N__17217\ : std_logic;
signal \N__17214\ : std_logic;
signal \N__17209\ : std_logic;
signal \N__17206\ : std_logic;
signal \N__17201\ : std_logic;
signal \N__17198\ : std_logic;
signal \N__17195\ : std_logic;
signal \N__17192\ : std_logic;
signal \N__17189\ : std_logic;
signal \N__17186\ : std_logic;
signal \N__17185\ : std_logic;
signal \N__17182\ : std_logic;
signal \N__17179\ : std_logic;
signal \N__17176\ : std_logic;
signal \N__17173\ : std_logic;
signal \N__17170\ : std_logic;
signal \N__17167\ : std_logic;
signal \N__17164\ : std_logic;
signal \N__17161\ : std_logic;
signal \N__17156\ : std_logic;
signal \N__17153\ : std_logic;
signal \N__17150\ : std_logic;
signal \N__17149\ : std_logic;
signal \N__17146\ : std_logic;
signal \N__17143\ : std_logic;
signal \N__17140\ : std_logic;
signal \N__17137\ : std_logic;
signal \N__17134\ : std_logic;
signal \N__17131\ : std_logic;
signal \N__17128\ : std_logic;
signal \N__17125\ : std_logic;
signal \N__17120\ : std_logic;
signal \N__17117\ : std_logic;
signal \N__17114\ : std_logic;
signal \N__17111\ : std_logic;
signal \N__17108\ : std_logic;
signal \N__17105\ : std_logic;
signal \N__17104\ : std_logic;
signal \N__17101\ : std_logic;
signal \N__17098\ : std_logic;
signal \N__17095\ : std_logic;
signal \N__17092\ : std_logic;
signal \N__17087\ : std_logic;
signal \N__17084\ : std_logic;
signal \N__17081\ : std_logic;
signal \N__17078\ : std_logic;
signal \N__17075\ : std_logic;
signal \N__17072\ : std_logic;
signal \N__17069\ : std_logic;
signal \N__17066\ : std_logic;
signal \N__17063\ : std_logic;
signal \N__17060\ : std_logic;
signal \N__17057\ : std_logic;
signal \N__17056\ : std_logic;
signal \N__17055\ : std_logic;
signal \N__17054\ : std_logic;
signal \N__17049\ : std_logic;
signal \N__17048\ : std_logic;
signal \N__17047\ : std_logic;
signal \N__17046\ : std_logic;
signal \N__17043\ : std_logic;
signal \N__17042\ : std_logic;
signal \N__17041\ : std_logic;
signal \N__17038\ : std_logic;
signal \N__17035\ : std_logic;
signal \N__17028\ : std_logic;
signal \N__17021\ : std_logic;
signal \N__17012\ : std_logic;
signal \N__17011\ : std_logic;
signal \N__17010\ : std_logic;
signal \N__17009\ : std_logic;
signal \N__17006\ : std_logic;
signal \N__17001\ : std_logic;
signal \N__17000\ : std_logic;
signal \N__16999\ : std_logic;
signal \N__16998\ : std_logic;
signal \N__16997\ : std_logic;
signal \N__16996\ : std_logic;
signal \N__16995\ : std_logic;
signal \N__16992\ : std_logic;
signal \N__16987\ : std_logic;
signal \N__16982\ : std_logic;
signal \N__16973\ : std_logic;
signal \N__16964\ : std_logic;
signal \N__16961\ : std_logic;
signal \N__16958\ : std_logic;
signal \N__16955\ : std_logic;
signal \N__16952\ : std_logic;
signal \N__16949\ : std_logic;
signal \N__16946\ : std_logic;
signal \N__16943\ : std_logic;
signal \N__16940\ : std_logic;
signal \N__16937\ : std_logic;
signal \N__16934\ : std_logic;
signal \N__16931\ : std_logic;
signal \N__16928\ : std_logic;
signal \N__16925\ : std_logic;
signal \N__16922\ : std_logic;
signal \N__16919\ : std_logic;
signal \N__16916\ : std_logic;
signal \N__16913\ : std_logic;
signal \N__16910\ : std_logic;
signal \N__16907\ : std_logic;
signal \N__16906\ : std_logic;
signal \N__16905\ : std_logic;
signal \N__16904\ : std_logic;
signal \N__16903\ : std_logic;
signal \N__16902\ : std_logic;
signal \N__16901\ : std_logic;
signal \N__16898\ : std_logic;
signal \N__16893\ : std_logic;
signal \N__16890\ : std_logic;
signal \N__16887\ : std_logic;
signal \N__16882\ : std_logic;
signal \N__16879\ : std_logic;
signal \N__16876\ : std_logic;
signal \N__16865\ : std_logic;
signal \N__16862\ : std_logic;
signal \N__16859\ : std_logic;
signal \N__16856\ : std_logic;
signal \N__16853\ : std_logic;
signal \N__16852\ : std_logic;
signal \N__16849\ : std_logic;
signal \N__16848\ : std_logic;
signal \N__16847\ : std_logic;
signal \N__16844\ : std_logic;
signal \N__16843\ : std_logic;
signal \N__16842\ : std_logic;
signal \N__16839\ : std_logic;
signal \N__16836\ : std_logic;
signal \N__16833\ : std_logic;
signal \N__16828\ : std_logic;
signal \N__16825\ : std_logic;
signal \N__16824\ : std_logic;
signal \N__16823\ : std_logic;
signal \N__16822\ : std_logic;
signal \N__16821\ : std_logic;
signal \N__16816\ : std_logic;
signal \N__16813\ : std_logic;
signal \N__16810\ : std_logic;
signal \N__16807\ : std_logic;
signal \N__16800\ : std_logic;
signal \N__16797\ : std_logic;
signal \N__16794\ : std_logic;
signal \N__16789\ : std_logic;
signal \N__16784\ : std_logic;
signal \N__16775\ : std_logic;
signal \N__16772\ : std_logic;
signal \N__16769\ : std_logic;
signal \N__16766\ : std_logic;
signal \N__16763\ : std_logic;
signal \N__16760\ : std_logic;
signal \N__16757\ : std_logic;
signal \N__16756\ : std_logic;
signal \N__16753\ : std_logic;
signal \N__16752\ : std_logic;
signal \N__16749\ : std_logic;
signal \N__16748\ : std_logic;
signal \N__16747\ : std_logic;
signal \N__16746\ : std_logic;
signal \N__16745\ : std_logic;
signal \N__16744\ : std_logic;
signal \N__16741\ : std_logic;
signal \N__16738\ : std_logic;
signal \N__16735\ : std_logic;
signal \N__16728\ : std_logic;
signal \N__16727\ : std_logic;
signal \N__16724\ : std_logic;
signal \N__16721\ : std_logic;
signal \N__16716\ : std_logic;
signal \N__16711\ : std_logic;
signal \N__16708\ : std_logic;
signal \N__16703\ : std_logic;
signal \N__16700\ : std_logic;
signal \N__16697\ : std_logic;
signal \N__16688\ : std_logic;
signal \N__16685\ : std_logic;
signal \N__16682\ : std_logic;
signal \N__16679\ : std_logic;
signal \N__16676\ : std_logic;
signal \N__16673\ : std_logic;
signal \N__16670\ : std_logic;
signal \N__16667\ : std_logic;
signal \N__16664\ : std_logic;
signal \N__16661\ : std_logic;
signal \N__16658\ : std_logic;
signal \N__16655\ : std_logic;
signal \N__16652\ : std_logic;
signal \N__16649\ : std_logic;
signal \N__16646\ : std_logic;
signal \N__16643\ : std_logic;
signal \N__16640\ : std_logic;
signal \N__16639\ : std_logic;
signal \N__16638\ : std_logic;
signal \N__16633\ : std_logic;
signal \N__16632\ : std_logic;
signal \N__16631\ : std_logic;
signal \N__16630\ : std_logic;
signal \N__16629\ : std_logic;
signal \N__16628\ : std_logic;
signal \N__16627\ : std_logic;
signal \N__16624\ : std_logic;
signal \N__16621\ : std_logic;
signal \N__16618\ : std_logic;
signal \N__16615\ : std_logic;
signal \N__16612\ : std_logic;
signal \N__16609\ : std_logic;
signal \N__16606\ : std_logic;
signal \N__16603\ : std_logic;
signal \N__16596\ : std_logic;
signal \N__16583\ : std_logic;
signal \N__16580\ : std_logic;
signal \N__16577\ : std_logic;
signal \N__16574\ : std_logic;
signal \N__16571\ : std_logic;
signal \N__16568\ : std_logic;
signal \N__16565\ : std_logic;
signal \N__16562\ : std_logic;
signal \N__16559\ : std_logic;
signal \N__16556\ : std_logic;
signal \N__16553\ : std_logic;
signal \N__16550\ : std_logic;
signal \N__16547\ : std_logic;
signal \N__16544\ : std_logic;
signal \N__16541\ : std_logic;
signal \N__16540\ : std_logic;
signal \N__16537\ : std_logic;
signal \N__16536\ : std_logic;
signal \N__16533\ : std_logic;
signal \N__16530\ : std_logic;
signal \N__16527\ : std_logic;
signal \N__16524\ : std_logic;
signal \N__16517\ : std_logic;
signal \N__16514\ : std_logic;
signal \N__16511\ : std_logic;
signal \N__16508\ : std_logic;
signal \N__16505\ : std_logic;
signal \N__16502\ : std_logic;
signal \N__16501\ : std_logic;
signal \N__16500\ : std_logic;
signal \N__16499\ : std_logic;
signal \N__16498\ : std_logic;
signal \N__16495\ : std_logic;
signal \N__16494\ : std_logic;
signal \N__16491\ : std_logic;
signal \N__16488\ : std_logic;
signal \N__16485\ : std_logic;
signal \N__16482\ : std_logic;
signal \N__16479\ : std_logic;
signal \N__16476\ : std_logic;
signal \N__16475\ : std_logic;
signal \N__16474\ : std_logic;
signal \N__16473\ : std_logic;
signal \N__16470\ : std_logic;
signal \N__16465\ : std_logic;
signal \N__16458\ : std_logic;
signal \N__16453\ : std_logic;
signal \N__16450\ : std_logic;
signal \N__16447\ : std_logic;
signal \N__16442\ : std_logic;
signal \N__16439\ : std_logic;
signal \N__16430\ : std_logic;
signal \N__16429\ : std_logic;
signal \N__16426\ : std_logic;
signal \N__16425\ : std_logic;
signal \N__16424\ : std_logic;
signal \N__16423\ : std_logic;
signal \N__16420\ : std_logic;
signal \N__16417\ : std_logic;
signal \N__16414\ : std_logic;
signal \N__16411\ : std_logic;
signal \N__16410\ : std_logic;
signal \N__16409\ : std_logic;
signal \N__16408\ : std_logic;
signal \N__16407\ : std_logic;
signal \N__16404\ : std_logic;
signal \N__16399\ : std_logic;
signal \N__16394\ : std_logic;
signal \N__16387\ : std_logic;
signal \N__16384\ : std_logic;
signal \N__16379\ : std_logic;
signal \N__16376\ : std_logic;
signal \N__16373\ : std_logic;
signal \N__16364\ : std_logic;
signal \N__16363\ : std_logic;
signal \N__16362\ : std_logic;
signal \N__16359\ : std_logic;
signal \N__16358\ : std_logic;
signal \N__16355\ : std_logic;
signal \N__16354\ : std_logic;
signal \N__16351\ : std_logic;
signal \N__16350\ : std_logic;
signal \N__16347\ : std_logic;
signal \N__16344\ : std_logic;
signal \N__16341\ : std_logic;
signal \N__16340\ : std_logic;
signal \N__16339\ : std_logic;
signal \N__16338\ : std_logic;
signal \N__16335\ : std_logic;
signal \N__16332\ : std_logic;
signal \N__16329\ : std_logic;
signal \N__16326\ : std_logic;
signal \N__16323\ : std_logic;
signal \N__16320\ : std_logic;
signal \N__16313\ : std_logic;
signal \N__16306\ : std_logic;
signal \N__16301\ : std_logic;
signal \N__16296\ : std_logic;
signal \N__16289\ : std_logic;
signal \N__16286\ : std_logic;
signal \N__16283\ : std_logic;
signal \N__16280\ : std_logic;
signal \N__16277\ : std_logic;
signal \N__16274\ : std_logic;
signal \N__16271\ : std_logic;
signal \N__16268\ : std_logic;
signal \N__16267\ : std_logic;
signal \N__16266\ : std_logic;
signal \N__16263\ : std_logic;
signal \N__16260\ : std_logic;
signal \N__16257\ : std_logic;
signal \N__16250\ : std_logic;
signal \N__16247\ : std_logic;
signal \N__16246\ : std_logic;
signal \N__16245\ : std_logic;
signal \N__16242\ : std_logic;
signal \N__16239\ : std_logic;
signal \N__16236\ : std_logic;
signal \N__16233\ : std_logic;
signal \N__16230\ : std_logic;
signal \N__16225\ : std_logic;
signal \N__16220\ : std_logic;
signal \N__16217\ : std_logic;
signal \N__16216\ : std_logic;
signal \N__16215\ : std_logic;
signal \N__16212\ : std_logic;
signal \N__16209\ : std_logic;
signal \N__16206\ : std_logic;
signal \N__16203\ : std_logic;
signal \N__16200\ : std_logic;
signal \N__16193\ : std_logic;
signal \N__16190\ : std_logic;
signal \N__16187\ : std_logic;
signal \N__16184\ : std_logic;
signal \N__16181\ : std_logic;
signal \N__16178\ : std_logic;
signal \N__16175\ : std_logic;
signal \N__16172\ : std_logic;
signal \N__16169\ : std_logic;
signal \N__16166\ : std_logic;
signal \N__16163\ : std_logic;
signal \N__16160\ : std_logic;
signal \N__16159\ : std_logic;
signal \N__16156\ : std_logic;
signal \N__16151\ : std_logic;
signal \N__16150\ : std_logic;
signal \N__16147\ : std_logic;
signal \N__16144\ : std_logic;
signal \N__16139\ : std_logic;
signal \N__16136\ : std_logic;
signal \N__16133\ : std_logic;
signal \N__16130\ : std_logic;
signal \N__16127\ : std_logic;
signal \N__16124\ : std_logic;
signal \N__16121\ : std_logic;
signal \N__16118\ : std_logic;
signal \N__16115\ : std_logic;
signal \N__16112\ : std_logic;
signal \N__16109\ : std_logic;
signal \N__16106\ : std_logic;
signal \N__16103\ : std_logic;
signal \N__16100\ : std_logic;
signal \N__16097\ : std_logic;
signal \N__16094\ : std_logic;
signal \N__16091\ : std_logic;
signal \N__16088\ : std_logic;
signal \N__16085\ : std_logic;
signal \N__16082\ : std_logic;
signal \N__16079\ : std_logic;
signal \N__16076\ : std_logic;
signal \N__16073\ : std_logic;
signal \N__16072\ : std_logic;
signal \N__16071\ : std_logic;
signal \N__16068\ : std_logic;
signal \N__16065\ : std_logic;
signal \N__16062\ : std_logic;
signal \N__16059\ : std_logic;
signal \N__16056\ : std_logic;
signal \N__16049\ : std_logic;
signal \N__16046\ : std_logic;
signal \N__16043\ : std_logic;
signal \N__16040\ : std_logic;
signal \N__16037\ : std_logic;
signal \N__16034\ : std_logic;
signal \N__16031\ : std_logic;
signal \N__16028\ : std_logic;
signal \N__16025\ : std_logic;
signal \N__16022\ : std_logic;
signal \N__16019\ : std_logic;
signal \N__16016\ : std_logic;
signal \N__16015\ : std_logic;
signal \N__16012\ : std_logic;
signal \N__16009\ : std_logic;
signal \N__16004\ : std_logic;
signal \N__16003\ : std_logic;
signal \N__16002\ : std_logic;
signal \N__15999\ : std_logic;
signal \N__15994\ : std_logic;
signal \N__15989\ : std_logic;
signal \N__15986\ : std_logic;
signal \N__15983\ : std_logic;
signal \N__15980\ : std_logic;
signal \N__15977\ : std_logic;
signal \N__15976\ : std_logic;
signal \N__15973\ : std_logic;
signal \N__15970\ : std_logic;
signal \N__15967\ : std_logic;
signal \N__15964\ : std_logic;
signal \N__15961\ : std_logic;
signal \N__15958\ : std_logic;
signal \N__15955\ : std_logic;
signal \N__15952\ : std_logic;
signal \N__15949\ : std_logic;
signal \N__15946\ : std_logic;
signal \N__15943\ : std_logic;
signal \N__15940\ : std_logic;
signal \N__15937\ : std_logic;
signal \N__15934\ : std_logic;
signal \N__15931\ : std_logic;
signal \N__15928\ : std_logic;
signal \N__15925\ : std_logic;
signal \N__15922\ : std_logic;
signal \N__15919\ : std_logic;
signal \N__15916\ : std_logic;
signal \N__15913\ : std_logic;
signal \N__15910\ : std_logic;
signal \N__15907\ : std_logic;
signal \N__15904\ : std_logic;
signal \N__15901\ : std_logic;
signal \N__15898\ : std_logic;
signal \N__15895\ : std_logic;
signal \N__15892\ : std_logic;
signal \N__15887\ : std_logic;
signal \N__15884\ : std_logic;
signal \N__15881\ : std_logic;
signal \N__15878\ : std_logic;
signal \N__15877\ : std_logic;
signal \N__15876\ : std_logic;
signal \N__15875\ : std_logic;
signal \N__15872\ : std_logic;
signal \N__15869\ : std_logic;
signal \N__15866\ : std_logic;
signal \N__15863\ : std_logic;
signal \N__15860\ : std_logic;
signal \N__15859\ : std_logic;
signal \N__15854\ : std_logic;
signal \N__15849\ : std_logic;
signal \N__15848\ : std_logic;
signal \N__15845\ : std_logic;
signal \N__15842\ : std_logic;
signal \N__15839\ : std_logic;
signal \N__15834\ : std_logic;
signal \N__15827\ : std_logic;
signal \N__15826\ : std_logic;
signal \N__15825\ : std_logic;
signal \N__15824\ : std_logic;
signal \N__15821\ : std_logic;
signal \N__15818\ : std_logic;
signal \N__15813\ : std_logic;
signal \N__15808\ : std_logic;
signal \N__15807\ : std_logic;
signal \N__15802\ : std_logic;
signal \N__15801\ : std_logic;
signal \N__15798\ : std_logic;
signal \N__15795\ : std_logic;
signal \N__15792\ : std_logic;
signal \N__15789\ : std_logic;
signal \N__15782\ : std_logic;
signal \N__15779\ : std_logic;
signal \N__15778\ : std_logic;
signal \N__15775\ : std_logic;
signal \N__15774\ : std_logic;
signal \N__15773\ : std_logic;
signal \N__15770\ : std_logic;
signal \N__15767\ : std_logic;
signal \N__15764\ : std_logic;
signal \N__15761\ : std_logic;
signal \N__15758\ : std_logic;
signal \N__15755\ : std_logic;
signal \N__15752\ : std_logic;
signal \N__15749\ : std_logic;
signal \N__15744\ : std_logic;
signal \N__15741\ : std_logic;
signal \N__15734\ : std_logic;
signal \N__15731\ : std_logic;
signal \N__15730\ : std_logic;
signal \N__15729\ : std_logic;
signal \N__15726\ : std_logic;
signal \N__15725\ : std_logic;
signal \N__15722\ : std_logic;
signal \N__15719\ : std_logic;
signal \N__15716\ : std_logic;
signal \N__15713\ : std_logic;
signal \N__15710\ : std_logic;
signal \N__15707\ : std_logic;
signal \N__15704\ : std_logic;
signal \N__15699\ : std_logic;
signal \N__15696\ : std_logic;
signal \N__15693\ : std_logic;
signal \N__15690\ : std_logic;
signal \N__15683\ : std_logic;
signal \N__15682\ : std_logic;
signal \N__15681\ : std_logic;
signal \N__15678\ : std_logic;
signal \N__15675\ : std_logic;
signal \N__15674\ : std_logic;
signal \N__15671\ : std_logic;
signal \N__15668\ : std_logic;
signal \N__15665\ : std_logic;
signal \N__15662\ : std_logic;
signal \N__15659\ : std_logic;
signal \N__15654\ : std_logic;
signal \N__15649\ : std_logic;
signal \N__15646\ : std_logic;
signal \N__15641\ : std_logic;
signal \N__15638\ : std_logic;
signal \N__15635\ : std_logic;
signal \N__15634\ : std_logic;
signal \N__15631\ : std_logic;
signal \N__15628\ : std_logic;
signal \N__15625\ : std_logic;
signal \N__15622\ : std_logic;
signal \N__15617\ : std_logic;
signal \N__15616\ : std_logic;
signal \N__15613\ : std_logic;
signal \N__15610\ : std_logic;
signal \N__15609\ : std_logic;
signal \N__15606\ : std_logic;
signal \N__15603\ : std_logic;
signal \N__15600\ : std_logic;
signal \N__15599\ : std_logic;
signal \N__15598\ : std_logic;
signal \N__15597\ : std_logic;
signal \N__15596\ : std_logic;
signal \N__15593\ : std_logic;
signal \N__15588\ : std_logic;
signal \N__15585\ : std_logic;
signal \N__15582\ : std_logic;
signal \N__15577\ : std_logic;
signal \N__15566\ : std_logic;
signal \N__15565\ : std_logic;
signal \N__15564\ : std_logic;
signal \N__15561\ : std_logic;
signal \N__15558\ : std_logic;
signal \N__15555\ : std_logic;
signal \N__15552\ : std_logic;
signal \N__15549\ : std_logic;
signal \N__15548\ : std_logic;
signal \N__15547\ : std_logic;
signal \N__15546\ : std_logic;
signal \N__15543\ : std_logic;
signal \N__15538\ : std_logic;
signal \N__15533\ : std_logic;
signal \N__15530\ : std_logic;
signal \N__15529\ : std_logic;
signal \N__15526\ : std_logic;
signal \N__15521\ : std_logic;
signal \N__15518\ : std_logic;
signal \N__15515\ : std_logic;
signal \N__15506\ : std_logic;
signal \N__15503\ : std_logic;
signal \N__15502\ : std_logic;
signal \N__15501\ : std_logic;
signal \N__15500\ : std_logic;
signal \N__15499\ : std_logic;
signal \N__15496\ : std_logic;
signal \N__15495\ : std_logic;
signal \N__15492\ : std_logic;
signal \N__15487\ : std_logic;
signal \N__15484\ : std_logic;
signal \N__15481\ : std_logic;
signal \N__15478\ : std_logic;
signal \N__15477\ : std_logic;
signal \N__15474\ : std_logic;
signal \N__15471\ : std_logic;
signal \N__15468\ : std_logic;
signal \N__15463\ : std_logic;
signal \N__15460\ : std_logic;
signal \N__15455\ : std_logic;
signal \N__15450\ : std_logic;
signal \N__15443\ : std_logic;
signal \N__15440\ : std_logic;
signal \N__15437\ : std_logic;
signal \N__15434\ : std_logic;
signal \N__15431\ : std_logic;
signal \N__15428\ : std_logic;
signal \N__15425\ : std_logic;
signal \N__15422\ : std_logic;
signal \N__15419\ : std_logic;
signal \N__15416\ : std_logic;
signal \N__15413\ : std_logic;
signal \N__15410\ : std_logic;
signal \N__15409\ : std_logic;
signal \N__15406\ : std_logic;
signal \N__15403\ : std_logic;
signal \N__15398\ : std_logic;
signal \N__15397\ : std_logic;
signal \N__15396\ : std_logic;
signal \N__15393\ : std_logic;
signal \N__15392\ : std_logic;
signal \N__15387\ : std_logic;
signal \N__15384\ : std_logic;
signal \N__15381\ : std_logic;
signal \N__15378\ : std_logic;
signal \N__15377\ : std_logic;
signal \N__15376\ : std_logic;
signal \N__15371\ : std_logic;
signal \N__15368\ : std_logic;
signal \N__15363\ : std_logic;
signal \N__15356\ : std_logic;
signal \N__15353\ : std_logic;
signal \N__15352\ : std_logic;
signal \N__15349\ : std_logic;
signal \N__15346\ : std_logic;
signal \N__15345\ : std_logic;
signal \N__15344\ : std_logic;
signal \N__15343\ : std_logic;
signal \N__15342\ : std_logic;
signal \N__15337\ : std_logic;
signal \N__15332\ : std_logic;
signal \N__15327\ : std_logic;
signal \N__15320\ : std_logic;
signal \N__15319\ : std_logic;
signal \N__15316\ : std_logic;
signal \N__15313\ : std_logic;
signal \N__15310\ : std_logic;
signal \N__15307\ : std_logic;
signal \N__15306\ : std_logic;
signal \N__15305\ : std_logic;
signal \N__15302\ : std_logic;
signal \N__15299\ : std_logic;
signal \N__15294\ : std_logic;
signal \N__15287\ : std_logic;
signal \N__15284\ : std_logic;
signal \N__15281\ : std_logic;
signal \N__15280\ : std_logic;
signal \N__15277\ : std_logic;
signal \N__15274\ : std_logic;
signal \N__15273\ : std_logic;
signal \N__15272\ : std_logic;
signal \N__15271\ : std_logic;
signal \N__15266\ : std_logic;
signal \N__15263\ : std_logic;
signal \N__15262\ : std_logic;
signal \N__15257\ : std_logic;
signal \N__15254\ : std_logic;
signal \N__15251\ : std_logic;
signal \N__15248\ : std_logic;
signal \N__15239\ : std_logic;
signal \N__15238\ : std_logic;
signal \N__15237\ : std_logic;
signal \N__15236\ : std_logic;
signal \N__15233\ : std_logic;
signal \N__15230\ : std_logic;
signal \N__15227\ : std_logic;
signal \N__15226\ : std_logic;
signal \N__15225\ : std_logic;
signal \N__15220\ : std_logic;
signal \N__15215\ : std_logic;
signal \N__15212\ : std_logic;
signal \N__15209\ : std_logic;
signal \N__15200\ : std_logic;
signal \N__15199\ : std_logic;
signal \N__15198\ : std_logic;
signal \N__15197\ : std_logic;
signal \N__15194\ : std_logic;
signal \N__15193\ : std_logic;
signal \N__15190\ : std_logic;
signal \N__15187\ : std_logic;
signal \N__15184\ : std_logic;
signal \N__15181\ : std_logic;
signal \N__15178\ : std_logic;
signal \N__15175\ : std_logic;
signal \N__15172\ : std_logic;
signal \N__15171\ : std_logic;
signal \N__15166\ : std_logic;
signal \N__15163\ : std_logic;
signal \N__15158\ : std_logic;
signal \N__15155\ : std_logic;
signal \N__15152\ : std_logic;
signal \N__15147\ : std_logic;
signal \N__15140\ : std_logic;
signal \N__15139\ : std_logic;
signal \N__15136\ : std_logic;
signal \N__15133\ : std_logic;
signal \N__15132\ : std_logic;
signal \N__15127\ : std_logic;
signal \N__15124\ : std_logic;
signal \N__15123\ : std_logic;
signal \N__15122\ : std_logic;
signal \N__15121\ : std_logic;
signal \N__15118\ : std_logic;
signal \N__15115\ : std_logic;
signal \N__15108\ : std_logic;
signal \N__15101\ : std_logic;
signal \N__15098\ : std_logic;
signal \N__15095\ : std_logic;
signal \N__15092\ : std_logic;
signal \N__15089\ : std_logic;
signal \N__15088\ : std_logic;
signal \N__15087\ : std_logic;
signal \N__15084\ : std_logic;
signal \N__15081\ : std_logic;
signal \N__15078\ : std_logic;
signal \N__15073\ : std_logic;
signal \N__15068\ : std_logic;
signal \N__15065\ : std_logic;
signal \N__15062\ : std_logic;
signal \N__15059\ : std_logic;
signal \N__15056\ : std_logic;
signal \N__15053\ : std_logic;
signal \N__15050\ : std_logic;
signal \N__15047\ : std_logic;
signal \N__15044\ : std_logic;
signal \N__15043\ : std_logic;
signal \N__15042\ : std_logic;
signal \N__15041\ : std_logic;
signal \N__15038\ : std_logic;
signal \N__15035\ : std_logic;
signal \N__15030\ : std_logic;
signal \N__15023\ : std_logic;
signal \N__15020\ : std_logic;
signal \N__15019\ : std_logic;
signal \N__15018\ : std_logic;
signal \N__15017\ : std_logic;
signal \N__15014\ : std_logic;
signal \N__15007\ : std_logic;
signal \N__15002\ : std_logic;
signal \N__14999\ : std_logic;
signal \N__14996\ : std_logic;
signal \N__14993\ : std_logic;
signal \N__14990\ : std_logic;
signal \N__14987\ : std_logic;
signal \N__14984\ : std_logic;
signal \N__14981\ : std_logic;
signal \N__14978\ : std_logic;
signal \N__14975\ : std_logic;
signal \N__14972\ : std_logic;
signal \N__14969\ : std_logic;
signal \N__14966\ : std_logic;
signal \N__14963\ : std_logic;
signal \N__14960\ : std_logic;
signal \N__14957\ : std_logic;
signal \N__14954\ : std_logic;
signal \N__14951\ : std_logic;
signal \N__14948\ : std_logic;
signal \N__14945\ : std_logic;
signal \N__14942\ : std_logic;
signal \N__14939\ : std_logic;
signal \N__14936\ : std_logic;
signal \N__14933\ : std_logic;
signal \N__14930\ : std_logic;
signal \N__14927\ : std_logic;
signal \N__14924\ : std_logic;
signal \N__14921\ : std_logic;
signal \N__14918\ : std_logic;
signal \N__14915\ : std_logic;
signal \N__14912\ : std_logic;
signal \N__14909\ : std_logic;
signal \N__14906\ : std_logic;
signal \N__14903\ : std_logic;
signal \N__14900\ : std_logic;
signal \N__14897\ : std_logic;
signal \N__14896\ : std_logic;
signal \N__14895\ : std_logic;
signal \N__14892\ : std_logic;
signal \N__14889\ : std_logic;
signal \N__14886\ : std_logic;
signal \N__14881\ : std_logic;
signal \N__14876\ : std_logic;
signal \N__14875\ : std_logic;
signal \N__14872\ : std_logic;
signal \N__14869\ : std_logic;
signal \N__14866\ : std_logic;
signal \N__14865\ : std_logic;
signal \N__14864\ : std_logic;
signal \N__14861\ : std_logic;
signal \N__14858\ : std_logic;
signal \N__14853\ : std_logic;
signal \N__14846\ : std_logic;
signal \N__14843\ : std_logic;
signal \N__14840\ : std_logic;
signal \N__14837\ : std_logic;
signal \N__14834\ : std_logic;
signal \N__14833\ : std_logic;
signal \N__14832\ : std_logic;
signal \N__14825\ : std_logic;
signal \N__14822\ : std_logic;
signal \N__14819\ : std_logic;
signal \N__14816\ : std_logic;
signal \N__14813\ : std_logic;
signal \N__14812\ : std_logic;
signal \N__14811\ : std_logic;
signal \N__14808\ : std_logic;
signal \N__14803\ : std_logic;
signal \N__14800\ : std_logic;
signal \N__14797\ : std_logic;
signal \N__14792\ : std_logic;
signal \N__14791\ : std_logic;
signal \N__14790\ : std_logic;
signal \N__14789\ : std_logic;
signal \N__14788\ : std_logic;
signal \N__14787\ : std_logic;
signal \N__14786\ : std_logic;
signal \N__14785\ : std_logic;
signal \N__14784\ : std_logic;
signal \N__14783\ : std_logic;
signal \N__14780\ : std_logic;
signal \N__14779\ : std_logic;
signal \N__14778\ : std_logic;
signal \N__14777\ : std_logic;
signal \N__14774\ : std_logic;
signal \N__14771\ : std_logic;
signal \N__14768\ : std_logic;
signal \N__14765\ : std_logic;
signal \N__14762\ : std_logic;
signal \N__14755\ : std_logic;
signal \N__14754\ : std_logic;
signal \N__14753\ : std_logic;
signal \N__14752\ : std_logic;
signal \N__14751\ : std_logic;
signal \N__14740\ : std_logic;
signal \N__14737\ : std_logic;
signal \N__14734\ : std_logic;
signal \N__14731\ : std_logic;
signal \N__14726\ : std_logic;
signal \N__14723\ : std_logic;
signal \N__14714\ : std_logic;
signal \N__14711\ : std_logic;
signal \N__14708\ : std_logic;
signal \N__14705\ : std_logic;
signal \N__14698\ : std_logic;
signal \N__14687\ : std_logic;
signal \N__14684\ : std_logic;
signal \N__14683\ : std_logic;
signal \N__14680\ : std_logic;
signal \N__14677\ : std_logic;
signal \N__14674\ : std_logic;
signal \N__14671\ : std_logic;
signal \N__14666\ : std_logic;
signal \N__14663\ : std_logic;
signal \N__14660\ : std_logic;
signal \N__14657\ : std_logic;
signal \N__14654\ : std_logic;
signal \N__14651\ : std_logic;
signal \N__14648\ : std_logic;
signal \N__14645\ : std_logic;
signal \N__14642\ : std_logic;
signal \N__14641\ : std_logic;
signal \N__14640\ : std_logic;
signal \N__14637\ : std_logic;
signal \N__14632\ : std_logic;
signal \N__14629\ : std_logic;
signal \N__14626\ : std_logic;
signal \N__14621\ : std_logic;
signal \N__14618\ : std_logic;
signal \N__14617\ : std_logic;
signal \N__14616\ : std_logic;
signal \N__14613\ : std_logic;
signal \N__14610\ : std_logic;
signal \N__14607\ : std_logic;
signal \N__14604\ : std_logic;
signal \N__14601\ : std_logic;
signal \N__14594\ : std_logic;
signal \N__14591\ : std_logic;
signal \N__14590\ : std_logic;
signal \N__14587\ : std_logic;
signal \N__14584\ : std_logic;
signal \N__14583\ : std_logic;
signal \N__14580\ : std_logic;
signal \N__14577\ : std_logic;
signal \N__14574\ : std_logic;
signal \N__14571\ : std_logic;
signal \N__14568\ : std_logic;
signal \N__14561\ : std_logic;
signal \N__14558\ : std_logic;
signal \N__14557\ : std_logic;
signal \N__14554\ : std_logic;
signal \N__14551\ : std_logic;
signal \N__14548\ : std_logic;
signal \N__14543\ : std_logic;
signal \N__14540\ : std_logic;
signal \N__14539\ : std_logic;
signal \N__14536\ : std_logic;
signal \N__14533\ : std_logic;
signal \N__14528\ : std_logic;
signal \N__14525\ : std_logic;
signal \N__14522\ : std_logic;
signal \N__14519\ : std_logic;
signal \N__14516\ : std_logic;
signal \N__14513\ : std_logic;
signal \N__14510\ : std_logic;
signal \N__14507\ : std_logic;
signal \N__14504\ : std_logic;
signal \N__14501\ : std_logic;
signal \N__14498\ : std_logic;
signal \N__14495\ : std_logic;
signal \N__14492\ : std_logic;
signal \N__14489\ : std_logic;
signal \N__14486\ : std_logic;
signal \N__14483\ : std_logic;
signal \N__14480\ : std_logic;
signal \N__14477\ : std_logic;
signal \N__14474\ : std_logic;
signal \N__14471\ : std_logic;
signal \N__14468\ : std_logic;
signal \N__14465\ : std_logic;
signal \N__14462\ : std_logic;
signal \N__14459\ : std_logic;
signal \N__14456\ : std_logic;
signal \N__14453\ : std_logic;
signal \N__14452\ : std_logic;
signal \N__14449\ : std_logic;
signal \N__14446\ : std_logic;
signal \N__14443\ : std_logic;
signal \N__14440\ : std_logic;
signal \N__14437\ : std_logic;
signal \N__14434\ : std_logic;
signal \N__14431\ : std_logic;
signal \N__14428\ : std_logic;
signal \N__14425\ : std_logic;
signal \N__14422\ : std_logic;
signal \N__14419\ : std_logic;
signal \N__14416\ : std_logic;
signal \N__14413\ : std_logic;
signal \N__14410\ : std_logic;
signal \N__14407\ : std_logic;
signal \N__14404\ : std_logic;
signal \N__14401\ : std_logic;
signal \N__14398\ : std_logic;
signal \N__14395\ : std_logic;
signal \N__14392\ : std_logic;
signal \N__14389\ : std_logic;
signal \N__14386\ : std_logic;
signal \N__14383\ : std_logic;
signal \N__14380\ : std_logic;
signal \N__14377\ : std_logic;
signal \N__14374\ : std_logic;
signal \N__14371\ : std_logic;
signal \N__14368\ : std_logic;
signal \N__14365\ : std_logic;
signal \N__14360\ : std_logic;
signal \N__14357\ : std_logic;
signal \N__14356\ : std_logic;
signal \N__14353\ : std_logic;
signal \N__14350\ : std_logic;
signal \N__14347\ : std_logic;
signal \N__14344\ : std_logic;
signal \N__14341\ : std_logic;
signal \N__14338\ : std_logic;
signal \N__14335\ : std_logic;
signal \N__14332\ : std_logic;
signal \N__14329\ : std_logic;
signal \N__14326\ : std_logic;
signal \N__14323\ : std_logic;
signal \N__14320\ : std_logic;
signal \N__14317\ : std_logic;
signal \N__14314\ : std_logic;
signal \N__14311\ : std_logic;
signal \N__14308\ : std_logic;
signal \N__14305\ : std_logic;
signal \N__14302\ : std_logic;
signal \N__14299\ : std_logic;
signal \N__14296\ : std_logic;
signal \N__14293\ : std_logic;
signal \N__14290\ : std_logic;
signal \N__14287\ : std_logic;
signal \N__14284\ : std_logic;
signal \N__14281\ : std_logic;
signal \N__14278\ : std_logic;
signal \N__14275\ : std_logic;
signal \N__14272\ : std_logic;
signal \N__14269\ : std_logic;
signal \N__14264\ : std_logic;
signal \N__14263\ : std_logic;
signal \N__14260\ : std_logic;
signal \N__14257\ : std_logic;
signal \N__14254\ : std_logic;
signal \N__14251\ : std_logic;
signal \N__14248\ : std_logic;
signal \N__14245\ : std_logic;
signal \N__14242\ : std_logic;
signal \N__14239\ : std_logic;
signal \N__14236\ : std_logic;
signal \N__14233\ : std_logic;
signal \N__14230\ : std_logic;
signal \N__14227\ : std_logic;
signal \N__14224\ : std_logic;
signal \N__14221\ : std_logic;
signal \N__14218\ : std_logic;
signal \N__14215\ : std_logic;
signal \N__14212\ : std_logic;
signal \N__14209\ : std_logic;
signal \N__14206\ : std_logic;
signal \N__14203\ : std_logic;
signal \N__14200\ : std_logic;
signal \N__14197\ : std_logic;
signal \N__14194\ : std_logic;
signal \N__14191\ : std_logic;
signal \N__14188\ : std_logic;
signal \N__14185\ : std_logic;
signal \N__14182\ : std_logic;
signal \N__14179\ : std_logic;
signal \N__14176\ : std_logic;
signal \N__14171\ : std_logic;
signal \N__14170\ : std_logic;
signal \N__14167\ : std_logic;
signal \N__14164\ : std_logic;
signal \N__14161\ : std_logic;
signal \N__14158\ : std_logic;
signal \N__14155\ : std_logic;
signal \N__14152\ : std_logic;
signal \N__14149\ : std_logic;
signal \N__14146\ : std_logic;
signal \N__14143\ : std_logic;
signal \N__14140\ : std_logic;
signal \N__14137\ : std_logic;
signal \N__14134\ : std_logic;
signal \N__14131\ : std_logic;
signal \N__14128\ : std_logic;
signal \N__14125\ : std_logic;
signal \N__14122\ : std_logic;
signal \N__14119\ : std_logic;
signal \N__14116\ : std_logic;
signal \N__14113\ : std_logic;
signal \N__14110\ : std_logic;
signal \N__14107\ : std_logic;
signal \N__14104\ : std_logic;
signal \N__14101\ : std_logic;
signal \N__14098\ : std_logic;
signal \N__14095\ : std_logic;
signal \N__14092\ : std_logic;
signal \N__14089\ : std_logic;
signal \N__14086\ : std_logic;
signal \N__14081\ : std_logic;
signal \N__14078\ : std_logic;
signal \N__14075\ : std_logic;
signal \N__14072\ : std_logic;
signal \N__14069\ : std_logic;
signal \N__14068\ : std_logic;
signal \N__14063\ : std_logic;
signal \N__14060\ : std_logic;
signal \N__14057\ : std_logic;
signal \N__14054\ : std_logic;
signal \N__14051\ : std_logic;
signal \N__14048\ : std_logic;
signal \N__14045\ : std_logic;
signal \N__14042\ : std_logic;
signal \N__14039\ : std_logic;
signal \N__14036\ : std_logic;
signal \N__14033\ : std_logic;
signal \N__14032\ : std_logic;
signal \N__14029\ : std_logic;
signal \N__14026\ : std_logic;
signal \N__14021\ : std_logic;
signal \N__14018\ : std_logic;
signal \N__14015\ : std_logic;
signal \N__14012\ : std_logic;
signal \N__14009\ : std_logic;
signal \N__14008\ : std_logic;
signal \N__14005\ : std_logic;
signal \N__14002\ : std_logic;
signal \N__13997\ : std_logic;
signal \N__13994\ : std_logic;
signal \N__13991\ : std_logic;
signal \N__13988\ : std_logic;
signal \N__13987\ : std_logic;
signal \N__13982\ : std_logic;
signal \N__13979\ : std_logic;
signal \N__13976\ : std_logic;
signal \N__13973\ : std_logic;
signal \N__13970\ : std_logic;
signal \N__13969\ : std_logic;
signal \N__13964\ : std_logic;
signal \N__13961\ : std_logic;
signal \N__13958\ : std_logic;
signal \N__13955\ : std_logic;
signal \N__13952\ : std_logic;
signal \N__13949\ : std_logic;
signal \N__13948\ : std_logic;
signal \N__13945\ : std_logic;
signal \N__13942\ : std_logic;
signal \N__13937\ : std_logic;
signal \N__13934\ : std_logic;
signal \N__13931\ : std_logic;
signal \N__13928\ : std_logic;
signal \N__13925\ : std_logic;
signal \N__13922\ : std_logic;
signal \N__13919\ : std_logic;
signal \N__13918\ : std_logic;
signal \N__13915\ : std_logic;
signal \N__13914\ : std_logic;
signal \N__13907\ : std_logic;
signal \N__13904\ : std_logic;
signal \N__13901\ : std_logic;
signal \N__13898\ : std_logic;
signal \N__13895\ : std_logic;
signal \N__13892\ : std_logic;
signal \N__13889\ : std_logic;
signal \N__13886\ : std_logic;
signal \N__13883\ : std_logic;
signal \N__13880\ : std_logic;
signal \N__13877\ : std_logic;
signal \N__13874\ : std_logic;
signal \N__13871\ : std_logic;
signal \N__13868\ : std_logic;
signal \N__13865\ : std_logic;
signal \N__13862\ : std_logic;
signal \N__13859\ : std_logic;
signal \N__13856\ : std_logic;
signal \N__13853\ : std_logic;
signal \N__13852\ : std_logic;
signal \N__13851\ : std_logic;
signal \N__13850\ : std_logic;
signal \N__13849\ : std_logic;
signal \N__13848\ : std_logic;
signal \N__13847\ : std_logic;
signal \N__13846\ : std_logic;
signal \N__13845\ : std_logic;
signal \N__13844\ : std_logic;
signal \N__13823\ : std_logic;
signal \N__13820\ : std_logic;
signal \N__13817\ : std_logic;
signal \N__13814\ : std_logic;
signal \N__13811\ : std_logic;
signal \N__13808\ : std_logic;
signal \N__13805\ : std_logic;
signal \N__13802\ : std_logic;
signal \N__13801\ : std_logic;
signal \N__13798\ : std_logic;
signal \N__13795\ : std_logic;
signal \N__13790\ : std_logic;
signal \N__13787\ : std_logic;
signal \N__13784\ : std_logic;
signal \N__13781\ : std_logic;
signal \N__13778\ : std_logic;
signal \N__13775\ : std_logic;
signal \N__13774\ : std_logic;
signal \N__13771\ : std_logic;
signal \N__13768\ : std_logic;
signal \N__13763\ : std_logic;
signal \N__13760\ : std_logic;
signal \N__13759\ : std_logic;
signal \N__13758\ : std_logic;
signal \N__13755\ : std_logic;
signal \N__13752\ : std_logic;
signal \N__13749\ : std_logic;
signal \N__13748\ : std_logic;
signal \N__13747\ : std_logic;
signal \N__13744\ : std_logic;
signal \N__13743\ : std_logic;
signal \N__13740\ : std_logic;
signal \N__13737\ : std_logic;
signal \N__13732\ : std_logic;
signal \N__13729\ : std_logic;
signal \N__13726\ : std_logic;
signal \N__13721\ : std_logic;
signal \N__13712\ : std_logic;
signal \N__13709\ : std_logic;
signal \N__13706\ : std_logic;
signal \N__13703\ : std_logic;
signal \N__13700\ : std_logic;
signal \N__13697\ : std_logic;
signal \N__13694\ : std_logic;
signal \N__13691\ : std_logic;
signal \N__13690\ : std_logic;
signal \N__13689\ : std_logic;
signal \N__13682\ : std_logic;
signal \N__13679\ : std_logic;
signal \N__13676\ : std_logic;
signal \N__13675\ : std_logic;
signal \N__13672\ : std_logic;
signal \N__13671\ : std_logic;
signal \N__13664\ : std_logic;
signal \N__13661\ : std_logic;
signal \N__13658\ : std_logic;
signal \N__13657\ : std_logic;
signal \N__13656\ : std_logic;
signal \N__13655\ : std_logic;
signal \N__13652\ : std_logic;
signal \N__13645\ : std_logic;
signal \N__13642\ : std_logic;
signal \N__13639\ : std_logic;
signal \N__13634\ : std_logic;
signal \N__13631\ : std_logic;
signal \N__13630\ : std_logic;
signal \N__13627\ : std_logic;
signal \N__13624\ : std_logic;
signal \N__13621\ : std_logic;
signal \N__13616\ : std_logic;
signal \N__13613\ : std_logic;
signal \N__13612\ : std_logic;
signal \N__13609\ : std_logic;
signal \N__13606\ : std_logic;
signal \N__13605\ : std_logic;
signal \N__13602\ : std_logic;
signal \N__13597\ : std_logic;
signal \N__13592\ : std_logic;
signal \N__13589\ : std_logic;
signal \N__13586\ : std_logic;
signal \N__13583\ : std_logic;
signal \N__13580\ : std_logic;
signal \N__13577\ : std_logic;
signal \N__13574\ : std_logic;
signal \N__13571\ : std_logic;
signal \N__13568\ : std_logic;
signal \N__13565\ : std_logic;
signal \N__13562\ : std_logic;
signal \N__13559\ : std_logic;
signal \N__13556\ : std_logic;
signal \N__13553\ : std_logic;
signal \N__13550\ : std_logic;
signal \N__13547\ : std_logic;
signal \N__13544\ : std_logic;
signal \N__13541\ : std_logic;
signal \N__13538\ : std_logic;
signal \N__13535\ : std_logic;
signal \N__13532\ : std_logic;
signal \N__13529\ : std_logic;
signal \N__13526\ : std_logic;
signal \N__13523\ : std_logic;
signal \N__13520\ : std_logic;
signal \N__13517\ : std_logic;
signal \N__13514\ : std_logic;
signal \N__13511\ : std_logic;
signal \N__13508\ : std_logic;
signal \N__13505\ : std_logic;
signal \N__13502\ : std_logic;
signal \N__13499\ : std_logic;
signal \N__13496\ : std_logic;
signal \N__13493\ : std_logic;
signal \N__13490\ : std_logic;
signal \N__13487\ : std_logic;
signal \N__13484\ : std_logic;
signal \N__13481\ : std_logic;
signal \N__13478\ : std_logic;
signal \N__13475\ : std_logic;
signal \N__13472\ : std_logic;
signal \N__13469\ : std_logic;
signal \N__13466\ : std_logic;
signal \N__13465\ : std_logic;
signal \N__13462\ : std_logic;
signal \N__13459\ : std_logic;
signal \N__13454\ : std_logic;
signal \N__13451\ : std_logic;
signal \N__13448\ : std_logic;
signal \N__13445\ : std_logic;
signal \N__13444\ : std_logic;
signal \N__13441\ : std_logic;
signal \N__13438\ : std_logic;
signal \N__13433\ : std_logic;
signal \N__13430\ : std_logic;
signal \N__13427\ : std_logic;
signal \N__13424\ : std_logic;
signal \N__13421\ : std_logic;
signal \N__13418\ : std_logic;
signal \N__13415\ : std_logic;
signal \N__13412\ : std_logic;
signal \N__13409\ : std_logic;
signal \N__13406\ : std_logic;
signal \N__13403\ : std_logic;
signal \N__13400\ : std_logic;
signal \N__13397\ : std_logic;
signal \N__13394\ : std_logic;
signal \N__13393\ : std_logic;
signal \N__13392\ : std_logic;
signal \N__13389\ : std_logic;
signal \N__13384\ : std_logic;
signal \N__13379\ : std_logic;
signal \N__13376\ : std_logic;
signal \N__13375\ : std_logic;
signal \N__13374\ : std_logic;
signal \N__13371\ : std_logic;
signal \N__13368\ : std_logic;
signal \N__13365\ : std_logic;
signal \N__13362\ : std_logic;
signal \N__13355\ : std_logic;
signal \N__13352\ : std_logic;
signal \N__13349\ : std_logic;
signal \N__13346\ : std_logic;
signal \N__13343\ : std_logic;
signal \N__13340\ : std_logic;
signal \N__13337\ : std_logic;
signal \N__13334\ : std_logic;
signal \N__13331\ : std_logic;
signal \N__13328\ : std_logic;
signal \N__13325\ : std_logic;
signal \N__13322\ : std_logic;
signal \N__13319\ : std_logic;
signal \N__13316\ : std_logic;
signal \N__13313\ : std_logic;
signal \N__13310\ : std_logic;
signal \N__13307\ : std_logic;
signal \N__13304\ : std_logic;
signal \N__13301\ : std_logic;
signal \N__13298\ : std_logic;
signal \N__13295\ : std_logic;
signal \N__13292\ : std_logic;
signal \N__13289\ : std_logic;
signal \N__13286\ : std_logic;
signal \N__13283\ : std_logic;
signal \N__13280\ : std_logic;
signal \N__13277\ : std_logic;
signal \N__13274\ : std_logic;
signal \N__13271\ : std_logic;
signal \N__13268\ : std_logic;
signal \N__13265\ : std_logic;
signal \N__13262\ : std_logic;
signal \N__13259\ : std_logic;
signal \N__13256\ : std_logic;
signal \N__13253\ : std_logic;
signal \N__13250\ : std_logic;
signal \N__13247\ : std_logic;
signal \N__13244\ : std_logic;
signal \N__13241\ : std_logic;
signal \N__13238\ : std_logic;
signal \N__13235\ : std_logic;
signal \N__13232\ : std_logic;
signal \N__13229\ : std_logic;
signal \N__13226\ : std_logic;
signal \N__13223\ : std_logic;
signal \N__13220\ : std_logic;
signal \N__13217\ : std_logic;
signal \N__13214\ : std_logic;
signal \N__13211\ : std_logic;
signal \N__13208\ : std_logic;
signal \N__13205\ : std_logic;
signal \N__13202\ : std_logic;
signal \N__13199\ : std_logic;
signal \N__13196\ : std_logic;
signal \N__13193\ : std_logic;
signal \N__13190\ : std_logic;
signal \N__13187\ : std_logic;
signal \N__13184\ : std_logic;
signal \N__13181\ : std_logic;
signal \N__13178\ : std_logic;
signal \N__13175\ : std_logic;
signal \N__13172\ : std_logic;
signal \N__13169\ : std_logic;
signal \N__13166\ : std_logic;
signal \N__13163\ : std_logic;
signal \N__13162\ : std_logic;
signal \N__13161\ : std_logic;
signal \N__13156\ : std_logic;
signal \N__13153\ : std_logic;
signal \N__13148\ : std_logic;
signal \N__13145\ : std_logic;
signal \N__13142\ : std_logic;
signal \N__13141\ : std_logic;
signal \N__13140\ : std_logic;
signal \N__13133\ : std_logic;
signal \N__13130\ : std_logic;
signal \N__13129\ : std_logic;
signal \N__13126\ : std_logic;
signal \N__13125\ : std_logic;
signal \N__13122\ : std_logic;
signal \N__13115\ : std_logic;
signal \N__13112\ : std_logic;
signal \N__13109\ : std_logic;
signal \N__13106\ : std_logic;
signal \N__13103\ : std_logic;
signal \N__13100\ : std_logic;
signal \N__13097\ : std_logic;
signal \N__13096\ : std_logic;
signal \N__13095\ : std_logic;
signal \N__13088\ : std_logic;
signal \N__13085\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \b2v_inst.N_4_i_i_a3_0_0_cascade_\ : std_logic;
signal \b2v_inst.un4_pix_count_intlto6_d_1_1_cascade_\ : std_logic;
signal b2v_inst4_pix_count_int_fast_1 : std_logic;
signal b2v_inst4_pix_count_int_fast_0 : std_logic;
signal \b2v_inst.N_13\ : std_logic;
signal b2v_inst4_pix_count_int_fast_2 : std_logic;
signal b2v_inst4_pix_count_int_fast_3 : std_logic;
signal \b2v_inst.pix_count_anteriorZ0Z_1\ : std_logic;
signal \b2v_inst.pix_count_anteriorZ0Z_4\ : std_logic;
signal \b2v_inst.un7_pix_count_int_0_I_1_c_RNOZ0\ : std_logic;
signal \bfn_2_11_0_\ : std_logic;
signal \b2v_inst.un7_pix_count_int_0_data_tmp_0\ : std_logic;
signal \b2v_inst.un7_pix_count_int_0_I_15_c_RNOZ0\ : std_logic;
signal \b2v_inst.un7_pix_count_int_0_data_tmp_1\ : std_logic;
signal \b2v_inst.un7_pix_count_int_0_data_tmp_2\ : std_logic;
signal \b2v_inst.un7_pix_count_int_0_data_tmp_3\ : std_logic;
signal \b2v_inst.un7_pix_count_int_0_data_tmp_4\ : std_logic;
signal \b2v_inst.un7_pix_count_int_0_data_tmp_5\ : std_logic;
signal \b2v_inst.un7_pix_count_int_0_data_tmp_6\ : std_logic;
signal \b2v_inst.un7_pix_count_int_0_data_tmp_7\ : std_logic;
signal \bfn_2_12_0_\ : std_logic;
signal \b2v_inst.un7_pix_count_int_0_data_tmp_8\ : std_logic;
signal \b2v_inst.un7_pix_count_int_0_N_2\ : std_logic;
signal \b2v_inst.un7_pix_count_int_0_I_57_c_RNOZ0\ : std_logic;
signal \b2v_inst4.un1_pix_count_int_0_sqmuxa_6\ : std_logic;
signal \b2v_inst.un7_pix_count_int_0_I_27_c_RNOZ0\ : std_logic;
signal \b2v_inst.pix_count_anteriorZ0Z_2\ : std_logic;
signal \b2v_inst.pix_count_anteriorZ0Z_3\ : std_logic;
signal \b2v_inst.pix_count_anteriorZ0Z_0\ : std_logic;
signal \b2v_inst.pix_count_anteriorZ0Z_5\ : std_logic;
signal \b2v_inst.un7_pix_count_int_0_I_33_c_RNOZ0\ : std_logic;
signal \b2v_inst.pix_count_anteriorZ0Z_18\ : std_logic;
signal \b2v_inst.un7_pix_count_int_0_I_39_c_RNOZ0\ : std_logic;
signal \b2v_inst.pix_count_anteriorZ0Z_12\ : std_logic;
signal \b2v_inst.pix_count_anteriorZ0Z_13\ : std_logic;
signal \b2v_inst.un7_pix_count_int_0_I_45_c_RNOZ0\ : std_logic;
signal \b2v_inst.pix_count_anteriorZ0Z_14\ : std_logic;
signal \b2v_inst4.un1_pix_count_int_0_sqmuxa_5_cascade_\ : std_logic;
signal \b2v_inst.pix_count_anteriorZ0Z_15\ : std_logic;
signal \b2v_inst.pix_count_anteriorZ0Z_19\ : std_logic;
signal \b2v_inst.pix_count_anteriorZ0Z_16\ : std_logic;
signal \b2v_inst.un1_state_36_0_a2_0_2_1_cascade_\ : std_logic;
signal \b2v_inst.N_305_2\ : std_logic;
signal \b2v_inst.N_305_2_cascade_\ : std_logic;
signal \b2v_inst.cuenta_pixelZ0Z_1\ : std_logic;
signal \bfn_3_10_0_\ : std_logic;
signal \b2v_inst.un1_cuenta_pixel_cry_1\ : std_logic;
signal \b2v_inst.un1_cuenta_pixel_cry_2\ : std_logic;
signal \b2v_inst.un1_cuenta_pixel_cry_3\ : std_logic;
signal \b2v_inst.un1_cuenta_pixel_cry_4\ : std_logic;
signal \b2v_inst.cuenta_pixelZ0Z_6\ : std_logic;
signal \b2v_inst.un1_cuenta_pixel_cry_5_c_RNIGL1IZ0\ : std_logic;
signal \b2v_inst.un1_cuenta_pixel_cry_5\ : std_logic;
signal \b2v_inst.cuenta_pixelZ0Z_7\ : std_logic;
signal \b2v_inst.un1_cuenta_pixel_cry_6_c_RNIIO2IZ0\ : std_logic;
signal \b2v_inst.un1_cuenta_pixel_cry_6\ : std_logic;
signal \b2v_inst.cuenta_pixelZ0Z_8\ : std_logic;
signal \b2v_inst.un1_cuenta_pixel_cry_7\ : std_logic;
signal \b2v_inst.un1_cuenta_pixel_cry_8\ : std_logic;
signal \b2v_inst.cuenta_pixelZ0Z_9\ : std_logic;
signal \bfn_3_11_0_\ : std_logic;
signal \b2v_inst.un1_cuenta_pixel_cry_9\ : std_logic;
signal \b2v_inst.cuenta_pixelZ0Z_10\ : std_logic;
signal \b2v_inst.pix_count_anteriorZ0Z_9\ : std_logic;
signal \b2v_inst.un7_pix_count_int_0_I_51_c_RNOZ0\ : std_logic;
signal \b2v_inst.N_1_0_0_cascade_\ : std_logic;
signal \b2v_inst.N_4_i_i_o6_2_cascade_\ : std_logic;
signal \b2v_inst.N_7\ : std_logic;
signal \b2v_inst.un7_pix_count_int_0_I_21_c_RNOZ0\ : std_logic;
signal \b2v_inst.pix_count_anteriorZ0Z_6\ : std_logic;
signal \b2v_inst.pix_count_anteriorZ0Z_7\ : std_logic;
signal \b2v_inst.pix_count_anteriorZ0Z_8\ : std_logic;
signal \b2v_inst4.un1_pix_count_int_0_sqmuxa_7\ : std_logic;
signal \b2v_inst4.un1_pix_count_int_0_sqmuxa_13\ : std_logic;
signal \b2v_inst4.un1_pix_count_int_0_sqmuxa_8_cascade_\ : std_logic;
signal \b2v_inst4.un1_pix_count_int_0_sqmuxa_14\ : std_logic;
signal \b2v_inst4.un1_pix_count_int_0_sqmuxa_10\ : std_logic;
signal \b2v_inst.cuenta_pixel_RNIT0FMZ0Z_1\ : std_logic;
signal \b2v_inst.cuenta_pixelZ0Z_0\ : std_logic;
signal \b2v_inst.cuenta_pixel_5_i_a2_0_2_5_cascade_\ : std_logic;
signal \b2v_inst.cuenta_pixelZ0Z_2\ : std_logic;
signal \b2v_inst.cuenta_pixelZ0Z_3\ : std_logic;
signal \b2v_inst.un1_cuenta_pixel_cry_1_c_RNI89THZ0\ : std_logic;
signal \b2v_inst.un1_cuenta_pixel_cry_2_c_RNIACUHZ0\ : std_logic;
signal \b2v_inst.un1_cuenta_pixel_cry_4_c_RNIEI0IZ0\ : std_logic;
signal \b2v_inst.cuenta_pixel_5_i_a2_0_2_5\ : std_logic;
signal \b2v_inst.cuenta_pixel_5_i_a2_0_1_5\ : std_logic;
signal \b2v_inst.cuenta_pixelZ0Z_5\ : std_logic;
signal \b2v_inst.un1_cuenta_pixel_cry_3_c_RNICFVHZ0\ : std_logic;
signal \b2v_inst.cuenta_pixelZ0Z_4\ : std_logic;
signal \b2v_inst.un7_pix_count_int_0_I_9_c_RNOZ0\ : std_logic;
signal \b2v_inst.pix_count_anteriorZ0Z_10\ : std_logic;
signal \b2v_inst.pix_count_anteriorZ0Z_11\ : std_logic;
signal \b2v_inst.pix_count_anteriorZ0Z_17\ : std_logic;
signal \b2v_inst.N_305_1_g\ : std_logic;
signal \b2v_inst.N_4_i_i_a6_1\ : std_logic;
signal \b2v_inst4.pix_count_int_RNI0EPTZ0Z_0\ : std_logic;
signal \bfn_5_13_0_\ : std_logic;
signal \b2v_inst4.un1_pix_count_int_cry_0_c_RNIIC2IZ0\ : std_logic;
signal \b2v_inst4.un1_pix_count_int_cry_0\ : std_logic;
signal \b2v_inst4.un1_pix_count_int_cry_1_c_RNIKF3IZ0\ : std_logic;
signal \b2v_inst4.un1_pix_count_int_cry_1\ : std_logic;
signal \b2v_inst4.un1_pix_count_int_cry_2_c_RNIMI4IZ0\ : std_logic;
signal \b2v_inst4.un1_pix_count_int_cry_2\ : std_logic;
signal \b2v_inst4.un1_pix_count_int_cry_3\ : std_logic;
signal \b2v_inst4.un1_pix_count_int_cry_4_c_RNIQO6IZ0\ : std_logic;
signal \b2v_inst4.un1_pix_count_int_cry_4\ : std_logic;
signal \b2v_inst4.un1_pix_count_int_cry_5_c_RNISR7IZ0\ : std_logic;
signal \b2v_inst4.un1_pix_count_int_cry_5\ : std_logic;
signal \b2v_inst4.un1_pix_count_int_cry_6\ : std_logic;
signal \b2v_inst4.un1_pix_count_int_cry_7\ : std_logic;
signal \bfn_5_14_0_\ : std_logic;
signal \b2v_inst4.un1_pix_count_int_cry_8\ : std_logic;
signal \b2v_inst4.un1_pix_count_int_cry_9\ : std_logic;
signal \b2v_inst4.un1_pix_count_int_cry_10\ : std_logic;
signal \b2v_inst4.un1_pix_count_int_cry_11_c_RNIMPVJZ0\ : std_logic;
signal \b2v_inst4.un1_pix_count_int_cry_11\ : std_logic;
signal \b2v_inst4.un1_pix_count_int_cry_12\ : std_logic;
signal \b2v_inst4.un1_pix_count_int_cry_13\ : std_logic;
signal \b2v_inst4.un1_pix_count_int_cry_14\ : std_logic;
signal \b2v_inst4.un1_pix_count_int_cry_15\ : std_logic;
signal \bfn_5_15_0_\ : std_logic;
signal \b2v_inst4.un1_pix_count_int_cry_16\ : std_logic;
signal \b2v_inst4.un1_pix_count_int_cry_17\ : std_logic;
signal \b2v_inst4.un1_pix_count_int_cry_18\ : std_logic;
signal \SYNTHESIZED_WIRE_12_1\ : std_logic;
signal \SYNTHESIZED_WIRE_12_7\ : std_logic;
signal \SYNTHESIZED_WIRE_12_0\ : std_logic;
signal \SYNTHESIZED_WIRE_12_8\ : std_logic;
signal \bfn_6_5_0_\ : std_logic;
signal \b2v_inst.un2_dir_mem_3_cry_0\ : std_logic;
signal \b2v_inst.un2_dir_mem_3_cry_1\ : std_logic;
signal \b2v_inst.un2_dir_mem_3_cry_2\ : std_logic;
signal \b2v_inst.un2_dir_mem_3_cry_3\ : std_logic;
signal \b2v_inst.un2_dir_mem_3_cry_4\ : std_logic;
signal \bfn_6_6_0_\ : std_logic;
signal \b2v_inst.un1_indice_cry_1\ : std_logic;
signal \b2v_inst.un1_indice_cry_2\ : std_logic;
signal \b2v_inst.un1_indice_cry_3\ : std_logic;
signal \b2v_inst.un1_indice_cry_4\ : std_logic;
signal \b2v_inst.un1_indice_cry_5\ : std_logic;
signal \b2v_inst.un1_indice_cry_6\ : std_logic;
signal \b2v_inst.un1_indice_cry_7\ : std_logic;
signal \b2v_inst.un1_indice_cry_8\ : std_logic;
signal \bfn_6_7_0_\ : std_logic;
signal \b2v_inst.un1_indice_cry_9\ : std_logic;
signal \b2v_inst.un1_indice_cry_10\ : std_logic;
signal \b2v_inst.ignorar_ancho_1_RNOZ0Z_1\ : std_logic;
signal \b2v_inst.ignorar_ancho_1_RNOZ0Z_2\ : std_logic;
signal \b2v_inst4.un1_pix_count_int_cry_9_c_RNIB86JZ0\ : std_logic;
signal \b2v_inst4.un1_pix_count_int_cry_8_c_RNI25BIZ0\ : std_logic;
signal \b2v_inst4.un1_pix_count_int_0_sqmuxa_0\ : std_logic;
signal \b2v_inst4.un1_pix_count_int_cry_10_c_RNIKMUJZ0\ : std_logic;
signal \b2v_inst.ignorar_ancho_1_RNOZ0Z_0\ : std_logic;
signal \b2v_inst.N_482_cascade_\ : std_logic;
signal \b2v_inst.un1_state_34_0\ : std_logic;
signal \b2v_inst.un1_cuenta_pixel_cry_8_c_RNIMU4IZ0\ : std_logic;
signal \b2v_inst.cuenta_pixel_RNIVBL9Z0Z_10\ : std_logic;
signal \b2v_inst.un1_cuenta_pixel_cry_7_c_RNIKR3IZ0\ : std_logic;
signal \b2v_inst.cuenta_pixel_5_i_a2_1_1_0_5\ : std_logic;
signal \b2v_inst.N_325\ : std_logic;
signal \b2v_inst.un1_state_36_0_rn_1\ : std_logic;
signal \b2v_inst.un1_state_36_0_sn\ : std_logic;
signal \b2v_inst.N_325_cascade_\ : std_logic;
signal \b2v_inst.N_305_1\ : std_logic;
signal \b2v_inst.un1_state_36_0\ : std_logic;
signal \b2v_inst4.stateZ0Z_0\ : std_logic;
signal \SYNTHESIZED_WIRE_9\ : std_logic;
signal \b2v_inst.un1_state_36_0_a2_0_1_mbZ0Z_1\ : std_logic;
signal \b2v_inst1.N_40\ : std_logic;
signal \bfn_7_6_0_\ : std_logic;
signal \b2v_inst.un8_dir_mem_1_cry_0\ : std_logic;
signal \b2v_inst.un8_dir_mem_1_cry_1\ : std_logic;
signal \b2v_inst.un8_dir_mem_1_cry_2\ : std_logic;
signal \b2v_inst.un8_dir_mem_1_cry_3\ : std_logic;
signal \b2v_inst.un8_dir_mem_1_cry_4\ : std_logic;
signal \b2v_inst.un8_dir_mem_1_cry_5\ : std_logic;
signal \b2v_inst.un8_dir_mem_1_cry_6\ : std_logic;
signal \b2v_inst.un8_dir_mem_1_cry_7\ : std_logic;
signal \bfn_7_7_0_\ : std_logic;
signal \b2v_inst.un8_dir_mem_1_cry_8\ : std_logic;
signal \b2v_inst.un8_dir_mem_1_cry_9\ : std_logic;
signal \b2v_inst.un8_dir_mem_1_cry_10\ : std_logic;
signal \b2v_inst.dir_mem_316lt6_0_cascade_\ : std_logic;
signal \b2v_inst.dir_mem_316lt7\ : std_logic;
signal \b2v_inst.un1_indice_cry_1_c_RNIUSJGZ0\ : std_logic;
signal \SYNTHESIZED_WIRE_4_fast_10\ : std_logic;
signal \SYNTHESIZED_WIRE_4_fast_9\ : std_logic;
signal \b2v_inst.N_9_cascade_\ : std_logic;
signal b2v_inst4_pix_count_int_fast_5 : std_logic;
signal b2v_inst4_pix_count_int_fast_6 : std_logic;
signal \b2v_inst.un4_pix_count_intlto6_1_xZ0Z1\ : std_logic;
signal \b2v_inst.un4_pix_count_intlto6_1_xZ0Z0\ : std_logic;
signal \b2v_inst.un4_pix_count_intlto6_dZ0Z_1\ : std_logic;
signal \b2v_inst.un4_pix_count_intlto10_1_0Z0Z_0\ : std_logic;
signal \b2v_inst.un4_pix_count_intlt8_cascade_\ : std_logic;
signal \b2v_inst.un4_pix_count_intlto15_1_aZ0Z0\ : std_logic;
signal \b2v_inst.un4_pix_count_intlt16\ : std_logic;
signal \SYNTHESIZED_WIRE_4_12\ : std_logic;
signal \SYNTHESIZED_WIRE_4_11\ : std_logic;
signal \SYNTHESIZED_WIRE_4_9_rep1\ : std_logic;
signal \b2v_inst1.r_RX_Bytece_0_4_cascade_\ : std_logic;
signal \b2v_inst.un4_pix_count_intlto10_1_d_0_xZ0Z1_cascade_\ : std_logic;
signal \SYNTHESIZED_WIRE_4_0\ : std_logic;
signal \SYNTHESIZED_WIRE_4_3\ : std_logic;
signal \SYNTHESIZED_WIRE_4_1\ : std_logic;
signal \SYNTHESIZED_WIRE_4_2\ : std_logic;
signal \SYNTHESIZED_WIRE_4_6\ : std_logic;
signal \SYNTHESIZED_WIRE_4_5\ : std_logic;
signal \b2v_inst.un4_pix_count_intlto6_d_1_0_cascade_\ : std_logic;
signal \SYNTHESIZED_WIRE_4_10_rep1\ : std_logic;
signal b2v_inst4_pix_count_int_fast_11 : std_logic;
signal b2v_inst4_pix_count_int_fast_12 : std_logic;
signal b2v_inst_un4_pix_count_intlto12_0 : std_logic;
signal \SYNTHESIZED_WIRE_4_10\ : std_logic;
signal \SYNTHESIZED_WIRE_4_9\ : std_logic;
signal \b2v_inst_un4_pix_count_intlto12_0_cascade_\ : std_logic;
signal \SYNTHESIZED_WIRE_4_8\ : std_logic;
signal \N_457_i\ : std_logic;
signal \b2v_inst1.N_48\ : std_logic;
signal \b2v_inst1.N_44_cascade_\ : std_logic;
signal \b2v_inst.N_8\ : std_logic;
signal \b2v_inst1.N_42\ : std_logic;
signal \b2v_inst1.r_SM_Main_d_4\ : std_logic;
signal \b2v_inst1.N_47\ : std_logic;
signal \b2v_inst1.r_SM_Main_d_4_cascade_\ : std_logic;
signal \b2v_inst1.N_51\ : std_logic;
signal \SYNTHESIZED_WIRE_12_9\ : std_logic;
signal \bfn_8_5_0_\ : std_logic;
signal \b2v_inst.un2_dir_mem_1_cry_0\ : std_logic;
signal \b2v_inst.un2_dir_mem_1_cry_1\ : std_logic;
signal \b2v_inst.un2_dir_mem_1_cry_2\ : std_logic;
signal \b2v_inst.un2_dir_mem_1_cry_3\ : std_logic;
signal \b2v_inst.un2_dir_mem_1_cry_4\ : std_logic;
signal \b2v_inst.un2_dir_mem_1_cry_5\ : std_logic;
signal \b2v_inst.un2_dir_mem_1_cry_6\ : std_logic;
signal \b2v_inst.un2_dir_mem_1_cry_7\ : std_logic;
signal \bfn_8_6_0_\ : std_logic;
signal \b2v_inst.un2_dir_mem_1_cry_8\ : std_logic;
signal \b2v_inst.un1_indice_cry_10_THRU_CO\ : std_logic;
signal \b2v_inst.dir_mem_3_RNO_0Z0Z_10\ : std_logic;
signal \b2v_inst.dir_mem_3_RNO_0Z0Z_7\ : std_logic;
signal \b2v_inst.dir_mem_3_RNO_0Z0Z_8\ : std_logic;
signal \b2v_inst.dir_mem_3_RNO_0Z0Z_9\ : std_logic;
signal \b2v_inst.un1_indice_cry_2_c_RNI00LGZ0\ : std_logic;
signal \b2v_inst.indice_RNIJFHBZ0Z_0\ : std_logic;
signal \b2v_inst.un1_indice_cry_5_c_RNI69OGZ0\ : std_logic;
signal \b2v_inst.dir_mem_3_RNO_0Z0Z_6\ : std_logic;
signal \bfn_8_9_0_\ : std_logic;
signal \b2v_inst.un3_dir_mem_cry_0\ : std_logic;
signal \b2v_inst.un3_dir_mem_cry_1\ : std_logic;
signal \b2v_inst.un3_dir_mem_cry_2\ : std_logic;
signal \b2v_inst.un3_dir_mem_cry_3\ : std_logic;
signal \b2v_inst.un3_dir_mem_cry_4\ : std_logic;
signal \b2v_inst.un3_dir_mem_cry_5\ : std_logic;
signal \b2v_inst.un3_dir_mem_cry_6\ : std_logic;
signal \b2v_inst.un3_dir_mem_cry_7\ : std_logic;
signal \bfn_8_10_0_\ : std_logic;
signal \b2v_inst.un3_dir_mem_cry_8\ : std_logic;
signal \b2v_inst.un3_dir_mem_cry_9\ : std_logic;
signal \SYNTHESIZED_WIRE_4_13\ : std_logic;
signal \SYNTHESIZED_WIRE_4_15\ : std_logic;
signal \SYNTHESIZED_WIRE_4_14\ : std_logic;
signal \b2v_inst.state_RNO_25Z0Z_29\ : std_logic;
signal \b2v_inst.g2_1_0\ : std_logic;
signal \b2v_inst.m29_2_cascade_\ : std_logic;
signal \b2v_inst.un4_pix_count_intlto10_1_d_0\ : std_logic;
signal \b2v_inst1.N_96_cascade_\ : std_logic;
signal \b2v_inst.g0_0_i_a4Z0Z_0\ : std_logic;
signal \b2v_inst.g0_0_iZ0Z_2\ : std_logic;
signal \b2v_inst.g2Z0Z_1\ : std_logic;
signal \b2v_inst1.N_58_i_cascade_\ : std_logic;
signal \b2v_inst1.un22_r_clk_count_ac0_3\ : std_logic;
signal \b2v_inst1.r_RX_Bytece_0_6\ : std_logic;
signal \b2v_inst1.r_Clk_CountZ0Z_2\ : std_logic;
signal \b2v_inst1.m16_0_o2_cascade_\ : std_logic;
signal \b2v_inst.g0_1_0_0\ : std_logic;
signal \SYNTHESIZED_WIRE_4_7\ : std_logic;
signal \b2v_inst.un4_pix_count_intlto6_d_1_2\ : std_logic;
signal \SYNTHESIZED_WIRE_4_4\ : std_logic;
signal \b2v_inst.g1_0_0\ : std_logic;
signal \b2v_inst.g1_0_0Z0Z_2\ : std_logic;
signal \b2v_inst.g1_0_a4Z0Z_0\ : std_logic;
signal swit_c_9 : std_logic;
signal \b2v_inst.addr_ram_energia_m0_9\ : std_logic;
signal \b2v_inst1.N_38_cascade_\ : std_logic;
signal \b2v_inst1.r_Bit_IndexZ0Z_2\ : std_logic;
signal \b2v_inst1.N_44\ : std_logic;
signal \b2v_inst1.N_36_cascade_\ : std_logic;
signal \b2v_inst1.r_Bit_IndexZ0Z_1\ : std_logic;
signal \b2v_inst1.r_Bit_IndexZ0Z_0\ : std_logic;
signal \b2v_inst1.N_50\ : std_logic;
signal \b2v_inst1.r_RX_Bytece_0_5\ : std_logic;
signal \N_460_i\ : std_logic;
signal \N_459_i\ : std_logic;
signal \bfn_9_5_0_\ : std_logic;
signal \b2v_inst.un8_dir_mem_2_cry_1\ : std_logic;
signal \b2v_inst.un8_dir_mem_2_cry_2\ : std_logic;
signal \b2v_inst.un8_dir_mem_2_cry_3\ : std_logic;
signal \b2v_inst.un8_dir_mem_2_cry_4\ : std_logic;
signal \b2v_inst.un8_dir_mem_2_cry_5\ : std_logic;
signal \b2v_inst.un8_dir_mem_2_cry_6\ : std_logic;
signal \b2v_inst.un8_dir_mem_2_cry_7\ : std_logic;
signal \b2v_inst.un8_dir_mem_2_cry_8\ : std_logic;
signal \bfn_9_6_0_\ : std_logic;
signal \b2v_inst.un8_dir_mem_2_cry_9\ : std_logic;
signal \b2v_inst.dir_mem_215lt6_0\ : std_logic;
signal leds_c_4 : std_logic;
signal leds_c_5 : std_logic;
signal \b2v_inst.dir_mem_115lt6_0\ : std_logic;
signal \b2v_inst.g0_1_0_cascade_\ : std_logic;
signal \b2v_inst.un7_pix_count_int_0_N_2_THRU_CO\ : std_logic;
signal \b2v_inst.g0_6_cascade_\ : std_logic;
signal \b2v_inst.o2\ : std_logic;
signal \b2v_inst.G_40_i_6_cascade_\ : std_logic;
signal \b2v_inst.state_ns_i_0_a2_11_a2_0_3_3\ : std_logic;
signal \b2v_inst.N_618_5\ : std_logic;
signal \b2v_inst1.N_49\ : std_logic;
signal \b2v_inst1.r_RX_Byte_1_sqmuxa\ : std_logic;
signal \b2v_inst.N_618_3\ : std_logic;
signal \b2v_inst.state_ns_i_0_a2_11_o2_4_0_3_3\ : std_logic;
signal \b2v_inst.un4_pix_count_intlto19_0_0\ : std_logic;
signal \b2v_inst.G_40_i_2\ : std_logic;
signal \b2v_inst.G_40_i_3\ : std_logic;
signal \SYNTHESIZED_WIRE_4_19\ : std_logic;
signal \SYNTHESIZED_WIRE_4_16\ : std_logic;
signal \b2v_inst.N_5\ : std_logic;
signal \b2v_inst.N_430_i_1_cascade_\ : std_logic;
signal \SYNTHESIZED_WIRE_4_18\ : std_logic;
signal \SYNTHESIZED_WIRE_4_17\ : std_logic;
signal \b2v_inst.g1Z0Z_0\ : std_logic;
signal \b2v_inst.pix_count_anterior5\ : std_logic;
signal \b2v_inst.state_ns_0_i_o2_6_23_cascade_\ : std_logic;
signal \b2v_inst.state_ns_0_i_o2_7_23\ : std_logic;
signal \b2v_inst.N_512_cascade_\ : std_logic;
signal \b2v_inst.N_430_tz\ : std_logic;
signal \b2v_inst.g0_4_4_cascade_\ : std_logic;
signal \b2v_inst.g3_0_0\ : std_logic;
signal \b2v_inst.un4_pix_count_intlto18Z0Z_0\ : std_logic;
signal \b2v_inst.g0_0_cascade_\ : std_logic;
signal \b2v_inst.g3_0\ : std_logic;
signal \b2v_inst.g0_4_5\ : std_logic;
signal leds_c_10 : std_logic;
signal leds_c_11 : std_logic;
signal leds_c_7 : std_logic;
signal \b2v_inst.un8_dir_mem_1_cry_2_c_RNI82QCZ0\ : std_logic;
signal \b2v_inst.un8_dir_mem_1_cry_3_c_RNIA5RCZ0\ : std_logic;
signal \b2v_inst.un8_dir_mem_1_cry_5_c_RNIEBTCZ0\ : std_logic;
signal \b2v_inst.dir_mem_1_RNO_0Z0Z_6\ : std_logic;
signal \b2v_inst.dir_mem_215lt7\ : std_logic;
signal \b2v_inst.dir_mem_115lt7\ : std_logic;
signal \b2v_inst.dir_mem_1_RNO_0Z0Z_10\ : std_logic;
signal \b2v_inst.dir_mem_115lt11_cascade_\ : std_logic;
signal \b2v_inst.dir_mem_115lto7\ : std_logic;
signal \b2v_inst.dir_mem_1_RNO_0Z0Z_7\ : std_logic;
signal \b2v_inst.un8_dir_mem_1_cry_7_c_RNIIHVCZ0\ : std_logic;
signal \b2v_inst.dir_mem_1_RNO_0Z0Z_8\ : std_logic;
signal \b2v_inst.un8_dir_mem_1_cry_8_c_RNIKK0DZ0\ : std_logic;
signal \b2v_inst.dir_mem_1_RNO_0Z0Z_9\ : std_logic;
signal \b2v_inst.un8_dir_mem_1_cry_4_c_RNIC8SCZ0\ : std_logic;
signal \b2v_inst.dir_mem_1_RNO_0Z0Z_5\ : std_logic;
signal \b2v_inst.dir_mem_1Z0Z_6\ : std_logic;
signal \b2v_inst.dir_mem_3Z0Z_6\ : std_logic;
signal \b2v_inst.dir_memZ0Z_7\ : std_logic;
signal \b2v_inst.N_450_i_1_cascade_\ : std_logic;
signal \b2v_inst.dir_memZ0Z_10\ : std_logic;
signal \b2v_inst.dir_mem_1Z0Z_5\ : std_logic;
signal \b2v_inst.dir_mem_3Z0Z_5\ : std_logic;
signal \SYNTHESIZED_WIRE_1_5\ : std_logic;
signal \b2v_inst.dir_memZ0Z_4\ : std_logic;
signal \b2v_inst.addr_ram_iv_i_0_4_cascade_\ : std_logic;
signal \indice_RNIN3333_4\ : std_logic;
signal \b2v_inst.dir_mem_1Z0Z_4\ : std_logic;
signal \b2v_inst.addr_ram_iv_i_1_4\ : std_logic;
signal \b2v_inst.un1_indice_cry_3_c_RNI23MGZ0\ : std_logic;
signal \b2v_inst.dir_mem_316lto11_0\ : std_logic;
signal \b2v_inst.dir_mem_316lt11\ : std_logic;
signal \b2v_inst.dir_mem_3Z0Z_4\ : std_logic;
signal \b2v_inst.N_362_i\ : std_logic;
signal \b2v_inst.state_ns_0_i_a2_0_0_23\ : std_logic;
signal \b2v_inst.state_ns_i_0_a2_11_o2_4_0_6_1_3_cascade_\ : std_logic;
signal \b2v_inst.state_ns_i_0_a2_11_o2_4_0_1_3\ : std_logic;
signal \b2v_inst.N_11\ : std_logic;
signal \b2v_inst.N_4_i_i_1_cascade_\ : std_logic;
signal \b2v_inst.g3_i_1\ : std_logic;
signal swit_c_8 : std_logic;
signal \b2v_inst.addr_ram_energia_m0_8\ : std_logic;
signal \b2v_inst.state_ns_i_0_a2_11_o2_4_0_5_3\ : std_logic;
signal \b2v_inst.state_RNO_2Z0Z_29\ : std_logic;
signal \b2v_inst.state_ns_i_0_a2_11_o2_4_0_7_3_cascade_\ : std_logic;
signal \b2v_inst.state_RNO_1Z0Z_29\ : std_logic;
signal \b2v_inst.dir_energia_RNO_0Z0Z_0\ : std_logic;
signal swit_c_6 : std_logic;
signal \b2v_inst.addr_ram_energia_m0_6_cascade_\ : std_logic;
signal \SYNTHESIZED_WIRE_12_6\ : std_logic;
signal swit_c_7 : std_logic;
signal \b2v_inst.addr_ram_energia_m0_7\ : std_logic;
signal leds_c_12 : std_logic;
signal \b2v_inst.un1_indice_cry_4_c_RNI46NGZ0\ : std_logic;
signal \b2v_inst.un1_indice_cry_8_c_RNICIRGZ0\ : std_logic;
signal \b2v_inst.dir_mem_316lto7\ : std_logic;
signal \b2v_inst.un8_dir_mem_2_cry_1_c_RNI88LLZ0\ : std_logic;
signal \b2v_inst.un8_dir_mem_2_cry_2_c_RNIABMLZ0\ : std_logic;
signal \b2v_inst.dir_mem_2Z0Z_4\ : std_logic;
signal \b2v_inst.un8_dir_mem_2_cry_3_c_RNICENLZ0\ : std_logic;
signal \b2v_inst.un8_dir_mem_2_cry_4_c_RNIEHOLZ0\ : std_logic;
signal \b2v_inst.un8_dir_mem_1_cry_10_THRU_CO\ : std_logic;
signal \b2v_inst.un8_dir_mem_1_cry_9_c_RNITCOLZ0\ : std_logic;
signal \b2v_inst.dir_mem_1Z0Z_8\ : std_logic;
signal \b2v_inst.dir_mem_3Z0Z_8\ : std_logic;
signal \b2v_inst.dir_mem_3Z0Z_1\ : std_logic;
signal \b2v_inst.dir_memZ0Z_1\ : std_logic;
signal \b2v_inst.dir_mem_2Z0Z_1\ : std_logic;
signal \b2v_inst.un8_dir_mem_1_cry_0_c_RNI4SNCZ0\ : std_logic;
signal \b2v_inst.dir_mem_1Z0Z_1\ : std_logic;
signal \b2v_inst.dir_mem_115lt11\ : std_logic;
signal \b2v_inst.indice_RNILHHBZ0Z_2\ : std_logic;
signal \b2v_inst.dir_mem_115lto11_0\ : std_logic;
signal \b2v_inst.un8_dir_mem_1_cry_1_c_RNI6VOCZ0\ : std_logic;
signal \b2v_inst.N_363_i\ : std_logic;
signal \b2v_inst.dir_mem_2Z0Z_6\ : std_logic;
signal \b2v_inst.N_489_cascade_\ : std_logic;
signal \b2v_inst.dir_mem_1Z0Z_7\ : std_logic;
signal \b2v_inst.dir_mem_3Z0Z_7\ : std_logic;
signal \b2v_inst.N_488_cascade_\ : std_logic;
signal \b2v_inst.addr_ram_iv_i_0_0_7\ : std_logic;
signal \b2v_inst.addr_ram_iv_i_0_1_7_cascade_\ : std_logic;
signal \indice_RNI6J333_7\ : std_logic;
signal \b2v_inst.state_RNO_0Z0Z_29\ : std_logic;
signal \b2v_inst.dir_mem_1Z0Z_0\ : std_logic;
signal \b2v_inst.dir_mem_3Z0Z_0\ : std_logic;
signal \b2v_inst.dir_mem_2Z0Z_3\ : std_logic;
signal \b2v_inst.dir_memZ0Z_3\ : std_logic;
signal \b2v_inst.addr_ram_iv_i_0_0_3_cascade_\ : std_logic;
signal \indice_RNIIU233_3\ : std_logic;
signal \b2v_inst.dir_mem_3Z0Z_3\ : std_logic;
signal \b2v_inst.dir_mem_1Z0Z_3\ : std_logic;
signal \b2v_inst.addr_ram_iv_i_0_1_3\ : std_logic;
signal \b2v_inst.dir_memZ0Z_0\ : std_logic;
signal \b2v_inst.N_618_6\ : std_logic;
signal \b2v_inst.N_514_cascade_\ : std_logic;
signal \N_116_i\ : std_logic;
signal \b2v_inst.stateZ0Z_16\ : std_logic;
signal \N_548_i\ : std_logic;
signal \b2v_inst.stateZ0Z_0\ : std_logic;
signal \b2v_inst.N_692_cascade_\ : std_logic;
signal \b2v_inst.N_477\ : std_logic;
signal swit_c_1 : std_logic;
signal \b2v_inst.N_494_cascade_\ : std_logic;
signal \b2v_inst.addr_ram_energia_m0_1\ : std_logic;
signal \SYNTHESIZED_WIRE_12_10\ : std_logic;
signal swit_c_2 : std_logic;
signal \b2v_inst.addr_ram_energia_m0_2_cascade_\ : std_logic;
signal \SYNTHESIZED_WIRE_12_2\ : std_logic;
signal swit_c_5 : std_logic;
signal \b2v_inst.addr_ram_energia_m0_5_cascade_\ : std_logic;
signal \SYNTHESIZED_WIRE_12_5\ : std_logic;
signal swit_c_10 : std_logic;
signal \b2v_inst.addr_ram_energia_m0_10\ : std_logic;
signal swit_c_3 : std_logic;
signal \b2v_inst.addr_ram_energia_m0_3_cascade_\ : std_logic;
signal \SYNTHESIZED_WIRE_12_3\ : std_logic;
signal leds_c_6 : std_logic;
signal swit_c_0 : std_logic;
signal \b2v_inst.addr_ram_energia_m0_0\ : std_logic;
signal \N_120_i\ : std_logic;
signal \b2v_inst.N_432_1_cascade_\ : std_logic;
signal \b2v_inst.un1_indice_cry_9_c_RNILAJPZ0\ : std_logic;
signal \b2v_inst.un1_indice_cry_7_c_RNIAFQGZ0\ : std_logic;
signal \b2v_inst.dir_mem_2Z0Z_0\ : std_logic;
signal \b2v_inst.un8_dir_mem_2_cry_9_THRU_CO\ : std_logic;
signal \b2v_inst.un8_dir_mem_2_cry_8_c_RNITIJEZ0\ : std_logic;
signal \b2v_inst.dir_mem_2Z0Z_10\ : std_logic;
signal \b2v_inst.dir_mem_215lto7\ : std_logic;
signal \b2v_inst.dir_mem_2Z0Z_7\ : std_logic;
signal \b2v_inst.un8_dir_mem_2_cry_6_c_RNIINQZ0Z5\ : std_logic;
signal \b2v_inst.dir_mem_2Z0Z_8\ : std_logic;
signal \b2v_inst.un8_dir_mem_2_cry_7_c_RNIKQRZ0Z5\ : std_logic;
signal \b2v_inst.dir_mem_215lto11_0\ : std_logic;
signal \b2v_inst.dir_mem_215lt11\ : std_logic;
signal \b2v_inst.N_463_i\ : std_logic;
signal \b2v_inst.indice_4_i_a2_0_7_3_1\ : std_logic;
signal \b2v_inst.N_432_1_tz\ : std_logic;
signal \N_556_i\ : std_logic;
signal \b2v_inst.indice_4_i_a2_0_7_2_1\ : std_logic;
signal \N_117_i\ : std_logic;
signal \b2v_inst.dir_mem_1Z0Z_9\ : std_logic;
signal \b2v_inst.dir_mem_3Z0Z_9\ : std_logic;
signal \N_554_i\ : std_logic;
signal \b2v_inst.dir_mem_2Z0Z_2\ : std_logic;
signal \b2v_inst.dir_memZ0Z_2\ : std_logic;
signal \b2v_inst.dir_mem_2Z0Z_9\ : std_logic;
signal \b2v_inst.dir_mem_1Z0Z_2\ : std_logic;
signal \b2v_inst.dir_mem_3Z0Z_2\ : std_logic;
signal \b2v_inst.N_829_cascade_\ : std_logic;
signal \b2v_inst.N_829\ : std_logic;
signal \b2v_inst.un1_state_23_i_a2_0_a2_0_a2_0_cascade_\ : std_logic;
signal \b2v_inst.stateZ0Z_22\ : std_logic;
signal \b2v_inst.stateZ0Z_26\ : std_logic;
signal \b2v_inst.un2_cuentalto10_i_a2_6\ : std_logic;
signal \b2v_inst1.m16_0_o2\ : std_logic;
signal \b2v_inst1.m16_0_a3_0_cascade_\ : std_logic;
signal \b2v_inst1.N_119\ : std_logic;
signal \b2v_inst1.r_Clk_Count_6_iv_0_a3_1_1_1_cascade_\ : std_logic;
signal \b2v_inst1.N_43\ : std_logic;
signal \b2v_inst1.r_Clk_Count_6_iv_0_0_1_cascade_\ : std_logic;
signal \b2v_inst1.r_Clk_CountZ0Z_0\ : std_logic;
signal \b2v_inst1.r_Clk_CountZ0Z_1\ : std_logic;
signal \b2v_inst.N_653_cascade_\ : std_logic;
signal \b2v_inst.stateZ0Z_17\ : std_logic;
signal \b2v_inst.state_ns_i_a2_1_15\ : std_logic;
signal \b2v_inst.cuenta_RNIKUJVZ0Z_0_cascade_\ : std_logic;
signal \b2v_inst.un20_cuentalto10_5_cascade_\ : std_logic;
signal \b2v_inst.un20_cuentalto10_sx\ : std_logic;
signal \b2v_inst.un20_cuentalto10_sx_cascade_\ : std_logic;
signal \b2v_inst.state18_li_0_cascade_\ : std_logic;
signal \N_130_i\ : std_logic;
signal \b2v_inst.N_512\ : std_logic;
signal \b2v_inst.stateZ0Z_30\ : std_logic;
signal \b2v_inst.N_828_cascade_\ : std_logic;
signal \N_552_i\ : std_logic;
signal \b2v_inst.state_ns_0_i_o2_8_23\ : std_logic;
signal \N_550_i\ : std_logic;
signal \b2v_inst.state_fastZ0Z_32\ : std_logic;
signal \b2v_inst.stateZ0Z_5\ : std_logic;
signal \b2v_inst.addr_ram_energia_ss0_0_i_o2_i_o2_0\ : std_logic;
signal \b2v_inst.dir_mem_RNO_0Z0Z_6\ : std_logic;
signal \b2v_inst.dir_memZ0Z_6\ : std_logic;
signal \b2v_inst.dir_mem_RNO_0Z0Z_8\ : std_logic;
signal \b2v_inst.dir_memZ0Z_8\ : std_logic;
signal \b2v_inst.dir_mem_RNO_0Z0Z_9\ : std_logic;
signal \b2v_inst.dir_memZ0Z_9\ : std_logic;
signal swit_c_4 : std_logic;
signal \b2v_inst.N_494\ : std_logic;
signal \b2v_inst.N_247\ : std_logic;
signal \b2v_inst.addr_ram_energia_m0_4_cascade_\ : std_logic;
signal \SYNTHESIZED_WIRE_12_4\ : std_logic;
signal uart_rx_i_c : std_logic;
signal \b2v_inst1.r_RX_Data_RZ0\ : std_logic;
signal \b2v_inst.un9_indice_0_a2_2\ : std_logic;
signal \b2v_inst.un9_indice_0_a2_3\ : std_logic;
signal \b2v_inst.dir_mem_RNO_0Z0Z_5\ : std_logic;
signal \b2v_inst.un9_indice_0_a2_2_cascade_\ : std_logic;
signal \b2v_inst.stateZ0Z_28\ : std_logic;
signal \b2v_inst.N_432_1\ : std_logic;
signal \bfn_13_6_0_\ : std_logic;
signal \b2v_inst.N_442_i\ : std_logic;
signal \b2v_inst.un2_dir_mem_2_cry_0_THRU_CO\ : std_logic;
signal \b2v_inst.un2_dir_mem_2_cry_0\ : std_logic;
signal \b2v_inst.dir_mem_2_RNO_0Z0Z_2\ : std_logic;
signal \b2v_inst.un2_dir_mem_2_cry_1\ : std_logic;
signal \b2v_inst.dir_mem_2_RNO_0Z0Z_3\ : std_logic;
signal \b2v_inst.un2_dir_mem_2_cry_2\ : std_logic;
signal \b2v_inst.dir_mem_2_RNO_0Z0Z_4\ : std_logic;
signal \b2v_inst.un2_dir_mem_2_cry_3\ : std_logic;
signal \b2v_inst.dir_mem_2_RNO_0Z0Z_5\ : std_logic;
signal \b2v_inst.un2_dir_mem_2_cry_4\ : std_logic;
signal \b2v_inst.dir_mem_2_RNO_0Z0Z_6\ : std_logic;
signal \b2v_inst.un2_dir_mem_2_cry_5\ : std_logic;
signal \b2v_inst.dir_mem_2_RNO_0Z0Z_7\ : std_logic;
signal \b2v_inst.un2_dir_mem_2_cry_6\ : std_logic;
signal \b2v_inst.un2_dir_mem_2_cry_7\ : std_logic;
signal \b2v_inst.dir_mem_2_RNO_0Z0Z_8\ : std_logic;
signal \bfn_13_7_0_\ : std_logic;
signal \b2v_inst.dir_mem_2_RNO_0Z0Z_9\ : std_logic;
signal \b2v_inst.un2_dir_mem_2_cry_8\ : std_logic;
signal \b2v_inst.un2_dir_mem_2_cry_9\ : std_logic;
signal \b2v_inst.dir_mem_2_RNO_0Z0Z_10\ : std_logic;
signal \b2v_inst1.r_SM_MainZ0Z_1\ : std_logic;
signal \b2v_inst1.r_RX_DataZ0\ : std_logic;
signal \b2v_inst1.r_SM_MainZ0Z_2\ : std_logic;
signal \b2v_inst1.m13_i_2\ : std_logic;
signal \b2v_inst1.N_95_cascade_\ : std_logic;
signal \b2v_inst1.N_96\ : std_logic;
signal \b2v_inst1.r_SM_MainZ0Z_0\ : std_logic;
signal \b2v_inst.dir_memZ0Z_5\ : std_logic;
signal \b2v_inst.N_450_i_1\ : std_logic;
signal \b2v_inst.dir_mem_2Z0Z_5\ : std_logic;
signal \b2v_inst.N_489\ : std_logic;
signal \b2v_inst9.data_to_send_10_0_0_0_5_cascade_\ : std_logic;
signal \b2v_inst9.data_to_sendZ0Z_5\ : std_logic;
signal \b2v_inst9.data_to_send_10_0_0_0_3_cascade_\ : std_logic;
signal \b2v_inst9.data_to_sendZ0Z_6\ : std_logic;
signal \b2v_inst.un1_data_a_escribir_0_sqmuxa_3_i_i_a2_0\ : std_logic;
signal \b2v_inst.N_655_cascade_\ : std_logic;
signal \b2v_inst.state18_li_0\ : std_logic;
signal \b2v_inst.cuenta_RNIR03AZ0Z_1\ : std_logic;
signal \b2v_inst.cuentaZ0Z_0\ : std_logic;
signal \b2v_inst.cuentaZ0Z_1\ : std_logic;
signal \bfn_13_12_0_\ : std_logic;
signal \b2v_inst.cuentaZ0Z_2\ : std_logic;
signal \b2v_inst.un4_cuenta_cry_1_c_RNI9VZ0Z48\ : std_logic;
signal \b2v_inst.un4_cuenta_cry_1\ : std_logic;
signal \b2v_inst.cuentaZ0Z_3\ : std_logic;
signal \b2v_inst.un4_cuenta_cry_2_c_RNIBZ0Z268\ : std_logic;
signal \b2v_inst.un4_cuenta_cry_2\ : std_logic;
signal \b2v_inst.cuentaZ0Z_4\ : std_logic;
signal \b2v_inst.un4_cuenta_cry_3_c_RNIDZ0Z578\ : std_logic;
signal \b2v_inst.un4_cuenta_cry_3\ : std_logic;
signal \b2v_inst.un4_cuenta_cry_4\ : std_logic;
signal \b2v_inst.cuentaZ0Z_6\ : std_logic;
signal \b2v_inst.un4_cuenta_cry_5_c_RNIHBZ0Z98\ : std_logic;
signal \b2v_inst.un4_cuenta_cry_5\ : std_logic;
signal \b2v_inst.cuentaZ0Z_7\ : std_logic;
signal \b2v_inst.un4_cuenta_cry_6_c_RNIJEAZ0Z8\ : std_logic;
signal \b2v_inst.un4_cuenta_cry_6\ : std_logic;
signal \b2v_inst.cuentaZ0Z_8\ : std_logic;
signal \b2v_inst.un4_cuenta_cry_7_c_RNILHBZ0Z8\ : std_logic;
signal \b2v_inst.un4_cuenta_cry_7\ : std_logic;
signal \b2v_inst.un4_cuenta_cry_8\ : std_logic;
signal \b2v_inst.cuentaZ0Z_9\ : std_logic;
signal \b2v_inst.un4_cuenta_cry_8_c_RNINKCZ0Z8\ : std_logic;
signal \bfn_13_13_0_\ : std_logic;
signal \b2v_inst.un4_cuenta_cry_9\ : std_logic;
signal \N_458_i\ : std_logic;
signal b2v_inst_state_4 : std_logic;
signal b2v_inst_state_8 : std_logic;
signal leds_c_0 : std_logic;
signal leds_c_1 : std_logic;
signal leds_c_13 : std_logic;
signal leds_c_2 : std_logic;
signal leds_c_3 : std_logic;
signal \N_546_i\ : std_logic;
signal \bfn_13_16_0_\ : std_logic;
signal \b2v_inst.dir_energia_s_1\ : std_logic;
signal \b2v_inst.dir_energia_cry_0\ : std_logic;
signal \b2v_inst.dir_energia_s_2\ : std_logic;
signal \b2v_inst.dir_energia_cry_1\ : std_logic;
signal \b2v_inst.dir_energia_s_3\ : std_logic;
signal \b2v_inst.dir_energia_cry_2\ : std_logic;
signal \b2v_inst.dir_energia_s_4\ : std_logic;
signal \b2v_inst.dir_energia_cry_3\ : std_logic;
signal \b2v_inst.dir_energia_s_5\ : std_logic;
signal \b2v_inst.dir_energia_cry_4\ : std_logic;
signal \b2v_inst.dir_energia_s_6\ : std_logic;
signal \b2v_inst.dir_energia_cry_5\ : std_logic;
signal \b2v_inst.dir_energia_s_7\ : std_logic;
signal \b2v_inst.dir_energia_cry_6\ : std_logic;
signal \b2v_inst.dir_energia_cry_7\ : std_logic;
signal \b2v_inst.dir_energia_s_8\ : std_logic;
signal \bfn_13_17_0_\ : std_logic;
signal \b2v_inst.dir_energia_s_9\ : std_logic;
signal \b2v_inst.dir_energia_cry_8\ : std_logic;
signal \b2v_inst.dir_energia_s_10\ : std_logic;
signal \b2v_inst.dir_energia_cry_9\ : std_logic;
signal \b2v_inst.stateZ0Z_19\ : std_logic;
signal \b2v_inst.N_352_0\ : std_logic;
signal \b2v_inst.dir_energia_cry_10\ : std_logic;
signal \b2v_inst.dir_energiaZ0Z_11\ : std_logic;
signal \b2v_inst.N_430_i\ : std_logic;
signal \b2v_inst.N_648_5\ : std_logic;
signal \b2v_inst.un9_indice_0_a2_5_1\ : std_logic;
signal \b2v_inst.un4_cuenta_cry_9_c_RNI01TZ0Z9\ : std_logic;
signal \b2v_inst.cuentaZ0Z_10\ : std_logic;
signal \b2v_inst.N_655\ : std_logic;
signal \b2v_inst.un4_cuenta_cry_4_c_RNIFZ0Z888\ : std_logic;
signal \b2v_inst.cuentaZ0Z_5\ : std_logic;
signal \b2v_inst.N_547_i_0\ : std_logic;
signal \b2v_inst9.data_to_send_10_0_0_0_4\ : std_logic;
signal \b2v_inst9.data_to_sendZ0Z_4\ : std_logic;
signal \b2v_inst9.data_to_send_10_0_0_1_4\ : std_logic;
signal \b2v_inst9.data_to_send_10_0_0_1_5\ : std_logic;
signal \b2v_inst9.fsm_state_ns_i_i_0_a2_2_2Z0Z_0\ : std_logic;
signal \b2v_inst9.N_583_cascade_\ : std_logic;
signal reset_c_i : std_logic;
signal \b2v_inst9.un2_n_fsm_state_0_sqmuxa_2_0_i_cascade_\ : std_logic;
signal \b2v_inst9.data_to_send_10_0_0_0_6\ : std_logic;
signal \b2v_inst9.data_to_send_10_0_0_0_7_cascade_\ : std_logic;
signal \b2v_inst9.data_to_sendZ0Z_7\ : std_logic;
signal \b2v_inst9.data_to_send_10_0_0_2_0\ : std_logic;
signal \b2v_inst9.data_to_send_10_0_0_1_0\ : std_logic;
signal \b2v_inst9.N_738_cascade_\ : std_logic;
signal \b2v_inst9.data_to_send_10_0_0_2_1\ : std_logic;
signal \b2v_inst9.data_to_sendZ0Z_1\ : std_logic;
signal \N_478_cascade_\ : std_logic;
signal \b2v_inst9.data_to_send_10_0_0_0_0\ : std_logic;
signal b2v_inst_state_15 : std_logic;
signal \b2v_inst9.N_832_cascade_\ : std_logic;
signal \b2v_inst9.data_to_send_10_0_0_0_1\ : std_logic;
signal \b2v_inst9.data_to_send_10_0_0_1_1\ : std_logic;
signal \b2v_inst9.data_to_send_10_0_0_2_2_cascade_\ : std_logic;
signal \b2v_inst9.data_to_sendZ0Z_2\ : std_logic;
signal \b2v_inst9.un2_n_fsm_state_0_sqmuxa_2_0_i_0\ : std_logic;
signal \b2v_inst9.N_740\ : std_logic;
signal \b2v_inst9.data_to_send_10_0_0_1_2\ : std_logic;
signal \b2v_inst9.N_738\ : std_logic;
signal \b2v_inst9.N_741\ : std_logic;
signal \b2v_inst9.data_to_send_10_0_0_1_3\ : std_logic;
signal b2v_inst_energia_temp_0 : std_logic;
signal \b2v_inst.un14_data_ram_energia_o_axb_0\ : std_logic;
signal \bfn_14_14_0_\ : std_logic;
signal b2v_inst_energia_temp_1 : std_logic;
signal \b2v_inst.un14_data_ram_energia_o_cry_0_c_RNIEI4MZ0\ : std_logic;
signal \b2v_inst.un14_data_ram_energia_o_cry_0\ : std_logic;
signal b2v_inst_energia_temp_2 : std_logic;
signal \b2v_inst.un14_data_ram_energia_o_cry_1_c_RNIHM5MZ0\ : std_logic;
signal \b2v_inst.un14_data_ram_energia_o_cry_1\ : std_logic;
signal b2v_inst_energia_temp_3 : std_logic;
signal \b2v_inst.un14_data_ram_energia_o_cry_2_c_RNIKQ6MZ0\ : std_logic;
signal \b2v_inst.un14_data_ram_energia_o_cry_2\ : std_logic;
signal \b2v_inst.pix_data_regZ0Z_4\ : std_logic;
signal b2v_inst_energia_temp_4 : std_logic;
signal \b2v_inst.un14_data_ram_energia_o_cry_3_c_RNINU7MZ0\ : std_logic;
signal \b2v_inst.un14_data_ram_energia_o_cry_3\ : std_logic;
signal b2v_inst_energia_temp_5 : std_logic;
signal \b2v_inst.un14_data_ram_energia_o_cry_4_c_RNIQ29MZ0\ : std_logic;
signal \b2v_inst.un14_data_ram_energia_o_cry_4\ : std_logic;
signal b2v_inst_energia_temp_6 : std_logic;
signal \b2v_inst.un14_data_ram_energia_o_cry_5_c_RNIT6AMZ0\ : std_logic;
signal \b2v_inst.un14_data_ram_energia_o_cry_5\ : std_logic;
signal b2v_inst_energia_temp_7 : std_logic;
signal \b2v_inst.un14_data_ram_energia_o_cry_6_c_RNI0BBMZ0\ : std_logic;
signal \b2v_inst.un14_data_ram_energia_o_cry_6\ : std_logic;
signal \b2v_inst.un14_data_ram_energia_o_cry_7\ : std_logic;
signal \b2v_inst.un14_data_ram_energia_o_cry_7_c_RNIN84CZ0\ : std_logic;
signal \bfn_14_15_0_\ : std_logic;
signal \b2v_inst.un14_data_ram_energia_o_cry_8_c_RNIPB5CZ0\ : std_logic;
signal \b2v_inst.un14_data_ram_energia_o_cry_8\ : std_logic;
signal b2v_inst_energia_temp_10 : std_logic;
signal \b2v_inst.un14_data_ram_energia_o_cry_9\ : std_logic;
signal b2v_inst_energia_temp_11 : std_logic;
signal \SYNTHESIZED_WIRE_13_11\ : std_logic;
signal \b2v_inst.un14_data_ram_energia_o_cry_10\ : std_logic;
signal b2v_inst_energia_temp_12 : std_logic;
signal \SYNTHESIZED_WIRE_13_12\ : std_logic;
signal \b2v_inst.un14_data_ram_energia_o_cry_11\ : std_logic;
signal b2v_inst_energia_temp_13 : std_logic;
signal \b2v_inst.un14_data_ram_energia_o_cry_12\ : std_logic;
signal \SYNTHESIZED_WIRE_13_13\ : std_logic;
signal leds_c_8 : std_logic;
signal b2v_inst_energia_temp_8 : std_logic;
signal \b2v_inst.un14_data_ram_energia_o_cry_9_c_RNI28GBZ0\ : std_logic;
signal \N_461_i\ : std_logic;
signal \bfn_15_8_0_\ : std_logic;
signal \b2v_inst.data_a_escribir11_0\ : std_logic;
signal \b2v_inst.data_a_escribir11_2_and\ : std_logic;
signal \b2v_inst.data_a_escribir11_1\ : std_logic;
signal \b2v_inst.data_a_escribir11_2\ : std_logic;
signal \b2v_inst.data_a_escribir11_4_and\ : std_logic;
signal \b2v_inst.data_a_escribir11_3\ : std_logic;
signal \b2v_inst.data_a_escribir11_4\ : std_logic;
signal \b2v_inst.data_a_escribir11_5\ : std_logic;
signal \b2v_inst.data_a_escribir11_6\ : std_logic;
signal \b2v_inst.data_a_escribir11_7\ : std_logic;
signal \bfn_15_9_0_\ : std_logic;
signal \b2v_inst.data_a_escribir11_8\ : std_logic;
signal \b2v_inst.data_a_escribir11_9\ : std_logic;
signal \b2v_inst.data_a_escribir12\ : std_logic;
signal \b2v_inst.data_a_escribir11_9_and\ : std_logic;
signal \b2v_inst.data_a_escribir11_8_and\ : std_logic;
signal \b2v_inst.dir_mem_1Z0Z_10\ : std_logic;
signal \b2v_inst.N_490\ : std_logic;
signal \b2v_inst.dir_mem_3Z0Z_10\ : std_logic;
signal \b2v_inst.N_488\ : std_logic;
signal \bfn_15_10_0_\ : std_logic;
signal \b2v_inst.eventos_cry_0\ : std_logic;
signal \b2v_inst.eventos_cry_1\ : std_logic;
signal \b2v_inst.eventos_cry_2\ : std_logic;
signal \b2v_inst.eventos_cry_3\ : std_logic;
signal \b2v_inst.eventos_cry_4\ : std_logic;
signal \b2v_inst.eventos_cry_5\ : std_logic;
signal \b2v_inst.eventos_cry_6\ : std_logic;
signal \b2v_inst.eventos_cry_7\ : std_logic;
signal \bfn_15_11_0_\ : std_logic;
signal \b2v_inst.eventos_cry_8\ : std_logic;
signal \b2v_inst.eventos_cry_9\ : std_logic;
signal \b2v_inst.state_ns_a3_i_0_a2_5_1\ : std_logic;
signal \b2v_inst.state_ns_a3_i_0_a2_4_1_cascade_\ : std_logic;
signal \b2v_inst.stateZ0Z_31\ : std_logic;
signal b2v_inst_state_7 : std_logic;
signal b2v_inst_state_1 : std_logic;
signal b2v_inst_state_2 : std_logic;
signal \b2v_inst.stateZ0Z_11\ : std_logic;
signal \b2v_inst.stateZ0Z_32\ : std_logic;
signal b2v_inst_state_14 : std_logic;
signal \b2v_inst.state_ns_a3_i_0_a2_6_1\ : std_logic;
signal \b2v_inst9.fsm_state_ns_i_0_i_0_1_cascade_\ : std_logic;
signal \b2v_inst9.N_832\ : std_logic;
signal \b2v_inst9.data_to_sendZ0Z_3\ : std_logic;
signal \b2v_inst9.data_to_send_10_0_0_0_2\ : std_logic;
signal b2v_inst_state_12 : std_logic;
signal b2v_inst_state_13 : std_logic;
signal \b2v_inst9.N_739\ : std_logic;
signal \b2v_inst.pix_data_regZ0Z_0\ : std_logic;
signal \b2v_inst.pix_data_regZ0Z_1\ : std_logic;
signal \b2v_inst.pix_data_regZ0Z_2\ : std_logic;
signal \b2v_inst.pix_data_regZ0Z_5\ : std_logic;
signal \b2v_inst.pix_data_regZ0Z_6\ : std_logic;
signal \b2v_inst.pix_data_regZ0Z_7\ : std_logic;
signal \b2v_inst9.N_583\ : std_logic;
signal leds_c_9 : std_logic;
signal b2v_inst_energia_temp_9 : std_logic;
signal \b2v_inst.N_577_i\ : std_logic;
signal \b2v_inst9.data_to_sendZ0Z_0\ : std_logic;
signal uart_tx_o_c : std_logic;
signal \b2v_inst.reg_ancho_1_i_0\ : std_logic;
signal \bfn_16_6_0_\ : std_logic;
signal \b2v_inst.reg_ancho_1_i_1\ : std_logic;
signal \b2v_inst.un2_valor_max1_cry_0\ : std_logic;
signal \b2v_inst.reg_ancho_1_i_2\ : std_logic;
signal \b2v_inst.un2_valor_max1_cry_1\ : std_logic;
signal \b2v_inst.reg_ancho_1_i_3\ : std_logic;
signal \b2v_inst.un2_valor_max1_cry_2\ : std_logic;
signal \b2v_inst.reg_ancho_1_i_4\ : std_logic;
signal \b2v_inst.un2_valor_max1_cry_3\ : std_logic;
signal \b2v_inst.reg_ancho_1_i_5\ : std_logic;
signal \b2v_inst.un2_valor_max1_cry_4\ : std_logic;
signal \b2v_inst.reg_ancho_1_i_6\ : std_logic;
signal \b2v_inst.un2_valor_max1_cry_5\ : std_logic;
signal \b2v_inst.reg_ancho_1_i_7\ : std_logic;
signal \b2v_inst.un2_valor_max1_cry_6\ : std_logic;
signal \b2v_inst.un2_valor_max1_cry_7\ : std_logic;
signal \b2v_inst.reg_ancho_1_i_8\ : std_logic;
signal \bfn_16_7_0_\ : std_logic;
signal \b2v_inst.reg_ancho_1_i_9\ : std_logic;
signal \b2v_inst.un2_valor_max1_cry_8\ : std_logic;
signal \b2v_inst.reg_ancho_1_i_10\ : std_logic;
signal \b2v_inst.un2_valor_max1_cry_9\ : std_logic;
signal \b2v_inst.un2_valor_max1\ : std_logic;
signal \b2v_inst.ignorar_anchoZ0Z_1\ : std_logic;
signal \b2v_inst.stateZ0Z_25\ : std_logic;
signal \b2v_inst.data_a_escribir11_0_and\ : std_logic;
signal \b2v_inst.eventosZ0Z_0\ : std_logic;
signal \b2v_inst.data_a_escribir_RNO_2Z0Z_0_cascade_\ : std_logic;
signal \b2v_inst.un1_reg_anterior_0_i_1_0_cascade_\ : std_logic;
signal \b2v_inst.eventosZ0Z_1\ : std_logic;
signal \b2v_inst.data_a_escribir_RNO_2Z0Z_1_cascade_\ : std_logic;
signal \b2v_inst.un1_reg_anterior_0_i_1_1_cascade_\ : std_logic;
signal \b2v_inst.eventosZ0Z_10\ : std_logic;
signal \b2v_inst.N_269\ : std_logic;
signal \b2v_inst.un1_reg_anterior_iv_0_0_10_cascade_\ : std_logic;
signal \b2v_inst.eventosZ0Z_6\ : std_logic;
signal \b2v_inst.un1_reg_anterior_iv_0_0_6_cascade_\ : std_logic;
signal \b2v_inst.N_272\ : std_logic;
signal \b2v_inst.data_a_escribir_1_sqmuxa\ : std_logic;
signal \b2v_inst.data_a_escribir11_1_and\ : std_logic;
signal \b2v_inst.eventosZ0Z_4\ : std_logic;
signal \b2v_inst.un1_reg_anterior_iv_0_0_4_cascade_\ : std_logic;
signal \b2v_inst.un1_reg_anterior_iv_0_1_4_cascade_\ : std_logic;
signal \b2v_inst.N_274\ : std_logic;
signal \b2v_inst.N_268\ : std_logic;
signal \b2v_inst.un1_reg_anterior_iv_0_1_10\ : std_logic;
signal \SYNTHESIZED_WIRE_10_3\ : std_logic;
signal \SYNTHESIZED_WIRE_10_4\ : std_logic;
signal \SYNTHESIZED_WIRE_10_6\ : std_logic;
signal \SYNTHESIZED_WIRE_10_7\ : std_logic;
signal \SYNTHESIZED_WIRE_10_0\ : std_logic;
signal \SYNTHESIZED_WIRE_5_0\ : std_logic;
signal \SYNTHESIZED_WIRE_5_4\ : std_logic;
signal \b2v_inst.un12_pix_count_intlto7_N_2LZ0Z1_cascade_\ : std_logic;
signal \b2v_inst.un13_pix_count_int_li_0\ : std_logic;
signal \b2v_inst.un13_pix_count_int_li_0_cascade_\ : std_logic;
signal \SYNTHESIZED_WIRE_10_1\ : std_logic;
signal \SYNTHESIZED_WIRE_5_1\ : std_logic;
signal \SYNTHESIZED_WIRE_10_2\ : std_logic;
signal \SYNTHESIZED_WIRE_5_2\ : std_logic;
signal \b2v_inst.state_fastZ0Z_19\ : std_logic;
signal \b2v_inst9.fsm_state_srsts_1_0\ : std_logic;
signal \b2v_inst9.N_522\ : std_logic;
signal \b2v_inst9.N_522_cascade_\ : std_logic;
signal \b2v_inst9.fsm_stateZ0Z_0\ : std_logic;
signal \b2v_inst9.fsm_stateZ0Z_1\ : std_logic;
signal \b2v_inst9.N_84_2_cascade_\ : std_logic;
signal \b2v_inst9.N_582\ : std_logic;
signal \bfn_17_5_0_\ : std_logic;
signal \b2v_inst.valor_max_final4_2_cry_0\ : std_logic;
signal \b2v_inst.valor_max_final4_2_cry_1\ : std_logic;
signal \b2v_inst.valor_max_final4_2_cry_2\ : std_logic;
signal \b2v_inst.valor_max_final4_2_cry_3\ : std_logic;
signal \b2v_inst.valor_max_final4_2_cry_4\ : std_logic;
signal \b2v_inst.valor_max_final4_2_cry_5\ : std_logic;
signal \b2v_inst.valor_max_final4_2_cry_6\ : std_logic;
signal \b2v_inst.valor_max_final4_2_cry_7\ : std_logic;
signal \bfn_17_6_0_\ : std_logic;
signal \b2v_inst.valor_max_final4_2_cry_8\ : std_logic;
signal \b2v_inst.valor_max_final4_2_cry_9\ : std_logic;
signal \b2v_inst.valor_max_final42\ : std_logic;
signal \b2v_inst.data_a_escribir11_7_and\ : std_logic;
signal \SYNTHESIZED_WIRE_3_7\ : std_logic;
signal \SYNTHESIZED_WIRE_3_8\ : std_logic;
signal \SYNTHESIZED_WIRE_3_0\ : std_logic;
signal \b2v_inst.reg_ancho_2Z0Z_0\ : std_logic;
signal \bfn_17_8_0_\ : std_logic;
signal \b2v_inst.valor_max_final4_3_cry_0\ : std_logic;
signal \b2v_inst.valor_max_final4_3_cry_1\ : std_logic;
signal \b2v_inst.valor_max_final4_3_cry_2\ : std_logic;
signal \b2v_inst.valor_max_final4_3_cry_3\ : std_logic;
signal \b2v_inst.reg_ancho_2Z0Z_5\ : std_logic;
signal \b2v_inst.valor_max_final4_3_cry_4\ : std_logic;
signal \b2v_inst.reg_ancho_2Z0Z_6\ : std_logic;
signal \b2v_inst.valor_max_final4_3_cry_5\ : std_logic;
signal \b2v_inst.reg_ancho_2Z0Z_7\ : std_logic;
signal \b2v_inst.valor_max_final4_3_cry_6\ : std_logic;
signal \b2v_inst.valor_max_final4_3_cry_7\ : std_logic;
signal \bfn_17_9_0_\ : std_logic;
signal \b2v_inst.valor_max_final4_3_cry_8\ : std_logic;
signal \b2v_inst.valor_max_final4_3_cry_9\ : std_logic;
signal \b2v_inst.valor_max_final43\ : std_logic;
signal \b2v_inst.data_a_escribir_RNO_0Z0Z_0\ : std_logic;
signal \b2v_inst.data_a_escribir_RNO_0Z0Z_1\ : std_logic;
signal \b2v_inst.eventosZ0Z_5\ : std_logic;
signal \b2v_inst.reg_anterior_i_0\ : std_logic;
signal \bfn_17_10_0_\ : std_logic;
signal \b2v_inst.reg_anterior_i_1\ : std_logic;
signal \b2v_inst.valor_max_final4_1_cry_0\ : std_logic;
signal \b2v_inst.reg_anterior_i_2\ : std_logic;
signal \b2v_inst.valor_max_final4_1_cry_1\ : std_logic;
signal \b2v_inst.reg_anterior_i_3\ : std_logic;
signal \b2v_inst.valor_max_final4_1_cry_2\ : std_logic;
signal \b2v_inst.reg_anterior_i_4\ : std_logic;
signal \b2v_inst.valor_max_final4_1_cry_3\ : std_logic;
signal \b2v_inst.reg_anterior_i_5\ : std_logic;
signal \b2v_inst.valor_max_final4_1_cry_4\ : std_logic;
signal \b2v_inst.reg_anterior_i_6\ : std_logic;
signal \b2v_inst.valor_max_final4_1_cry_5\ : std_logic;
signal \b2v_inst.reg_anterior_i_7\ : std_logic;
signal \b2v_inst.valor_max_final4_1_cry_6\ : std_logic;
signal \b2v_inst.valor_max_final4_1_cry_7\ : std_logic;
signal \b2v_inst.reg_anterior_i_8\ : std_logic;
signal \bfn_17_11_0_\ : std_logic;
signal \b2v_inst.reg_anterior_i_9\ : std_logic;
signal \b2v_inst.valor_max_final4_1_cry_8\ : std_logic;
signal \b2v_inst.reg_anterior_i_10\ : std_logic;
signal \b2v_inst.valor_max_final4_1_cry_9\ : std_logic;
signal \b2v_inst.valor_max_final43_THRU_CO\ : std_logic;
signal \b2v_inst.m54_ns_1\ : std_logic;
signal \b2v_inst.valor_max_final41\ : std_logic;
signal \b2v_inst.stateZ0Z_6\ : std_logic;
signal \b2v_inst.stateZ0Z_10\ : std_logic;
signal \b2v_inst.stateZ0Z_29\ : std_logic;
signal \b2v_inst.state_ns_a3_i_0_a2_1_4_1\ : std_logic;
signal b2v_inst_state_3 : std_logic;
signal \b2v_inst.N_694\ : std_logic;
signal \b2v_inst.N_695_cascade_\ : std_logic;
signal \b2v_inst.state_ns_a3_i_0_1_1\ : std_logic;
signal \b2v_inst.un2_cuentalto10_i_a2_8\ : std_logic;
signal \b2v_inst.un2_cuentalto10_i_a2_7\ : std_logic;
signal \b2v_inst.state_32_repZ0Z1\ : std_logic;
signal reset_c : std_logic;
signal \b2v_inst.N_654_2\ : std_logic;
signal \b2v_inst.un1_reset_inv_0_0_tz_cascade_\ : std_logic;
signal \b2v_inst.N_482\ : std_logic;
signal \b2v_inst.eventosZ0Z_7\ : std_logic;
signal \b2v_inst.data_a_escribir_RNO_2Z0Z_7\ : std_logic;
signal \bfn_17_13_0_\ : std_logic;
signal \b2v_inst9.un1_cycle_counter_2_cry_0\ : std_logic;
signal \b2v_inst9.un1_cycle_counter_2_cry_1\ : std_logic;
signal \b2v_inst9.un1_cycle_counter_2_cry_2\ : std_logic;
signal \b2v_inst9.cycle_counterZ0Z_3\ : std_logic;
signal \b2v_inst9.cycle_counter_RNIQAGDZ0Z_3_cascade_\ : std_logic;
signal \b2v_inst9.un1_cycle_counter_2_cry_0_THRU_CO\ : std_logic;
signal \b2v_inst9.cycle_counterZ0Z_1\ : std_logic;
signal \SYNTHESIZED_WIRE_5_7\ : std_logic;
signal \SYNTHESIZED_WIRE_5_6\ : std_logic;
signal \b2v_inst.un12_pix_count_intlto7_N_3LZ0Z3\ : std_logic;
signal \SYNTHESIZED_WIRE_10_5\ : std_logic;
signal \SYNTHESIZED_WIRE_5_5\ : std_logic;
signal \b2v_inst4.pix_count_int_0_sqmuxa\ : std_logic;
signal \b2v_inst9.N_175_i\ : std_logic;
signal \b2v_inst9.bit_counterZ0Z_0\ : std_logic;
signal \bfn_17_16_0_\ : std_logic;
signal \b2v_inst9.bit_counterZ1Z_1\ : std_logic;
signal \b2v_inst9.un1_bit_counter_3_cry_0\ : std_logic;
signal \b2v_inst9.bit_counterZ0Z_2\ : std_logic;
signal \b2v_inst9.un1_bit_counter_3_cry_1\ : std_logic;
signal \b2v_inst9.fsm_state_RNIND1P1Z0Z_0\ : std_logic;
signal \b2v_inst9.un1_bit_counter_3_cry_2\ : std_logic;
signal \b2v_inst9.bit_counterZ0Z_3\ : std_logic;
signal \b2v_inst.reg_anteriorZ0Z_0\ : std_logic;
signal \bfn_18_6_0_\ : std_logic;
signal \b2v_inst.reg_anteriorZ0Z_1\ : std_logic;
signal \b2v_inst.un2_valor_max2_cry_0\ : std_logic;
signal \b2v_inst.un2_valor_max2_cry_1\ : std_logic;
signal \b2v_inst.un2_valor_max2_cry_2\ : std_logic;
signal \b2v_inst.un2_valor_max2_cry_3\ : std_logic;
signal \b2v_inst.un2_valor_max2_cry_4\ : std_logic;
signal \b2v_inst.un2_valor_max2_cry_5\ : std_logic;
signal \b2v_inst.un2_valor_max2_cry_6\ : std_logic;
signal \b2v_inst.un2_valor_max2_cry_7\ : std_logic;
signal \bfn_18_7_0_\ : std_logic;
signal \b2v_inst.un2_valor_max2_cry_8\ : std_logic;
signal \b2v_inst.un2_valor_max2_cry_9\ : std_logic;
signal \b2v_inst.un2_valor_max2\ : std_logic;
signal \b2v_inst.reg_anteriorZ0Z_3\ : std_logic;
signal \b2v_inst.data_a_escribir_RNO_0Z0Z_3\ : std_logic;
signal \b2v_inst.reg_anteriorZ0Z_5\ : std_logic;
signal \b2v_inst.reg_ancho_1Z0Z_0\ : std_logic;
signal \b2v_inst.reg_ancho_3_i_0\ : std_logic;
signal \bfn_18_8_0_\ : std_logic;
signal \b2v_inst.reg_ancho_1Z0Z_1\ : std_logic;
signal \b2v_inst.reg_ancho_3_i_1\ : std_logic;
signal \b2v_inst.valor_max_final4_0_cry_0\ : std_logic;
signal \b2v_inst.reg_ancho_3_i_2\ : std_logic;
signal \b2v_inst.valor_max_final4_0_cry_1\ : std_logic;
signal \b2v_inst.reg_ancho_3_i_3\ : std_logic;
signal \b2v_inst.valor_max_final4_0_cry_2\ : std_logic;
signal \b2v_inst.reg_ancho_1Z0Z_4\ : std_logic;
signal \b2v_inst.reg_ancho_3_i_4\ : std_logic;
signal \b2v_inst.valor_max_final4_0_cry_3\ : std_logic;
signal \b2v_inst.reg_ancho_1Z0Z_5\ : std_logic;
signal \b2v_inst.reg_ancho_3_i_5\ : std_logic;
signal \b2v_inst.valor_max_final4_0_cry_4\ : std_logic;
signal \b2v_inst.reg_ancho_1Z0Z_6\ : std_logic;
signal \b2v_inst.reg_ancho_3Z0Z_6\ : std_logic;
signal \b2v_inst.reg_ancho_3_i_6\ : std_logic;
signal \b2v_inst.valor_max_final4_0_cry_5\ : std_logic;
signal \b2v_inst.reg_ancho_1Z0Z_7\ : std_logic;
signal \b2v_inst.reg_ancho_3_i_7\ : std_logic;
signal \b2v_inst.valor_max_final4_0_cry_6\ : std_logic;
signal \b2v_inst.valor_max_final4_0_cry_7\ : std_logic;
signal \b2v_inst.reg_ancho_3_i_8\ : std_logic;
signal \bfn_18_9_0_\ : std_logic;
signal \b2v_inst.reg_ancho_3_i_9\ : std_logic;
signal \b2v_inst.valor_max_final4_0_cry_8\ : std_logic;
signal \b2v_inst.reg_ancho_1Z0Z_10\ : std_logic;
signal \b2v_inst.reg_ancho_3_i_10\ : std_logic;
signal \b2v_inst.valor_max_final4_0_cry_9\ : std_logic;
signal \b2v_inst.valor_max_final40\ : std_logic;
signal \b2v_inst.valor_max_final40_THRU_CO\ : std_logic;
signal \b2v_inst.reg_ancho_1Z0Z_9\ : std_logic;
signal \b2v_inst.reg_ancho_1Z0Z_8\ : std_logic;
signal \b2v_inst.reg_ancho_2Z0Z_8\ : std_logic;
signal \b2v_inst.eventosZ0Z_3\ : std_logic;
signal \b2v_inst.un1_reg_anterior_0_i_1_3\ : std_logic;
signal \b2v_inst.reg_anteriorZ0Z_2\ : std_logic;
signal \b2v_inst.data_a_escribir11_6_and\ : std_logic;
signal \b2v_inst.N_273\ : std_logic;
signal \b2v_inst.un1_reg_anterior_iv_0_0_5\ : std_logic;
signal \b2v_inst.N_267\ : std_logic;
signal \b2v_inst.un1_reg_anterior_iv_0_1_5_cascade_\ : std_logic;
signal \b2v_inst.data_a_escribir_RNO_0Z0Z_2\ : std_logic;
signal \b2v_inst.reg_ancho_2Z0Z_9\ : std_logic;
signal \b2v_inst.reg_ancho_3Z0Z_1\ : std_logic;
signal \b2v_inst.reg_ancho_3Z0Z_0\ : std_logic;
signal \b2v_inst.data_a_escribir11_5_and\ : std_logic;
signal \b2v_inst.reg_ancho_3Z0Z_9\ : std_logic;
signal \b2v_inst.eventosZ0Z_9\ : std_logic;
signal \b2v_inst.N_545\ : std_logic;
signal \b2v_inst.un1_reg_anterior_iv_0_0_0_9_cascade_\ : std_logic;
signal \b2v_inst.N_543\ : std_logic;
signal \b2v_inst.un1_reg_anterior_iv_0_0_1_9_cascade_\ : std_logic;
signal \b2v_inst.valor_max2_6\ : std_logic;
signal \b2v_inst.un1_reg_anterior_iv_0_1_6\ : std_logic;
signal \b2v_inst.data_a_escribir11_10_and\ : std_logic;
signal \b2v_inst.eventosZ0Z_8\ : std_logic;
signal \b2v_inst.un1_reg_anterior_iv_0_0_0_8_cascade_\ : std_logic;
signal \b2v_inst.N_542\ : std_logic;
signal \b2v_inst.un1_reg_anterior_iv_0_0_1_8_cascade_\ : std_logic;
signal \b2v_inst.reg_anteriorZ0Z_8\ : std_logic;
signal \b2v_inst.reg_ancho_3Z0Z_8\ : std_logic;
signal \b2v_inst.N_544\ : std_logic;
signal \b2v_inst.reg_ancho_3Z0Z_7\ : std_logic;
signal \b2v_inst.reg_anteriorZ0Z_7\ : std_logic;
signal \b2v_inst.un1_reg_anterior_0_i_1_7\ : std_logic;
signal \b2v_inst.data_a_escribir_RNO_0Z0Z_7_cascade_\ : std_logic;
signal \b2v_inst.N_711\ : std_logic;
signal \b2v_inst.un1_reset_inv_0\ : std_logic;
signal \b2v_inst9.un1_cycle_counter_2_cry_1_THRU_CO\ : std_logic;
signal \b2v_inst9.cycle_counterZ0Z_2\ : std_logic;
signal \b2v_inst9.cycle_counter_RNIQAGDZ0Z_3\ : std_logic;
signal \N_478\ : std_logic;
signal \b2v_inst9.cycle_counterZ0Z_0\ : std_logic;
signal \SYNTHESIZED_WIRE_5_3\ : std_logic;
signal \b2v_inst.pix_data_regZ0Z_3\ : std_logic;
signal \b2v_inst.stateZ0Z_24\ : std_logic;
signal \SYNTHESIZED_WIRE_1_2\ : std_logic;
signal \b2v_inst.reg_anteriorZ0Z_4\ : std_logic;
signal \SYNTHESIZED_WIRE_3_6\ : std_logic;
signal \b2v_inst.reg_anteriorZ0Z_6\ : std_logic;
signal \b2v_inst.reg_ancho_2Z0Z_10\ : std_logic;
signal \b2v_inst.reg_ancho_3Z0Z_4\ : std_logic;
signal \b2v_inst.data_a_escribir11_3_and\ : std_logic;
signal \SYNTHESIZED_WIRE_3_1\ : std_logic;
signal \b2v_inst.reg_ancho_2Z0Z_1\ : std_logic;
signal \b2v_inst.reg_ancho_2Z0Z_2\ : std_logic;
signal \b2v_inst.reg_ancho_1Z0Z_2\ : std_logic;
signal \b2v_inst.eventosZ0Z_2\ : std_logic;
signal \b2v_inst.data_a_escribir_RNO_2Z0Z_2_cascade_\ : std_logic;
signal \b2v_inst.data_a_escribir12_THRU_CO\ : std_logic;
signal \b2v_inst.un1_reg_anterior_0_i_1_2\ : std_logic;
signal \b2v_inst.reg_ancho_1Z0Z_3\ : std_logic;
signal \b2v_inst.stateZ0Z_20\ : std_logic;
signal \b2v_inst.un2_valor_max1_THRU_CO\ : std_logic;
signal \b2v_inst.data_a_escribir_RNO_2Z0Z_3\ : std_logic;
signal \b2v_inst.reg_ancho_2Z0Z_3\ : std_logic;
signal \b2v_inst.un2_valor_max2_THRU_CO\ : std_logic;
signal \b2v_inst.N_264\ : std_logic;
signal \b2v_inst.reg_ancho_3Z0Z_10\ : std_logic;
signal \SYNTHESIZED_WIRE_3_3\ : std_logic;
signal \b2v_inst.reg_ancho_3Z0Z_3\ : std_logic;
signal \SYNTHESIZED_WIRE_3_2\ : std_logic;
signal \b2v_inst.reg_ancho_3Z0Z_2\ : std_logic;
signal \SYNTHESIZED_WIRE_3_5\ : std_logic;
signal \b2v_inst.reg_ancho_3Z0Z_5\ : std_logic;
signal \b2v_inst.stateZ0Z_21\ : std_logic;
signal \SYNTHESIZED_WIRE_3_9\ : std_logic;
signal \b2v_inst.reg_anteriorZ0Z_9\ : std_logic;
signal \b2v_inst.ignorar_anteriorZ0\ : std_logic;
signal \SYNTHESIZED_WIRE_3_10\ : std_logic;
signal \b2v_inst.reg_anteriorZ0Z_10\ : std_logic;
signal \b2v_inst.stateZ0Z_27\ : std_logic;
signal \SYNTHESIZED_WIRE_1_0\ : std_logic;
signal \SYNTHESIZED_WIRE_1_1\ : std_logic;
signal \SYNTHESIZED_WIRE_1_4\ : std_logic;
signal \bfn_19_14_0_\ : std_logic;
signal b2v_inst_cantidad_temp_2 : std_logic;
signal \b2v_inst.un16_data_ram_cantidad_o_cry_1\ : std_logic;
signal \b2v_inst.un16_data_ram_cantidad_o_cry_2\ : std_logic;
signal b2v_inst_cantidad_temp_4 : std_logic;
signal \b2v_inst.un16_data_ram_cantidad_o_cry_3\ : std_logic;
signal b2v_inst_cantidad_temp_5 : std_logic;
signal \b2v_inst.un16_data_ram_cantidad_o_cry_4\ : std_logic;
signal \b2v_inst.un16_data_ram_cantidad_o_cry_1_c_RNI77COZ0\ : std_logic;
signal \N_553_i\ : std_logic;
signal \b2v_inst.un16_data_ram_cantidad_o_cry_3_c_RNIBDEOZ0\ : std_logic;
signal b2v_inst_data_a_escribir_4 : std_logic;
signal \N_549_i\ : std_logic;
signal \b2v_inst.un16_data_ram_cantidad_o_cry_2_c_RNI9ADOZ0\ : std_logic;
signal b2v_inst_data_a_escribir_3 : std_logic;
signal \N_551_i\ : std_logic;
signal \b2v_inst.N_481\ : std_logic;
signal \N_121_i\ : std_logic;
signal b2v_inst_data_a_escribir_2 : std_logic;
signal \N_118_i\ : std_logic;
signal \SYNTHESIZED_WIRE_3_4\ : std_logic;
signal \b2v_inst.reg_ancho_2Z0Z_4\ : std_logic;
signal \b2v_inst.stateZ0Z_23\ : std_logic;
signal b2v_inst_data_a_escribir_9 : std_logic;
signal \N_111_i\ : std_logic;
signal \b2v_inst.addr_ram_iv_i_1_6\ : std_logic;
signal \b2v_inst.addr_ram_iv_i_0_6\ : std_logic;
signal \N_298\ : std_logic;
signal \b2v_inst.addr_ram_iv_i_0_5\ : std_logic;
signal \b2v_inst.addr_ram_iv_i_1_5\ : std_logic;
signal \indice_RNIS8333_5\ : std_logic;
signal \b2v_inst.addr_ram_iv_i_0_8\ : std_logic;
signal \b2v_inst.addr_ram_iv_i_1_8\ : std_logic;
signal \indice_RNIBO333_8\ : std_logic;
signal \b2v_inst.addr_ram_iv_i_0_9\ : std_logic;
signal \b2v_inst.addr_ram_iv_i_1_9\ : std_logic;
signal \indice_RNIGT333_9\ : std_logic;
signal \N_115_i\ : std_logic;
signal b2v_inst_data_a_escribir_10 : std_logic;
signal \N_110_i\ : std_logic;
signal \b2v_inst.addr_ram_iv_i_0_0\ : std_logic;
signal \b2v_inst.addr_ram_iv_i_1_0\ : std_logic;
signal \indice_RNI3F233_0\ : std_logic;
signal \b2v_inst.addr_ram_iv_i_0_10\ : std_logic;
signal \b2v_inst.addr_ram_iv_i_1_10\ : std_logic;
signal \N_37\ : std_logic;
signal b2v_inst_data_a_escribir_8 : std_logic;
signal \N_112_i\ : std_logic;
signal b2v_inst_data_a_escribir_7 : std_logic;
signal \N_113_i\ : std_logic;
signal \b2v_inst.addr_ram_iv_i_0_0_1\ : std_logic;
signal \b2v_inst.addr_ram_iv_i_0_1_1\ : std_logic;
signal \indice_RNI8K233_1\ : std_logic;
signal b2v_inst_data_a_escribir_6 : std_logic;
signal \N_114_i\ : std_logic;
signal \b2v_inst.addr_ram_iv_i_0_2\ : std_logic;
signal \b2v_inst.N_480\ : std_logic;
signal \b2v_inst.addr_ram_iv_i_1_2\ : std_logic;
signal \indice_RNIDP233_2\ : std_logic;
signal b2v_inst_data_a_escribir_0 : std_logic;
signal \N_557_i\ : std_logic;
signal b2v_inst_cantidad_temp_0 : std_logic;
signal b2v_inst_cantidad_temp_1 : std_logic;
signal b2v_inst_data_a_escribir_1 : std_logic;
signal \b2v_inst.cantidad_temp_RNILL3KZ0Z_1_cascade_\ : std_logic;
signal \N_555_i\ : std_logic;
signal \b2v_inst.stateZ0Z_18\ : std_logic;
signal \SYNTHESIZED_WIRE_1_3\ : std_logic;
signal \b2v_inst.stateZ0Z_9\ : std_logic;
signal b2v_inst_cantidad_temp_3 : std_logic;
signal clk_c_g : std_logic;
signal reset_c_i_g : std_logic;
signal \b2v_inst.N_828\ : std_logic;
signal \b2v_inst.un16_data_ram_cantidad_o_cry_4_c_RNIDGFOZ0\ : std_logic;
signal b2v_inst_data_a_escribir_5 : std_logic;
signal \b2v_inst.N_514\ : std_logic;
signal \N_547_i\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \b2v_inst.dir_energiaZ0Z_10\ : std_logic;
signal \b2v_inst.indiceZ0Z_10\ : std_logic;
signal \N_445_i\ : std_logic;
signal \b2v_inst.indiceZ0Z_3\ : std_logic;
signal \b2v_inst.dir_energiaZ0Z_3\ : std_logic;
signal \N_357_i\ : std_logic;
signal \b2v_inst.indiceZ0Z_4\ : std_logic;
signal \b2v_inst.dir_energiaZ0Z_4\ : std_logic;
signal \N_356_i\ : std_logic;
signal \b2v_inst.dir_energiaZ0Z_2\ : std_logic;
signal \b2v_inst.indiceZ0Z_2\ : std_logic;
signal \N_358_i\ : std_logic;
signal \b2v_inst.indiceZ0Z_9\ : std_logic;
signal \b2v_inst.dir_energiaZ0Z_9\ : std_logic;
signal \N_444_i\ : std_logic;
signal \b2v_inst.indiceZ0Z_5\ : std_logic;
signal \b2v_inst.dir_energiaZ0Z_5\ : std_logic;
signal \N_355_i\ : std_logic;
signal \b2v_inst.dir_energiaZ0Z_0\ : std_logic;
signal \b2v_inst.indiceZ0Z_0\ : std_logic;
signal \N_360_i\ : std_logic;
signal \b2v_inst.dir_energiaZ0Z_8\ : std_logic;
signal \b2v_inst.indiceZ0Z_8\ : std_logic;
signal \N_443_i\ : std_logic;
signal \b2v_inst.dir_energiaZ0Z_7\ : std_logic;
signal \b2v_inst.indiceZ0Z_7\ : std_logic;
signal \N_353_i\ : std_logic;
signal \b2v_inst.dir_energiaZ0Z_1\ : std_logic;
signal \b2v_inst.indiceZ0Z_1\ : std_logic;
signal \N_359_i\ : std_logic;
signal \b2v_inst.N_645\ : std_logic;
signal \b2v_inst.dir_energiaZ0Z_6\ : std_logic;
signal \b2v_inst.indiceZ0Z_6\ : std_logic;
signal \b2v_inst.N_484\ : std_logic;
signal \N_354_i\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal clk_wire : std_logic;
signal leds_wire : std_logic_vector(13 downto 0);
signal swit_wire : std_logic_vector(10 downto 0);
signal uart_rx_i_wire : std_logic;
signal reset_wire : std_logic;
signal uart_tx_o_wire : std_logic;
signal \b2v_inst2.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \b2v_inst2.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \b2v_inst2.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \b2v_inst2.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \b2v_inst2.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \b2v_inst8.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \b2v_inst8.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \b2v_inst8.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \b2v_inst8.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \b2v_inst8.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \b2v_inst7.mem_mem_0_2_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \b2v_inst7.mem_mem_0_2_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \b2v_inst7.mem_mem_0_2_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \b2v_inst7.mem_mem_0_2_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \b2v_inst7.mem_mem_0_2_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \b2v_inst2.mem_mem_0_2_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \b2v_inst2.mem_mem_0_2_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \b2v_inst2.mem_mem_0_2_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \b2v_inst2.mem_mem_0_2_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \b2v_inst2.mem_mem_0_2_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \b2v_inst2.mem_mem_0_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \b2v_inst2.mem_mem_0_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \b2v_inst2.mem_mem_0_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \b2v_inst2.mem_mem_0_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \b2v_inst2.mem_mem_0_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \b2v_inst8.mem_mem_0_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \b2v_inst8.mem_mem_0_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \b2v_inst8.mem_mem_0_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \b2v_inst8.mem_mem_0_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \b2v_inst8.mem_mem_0_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \b2v_inst7.mem_mem_0_4_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \b2v_inst7.mem_mem_0_4_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \b2v_inst7.mem_mem_0_4_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \b2v_inst7.mem_mem_0_4_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \b2v_inst7.mem_mem_0_4_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \b2v_inst7.mem_mem_0_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \b2v_inst7.mem_mem_0_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \b2v_inst7.mem_mem_0_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \b2v_inst7.mem_mem_0_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \b2v_inst7.mem_mem_0_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \b2v_inst2.mem_mem_0_4_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \b2v_inst2.mem_mem_0_4_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \b2v_inst2.mem_mem_0_4_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \b2v_inst2.mem_mem_0_4_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \b2v_inst2.mem_mem_0_4_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \b2v_inst2.mem_mem_0_3_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \b2v_inst2.mem_mem_0_3_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \b2v_inst2.mem_mem_0_3_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \b2v_inst2.mem_mem_0_3_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \b2v_inst2.mem_mem_0_3_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \b2v_inst7.mem_mem_0_6_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \b2v_inst7.mem_mem_0_6_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \b2v_inst7.mem_mem_0_6_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \b2v_inst7.mem_mem_0_6_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \b2v_inst7.mem_mem_0_6_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \b2v_inst8.mem_mem_0_2_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \b2v_inst8.mem_mem_0_2_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \b2v_inst8.mem_mem_0_2_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \b2v_inst8.mem_mem_0_2_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \b2v_inst8.mem_mem_0_2_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \b2v_inst7.mem_mem_0_3_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \b2v_inst7.mem_mem_0_3_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \b2v_inst7.mem_mem_0_3_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \b2v_inst7.mem_mem_0_3_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \b2v_inst7.mem_mem_0_3_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \b2v_inst7.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \b2v_inst7.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \b2v_inst7.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \b2v_inst7.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \b2v_inst7.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \b2v_inst2.mem_mem_0_5_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \b2v_inst2.mem_mem_0_5_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \b2v_inst2.mem_mem_0_5_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \b2v_inst2.mem_mem_0_5_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \b2v_inst2.mem_mem_0_5_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \b2v_inst7.mem_mem_0_5_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \b2v_inst7.mem_mem_0_5_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \b2v_inst7.mem_mem_0_5_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \b2v_inst7.mem_mem_0_5_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \b2v_inst7.mem_mem_0_5_physical_WDATA_wire\ : std_logic_vector(15 downto 0);

begin
    clk_wire <= clk;
    leds <= leds_wire;
    swit_wire <= swit;
    uart_rx_i_wire <= uart_rx_i;
    reset_wire <= reset;
    uart_tx_o <= uart_tx_o_wire;
    \SYNTHESIZED_WIRE_3_1\ <= \b2v_inst2.mem_mem_0_0_physical_RDATA_wire\(11);
    \SYNTHESIZED_WIRE_3_0\ <= \b2v_inst2.mem_mem_0_0_physical_RDATA_wire\(3);
    \b2v_inst2.mem_mem_0_0_physical_RADDR_wire\ <= \N__33476\&\N__33778\&\N__33892\&\N__19472\&\N__32785\&\N__34009\&\N__18469\&\N__19651\&\N__35057\&\N__35410\&\N__33590\;
    \b2v_inst2.mem_mem_0_0_physical_WADDR_wire\ <= \N__33475\&\N__33779\&\N__33893\&\N__19471\&\N__32786\&\N__34010\&\N__18473\&\N__19658\&\N__35056\&\N__35411\&\N__33589\;
    \b2v_inst2.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \b2v_inst2.mem_mem_0_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__20372\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__33146\&'0'&'0'&'0';
    \SYNTHESIZED_WIRE_1_1\ <= \b2v_inst8.mem_mem_0_0_physical_RDATA_wire\(11);
    \SYNTHESIZED_WIRE_1_0\ <= \b2v_inst8.mem_mem_0_0_physical_RDATA_wire\(3);
    \b2v_inst8.mem_mem_0_0_physical_RADDR_wire\ <= \N__36625\&\N__35770\&\N__38969\&\N__38756\&\N__38198\&\N__35548\&\N__36208\&\N__36421\&\N__35998\&\N__38510\&\N__39188\;
    \b2v_inst8.mem_mem_0_0_physical_WADDR_wire\ <= \N__36629\&\N__35771\&\N__38968\&\N__38755\&\N__38197\&\N__35549\&\N__36209\&\N__36422\&\N__35999\&\N__38509\&\N__39187\;
    \b2v_inst8.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \b2v_inst8.mem_mem_0_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__34772\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__34916\&'0'&'0'&'0';
    leds_c_5 <= \b2v_inst7.mem_mem_0_2_physical_RDATA_wire\(11);
    leds_c_4 <= \b2v_inst7.mem_mem_0_2_physical_RDATA_wire\(3);
    \b2v_inst7.mem_mem_0_2_physical_RADDR_wire\ <= \N__20128\&\N__15955\&\N__14149\&\N__14332\&\N__18703\&\N__19879\&\N__21574\&\N__20512\&\N__19996\&\N__14428\&\N__14239\;
    \b2v_inst7.mem_mem_0_2_physical_WADDR_wire\ <= \N__20125\&\N__15952\&\N__14146\&\N__14341\&\N__18700\&\N__19876\&\N__21571\&\N__20509\&\N__19993\&\N__14431\&\N__14242\;
    \b2v_inst7.mem_mem_0_2_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \b2v_inst7.mem_mem_0_2_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__23621\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19715\&'0'&'0'&'0';
    \SYNTHESIZED_WIRE_3_5\ <= \b2v_inst2.mem_mem_0_2_physical_RDATA_wire\(11);
    \SYNTHESIZED_WIRE_3_4\ <= \b2v_inst2.mem_mem_0_2_physical_RDATA_wire\(3);
    \b2v_inst2.mem_mem_0_2_physical_RADDR_wire\ <= \N__33454\&\N__33754\&\N__33868\&\N__19450\&\N__32761\&\N__33985\&\N__18445\&\N__19627\&\N__35035\&\N__35386\&\N__33568\;
    \b2v_inst2.mem_mem_0_2_physical_WADDR_wire\ <= \N__33451\&\N__33757\&\N__33871\&\N__19447\&\N__32764\&\N__33988\&\N__18454\&\N__19642\&\N__35032\&\N__35389\&\N__33565\;
    \b2v_inst2.mem_mem_0_2_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \b2v_inst2.mem_mem_0_2_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__33698\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19754\&'0'&'0'&'0';
    \SYNTHESIZED_WIRE_3_3\ <= \b2v_inst2.mem_mem_0_1_physical_RDATA_wire\(11);
    \SYNTHESIZED_WIRE_3_2\ <= \b2v_inst2.mem_mem_0_1_physical_RDATA_wire\(3);
    \b2v_inst2.mem_mem_0_1_physical_RADDR_wire\ <= \N__33466\&\N__33766\&\N__33880\&\N__19462\&\N__32773\&\N__33997\&\N__18457\&\N__19639\&\N__35047\&\N__35398\&\N__33580\;
    \b2v_inst2.mem_mem_0_1_physical_WADDR_wire\ <= \N__33463\&\N__33769\&\N__33883\&\N__19459\&\N__32776\&\N__34000\&\N__18466\&\N__19652\&\N__35044\&\N__35401\&\N__33577\;
    \b2v_inst2.mem_mem_0_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \b2v_inst2.mem_mem_0_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__20555\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__33071\&'0'&'0'&'0';
    \SYNTHESIZED_WIRE_1_3\ <= \b2v_inst8.mem_mem_0_1_physical_RDATA_wire\(11);
    \SYNTHESIZED_WIRE_1_2\ <= \b2v_inst8.mem_mem_0_1_physical_RDATA_wire\(3);
    \b2v_inst8.mem_mem_0_1_physical_RADDR_wire\ <= \N__36613\&\N__35758\&\N__38959\&\N__38746\&\N__38188\&\N__35536\&\N__36196\&\N__36409\&\N__35986\&\N__38500\&\N__39178\;
    \b2v_inst8.mem_mem_0_1_physical_WADDR_wire\ <= \N__36622\&\N__35761\&\N__38956\&\N__38743\&\N__38185\&\N__35539\&\N__36199\&\N__36412\&\N__35989\&\N__38497\&\N__39175\;
    \b2v_inst8.mem_mem_0_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \b2v_inst8.mem_mem_0_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__33197\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__32558\&'0'&'0'&'0';
    leds_c_9 <= \b2v_inst7.mem_mem_0_4_physical_RDATA_wire\(11);
    leds_c_8 <= \b2v_inst7.mem_mem_0_4_physical_RDATA_wire\(3);
    \b2v_inst7.mem_mem_0_4_physical_RADDR_wire\ <= \N__20104\&\N__15931\&\N__14125\&\N__14308\&\N__18679\&\N__19855\&\N__21550\&\N__20488\&\N__19972\&\N__14404\&\N__14215\;
    \b2v_inst7.mem_mem_0_4_physical_WADDR_wire\ <= \N__20101\&\N__15928\&\N__14122\&\N__14317\&\N__18676\&\N__19852\&\N__21547\&\N__20485\&\N__19969\&\N__14407\&\N__14218\;
    \b2v_inst7.mem_mem_0_4_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \b2v_inst7.mem_mem_0_4_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__16949\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__16940\&'0'&'0'&'0';
    leds_c_3 <= \b2v_inst7.mem_mem_0_1_physical_RDATA_wire\(11);
    leds_c_2 <= \b2v_inst7.mem_mem_0_1_physical_RDATA_wire\(3);
    \b2v_inst7.mem_mem_0_1_physical_RADDR_wire\ <= \N__20140\&\N__15967\&\N__14161\&\N__14344\&\N__18715\&\N__19891\&\N__21586\&\N__20524\&\N__20008\&\N__14440\&\N__14251\;
    \b2v_inst7.mem_mem_0_1_physical_WADDR_wire\ <= \N__20137\&\N__15964\&\N__14158\&\N__14353\&\N__18712\&\N__19888\&\N__21583\&\N__20521\&\N__20005\&\N__14443\&\N__14254\;
    \b2v_inst7.mem_mem_0_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \b2v_inst7.mem_mem_0_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__21917\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__21206\&'0'&'0'&'0';
    \SYNTHESIZED_WIRE_3_9\ <= \b2v_inst2.mem_mem_0_4_physical_RDATA_wire\(11);
    \SYNTHESIZED_WIRE_3_8\ <= \b2v_inst2.mem_mem_0_4_physical_RDATA_wire\(3);
    \b2v_inst2.mem_mem_0_4_physical_RADDR_wire\ <= \N__33430\&\N__33730\&\N__33844\&\N__19426\&\N__32737\&\N__33961\&\N__18421\&\N__19603\&\N__35011\&\N__35362\&\N__33544\;
    \b2v_inst2.mem_mem_0_4_physical_WADDR_wire\ <= \N__33427\&\N__33733\&\N__33847\&\N__19423\&\N__32740\&\N__33964\&\N__18430\&\N__19618\&\N__35008\&\N__35365\&\N__33541\;
    \b2v_inst2.mem_mem_0_4_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \b2v_inst2.mem_mem_0_4_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__32825\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__33356\&'0'&'0'&'0';
    \SYNTHESIZED_WIRE_3_7\ <= \b2v_inst2.mem_mem_0_3_physical_RDATA_wire\(11);
    \SYNTHESIZED_WIRE_3_6\ <= \b2v_inst2.mem_mem_0_3_physical_RDATA_wire\(3);
    \b2v_inst2.mem_mem_0_3_physical_RADDR_wire\ <= \N__33442\&\N__33742\&\N__33856\&\N__19438\&\N__32749\&\N__33973\&\N__18433\&\N__19615\&\N__35023\&\N__35374\&\N__33556\;
    \b2v_inst2.mem_mem_0_3_physical_WADDR_wire\ <= \N__33439\&\N__33745\&\N__33859\&\N__19435\&\N__32752\&\N__33976\&\N__18442\&\N__19630\&\N__35020\&\N__35377\&\N__33553\;
    \b2v_inst2.mem_mem_0_3_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \b2v_inst2.mem_mem_0_3_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__35462\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__35270\&'0'&'0'&'0';
    leds_c_13 <= \b2v_inst7.mem_mem_0_6_physical_RDATA_wire\(11);
    leds_c_12 <= \b2v_inst7.mem_mem_0_6_physical_RDATA_wire\(3);
    \b2v_inst7.mem_mem_0_6_physical_RADDR_wire\ <= \N__20080\&\N__15907\&\N__14101\&\N__14284\&\N__18655\&\N__19831\&\N__21526\&\N__20464\&\N__19948\&\N__14380\&\N__14191\;
    \b2v_inst7.mem_mem_0_6_physical_WADDR_wire\ <= \N__20077\&\N__15904\&\N__14098\&\N__14293\&\N__18652\&\N__19828\&\N__21523\&\N__20461\&\N__19945\&\N__14383\&\N__14194\;
    \b2v_inst7.mem_mem_0_6_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \b2v_inst7.mem_mem_0_6_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__24992\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__25034\&'0'&'0'&'0';
    \SYNTHESIZED_WIRE_1_5\ <= \b2v_inst8.mem_mem_0_2_physical_RDATA_wire\(11);
    \SYNTHESIZED_WIRE_1_4\ <= \b2v_inst8.mem_mem_0_2_physical_RDATA_wire\(3);
    \b2v_inst8.mem_mem_0_2_physical_RADDR_wire\ <= \N__36601\&\N__35746\&\N__38947\&\N__38734\&\N__38176\&\N__35524\&\N__36184\&\N__36397\&\N__35974\&\N__38488\&\N__39166\;
    \b2v_inst8.mem_mem_0_2_physical_WADDR_wire\ <= \N__36610\&\N__35749\&\N__38944\&\N__38731\&\N__38173\&\N__35527\&\N__36187\&\N__36400\&\N__35977\&\N__38485\&\N__39163\;
    \b2v_inst8.mem_mem_0_2_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \b2v_inst8.mem_mem_0_2_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__37316\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__33275\&'0'&'0'&'0';
    leds_c_7 <= \b2v_inst7.mem_mem_0_3_physical_RDATA_wire\(11);
    leds_c_6 <= \b2v_inst7.mem_mem_0_3_physical_RDATA_wire\(3);
    \b2v_inst7.mem_mem_0_3_physical_RADDR_wire\ <= \N__20116\&\N__15943\&\N__14137\&\N__14320\&\N__18691\&\N__19867\&\N__21562\&\N__20500\&\N__19984\&\N__14416\&\N__14227\;
    \b2v_inst7.mem_mem_0_3_physical_WADDR_wire\ <= \N__20113\&\N__15940\&\N__14134\&\N__14329\&\N__18688\&\N__19864\&\N__21559\&\N__20497\&\N__19981\&\N__14419\&\N__14230\;
    \b2v_inst7.mem_mem_0_3_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \b2v_inst7.mem_mem_0_3_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__23477\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__15443\&'0'&'0'&'0';
    leds_c_1 <= \b2v_inst7.mem_mem_0_0_physical_RDATA_wire\(11);
    leds_c_0 <= \b2v_inst7.mem_mem_0_0_physical_RDATA_wire\(3);
    \b2v_inst7.mem_mem_0_0_physical_RADDR_wire\ <= \N__20150\&\N__15977\&\N__14171\&\N__14356\&\N__18725\&\N__19901\&\N__21596\&\N__20534\&\N__20018\&\N__14452\&\N__14263\;
    \b2v_inst7.mem_mem_0_0_physical_WADDR_wire\ <= \N__20149\&\N__15976\&\N__14170\&\N__14360\&\N__18724\&\N__19900\&\N__21595\&\N__20533\&\N__20017\&\N__14453\&\N__14264\;
    \b2v_inst7.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \b2v_inst7.mem_mem_0_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__20858\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__20576\&'0'&'0'&'0';
    \SYNTHESIZED_WIRE_3_10\ <= \b2v_inst2.mem_mem_0_5_physical_RDATA_wire\(3);
    \b2v_inst2.mem_mem_0_5_physical_RADDR_wire\ <= \N__33418\&\N__33718\&\N__33832\&\N__19414\&\N__32725\&\N__33949\&\N__18409\&\N__19591\&\N__34999\&\N__35350\&\N__33532\;
    \b2v_inst2.mem_mem_0_5_physical_WADDR_wire\ <= \N__33415\&\N__33721\&\N__33835\&\N__19411\&\N__32728\&\N__33952\&\N__18418\&\N__19606\&\N__34996\&\N__35353\&\N__33529\;
    \b2v_inst2.mem_mem_0_5_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \b2v_inst2.mem_mem_0_5_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__33632\&'0'&'0'&'0';
    leds_c_11 <= \b2v_inst7.mem_mem_0_5_physical_RDATA_wire\(11);
    leds_c_10 <= \b2v_inst7.mem_mem_0_5_physical_RDATA_wire\(3);
    \b2v_inst7.mem_mem_0_5_physical_RADDR_wire\ <= \N__20092\&\N__15919\&\N__14113\&\N__14296\&\N__18667\&\N__19843\&\N__21538\&\N__20476\&\N__19960\&\N__14392\&\N__14203\;
    \b2v_inst7.mem_mem_0_5_physical_WADDR_wire\ <= \N__20089\&\N__15916\&\N__14110\&\N__14305\&\N__18664\&\N__19840\&\N__21535\&\N__20473\&\N__19957\&\N__14395\&\N__14206\;
    \b2v_inst7.mem_mem_0_5_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \b2v_inst7.mem_mem_0_5_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__25082\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__24926\&'0'&'0'&'0';

    \b2v_inst2.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \b2v_inst2.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \b2v_inst2.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \b2v_inst2.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \b2v_inst2.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \b2v_inst2.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__34435\,
            RE => \N__37212\,
            WCLKE => \N__21473\,
            WCLK => \N__34436\,
            WE => \N__37292\
        );

    \b2v_inst8.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \b2v_inst8.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \b2v_inst8.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \b2v_inst8.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \b2v_inst8.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \b2v_inst8.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__34376\,
            RE => \N__36996\,
            WCLKE => \N__21453\,
            WCLK => \N__34377\,
            WE => \N__36847\
        );

    \b2v_inst7.mem_mem_0_2_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \b2v_inst7.mem_mem_0_2_physical_RDATA_wire\,
            RADDR => \b2v_inst7.mem_mem_0_2_physical_RADDR_wire\,
            WADDR => \b2v_inst7.mem_mem_0_2_physical_WADDR_wire\,
            MASK => \b2v_inst7.mem_mem_0_2_physical_MASK_wire\,
            WDATA => \b2v_inst7.mem_mem_0_2_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__34486\,
            RE => \N__37231\,
            WCLKE => \N__21447\,
            WCLK => \N__34487\,
            WE => \N__37242\
        );

    \b2v_inst2.mem_mem_0_2_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \b2v_inst2.mem_mem_0_2_physical_RDATA_wire\,
            RADDR => \b2v_inst2.mem_mem_0_2_physical_RADDR_wire\,
            WADDR => \b2v_inst2.mem_mem_0_2_physical_WADDR_wire\,
            MASK => \b2v_inst2.mem_mem_0_2_physical_MASK_wire\,
            WDATA => \b2v_inst2.mem_mem_0_2_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__34400\,
            RE => \N__37129\,
            WCLKE => \N__21468\,
            WCLK => \N__34401\,
            WE => \N__37198\
        );

    \b2v_inst2.mem_mem_0_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \b2v_inst2.mem_mem_0_1_physical_RDATA_wire\,
            RADDR => \b2v_inst2.mem_mem_0_1_physical_RADDR_wire\,
            WADDR => \b2v_inst2.mem_mem_0_1_physical_WADDR_wire\,
            MASK => \b2v_inst2.mem_mem_0_1_physical_MASK_wire\,
            WDATA => \b2v_inst2.mem_mem_0_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__34419\,
            RE => \N__37256\,
            WCLKE => \N__21469\,
            WCLK => \N__34418\,
            WE => \N__37199\
        );

    \b2v_inst8.mem_mem_0_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \b2v_inst8.mem_mem_0_1_physical_RDATA_wire\,
            RADDR => \b2v_inst8.mem_mem_0_1_physical_RADDR_wire\,
            WADDR => \b2v_inst8.mem_mem_0_1_physical_WADDR_wire\,
            MASK => \b2v_inst8.mem_mem_0_1_physical_MASK_wire\,
            WDATA => \b2v_inst8.mem_mem_0_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__34389\,
            RE => \N__36836\,
            WCLKE => \N__21454\,
            WCLK => \N__34390\,
            WE => \N__36837\
        );

    \b2v_inst7.mem_mem_0_4_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \b2v_inst7.mem_mem_0_4_physical_RDATA_wire\,
            RADDR => \b2v_inst7.mem_mem_0_4_physical_RADDR_wire\,
            WADDR => \b2v_inst7.mem_mem_0_4_physical_WADDR_wire\,
            MASK => \b2v_inst7.mem_mem_0_4_physical_MASK_wire\,
            WDATA => \b2v_inst7.mem_mem_0_4_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__34520\,
            RE => \N__37213\,
            WCLKE => \N__21448\,
            WCLK => \N__34521\,
            WE => \N__37226\
        );

    \b2v_inst7.mem_mem_0_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \b2v_inst7.mem_mem_0_1_physical_RDATA_wire\,
            RADDR => \b2v_inst7.mem_mem_0_1_physical_RADDR_wire\,
            WADDR => \b2v_inst7.mem_mem_0_1_physical_WADDR_wire\,
            MASK => \b2v_inst7.mem_mem_0_1_physical_MASK_wire\,
            WDATA => \b2v_inst7.mem_mem_0_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__34504\,
            RE => \N__37286\,
            WCLKE => \N__21391\,
            WCLK => \N__34505\,
            WE => \N__37249\
        );

    \b2v_inst2.mem_mem_0_4_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \b2v_inst2.mem_mem_0_4_physical_RDATA_wire\,
            RADDR => \b2v_inst2.mem_mem_0_4_physical_RADDR_wire\,
            WADDR => \b2v_inst2.mem_mem_0_4_physical_WADDR_wire\,
            MASK => \b2v_inst2.mem_mem_0_4_physical_MASK_wire\,
            WDATA => \b2v_inst2.mem_mem_0_4_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__34374\,
            RE => \N__37014\,
            WCLKE => \N__21456\,
            WCLK => \N__34375\,
            WE => \N__37015\
        );

    \b2v_inst2.mem_mem_0_3_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \b2v_inst2.mem_mem_0_3_physical_RDATA_wire\,
            RADDR => \b2v_inst2.mem_mem_0_3_physical_RADDR_wire\,
            WADDR => \b2v_inst2.mem_mem_0_3_physical_WADDR_wire\,
            MASK => \b2v_inst2.mem_mem_0_3_physical_MASK_wire\,
            WDATA => \b2v_inst2.mem_mem_0_3_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__34387\,
            RE => \N__37112\,
            WCLKE => \N__21457\,
            WCLK => \N__34388\,
            WE => \N__37029\
        );

    \b2v_inst7.mem_mem_0_6_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \b2v_inst7.mem_mem_0_6_physical_RDATA_wire\,
            RADDR => \b2v_inst7.mem_mem_0_6_physical_RADDR_wire\,
            WADDR => \b2v_inst7.mem_mem_0_6_physical_WADDR_wire\,
            MASK => \b2v_inst7.mem_mem_0_6_physical_MASK_wire\,
            WDATA => \b2v_inst7.mem_mem_0_6_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__34528\,
            RE => \N__37282\,
            WCLKE => \N__21467\,
            WCLK => \N__34529\,
            WE => \N__37285\
        );

    \b2v_inst8.mem_mem_0_2_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \b2v_inst8.mem_mem_0_2_physical_RDATA_wire\,
            RADDR => \b2v_inst8.mem_mem_0_2_physical_RADDR_wire\,
            WADDR => \b2v_inst8.mem_mem_0_2_physical_WADDR_wire\,
            MASK => \b2v_inst8.mem_mem_0_2_physical_MASK_wire\,
            WDATA => \b2v_inst8.mem_mem_0_2_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__34402\,
            RE => \N__36921\,
            WCLKE => \N__21455\,
            WCLK => \N__34403\,
            WE => \N__37012\
        );

    \b2v_inst7.mem_mem_0_3_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \b2v_inst7.mem_mem_0_3_physical_RDATA_wire\,
            RADDR => \b2v_inst7.mem_mem_0_3_physical_RADDR_wire\,
            WADDR => \b2v_inst7.mem_mem_0_3_physical_WADDR_wire\,
            MASK => \b2v_inst7.mem_mem_0_3_physical_MASK_wire\,
            WDATA => \b2v_inst7.mem_mem_0_3_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__34506\,
            RE => \N__37160\,
            WCLKE => \N__21410\,
            WCLK => \N__34507\,
            WE => \N__37235\
        );

    \b2v_inst7.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \b2v_inst7.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \b2v_inst7.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \b2v_inst7.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \b2v_inst7.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \b2v_inst7.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__34518\,
            RE => \N__37287\,
            WCLKE => \N__21426\,
            WCLK => \N__34519\,
            WE => \N__37283\
        );

    \b2v_inst2.mem_mem_0_5_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \b2v_inst2.mem_mem_0_5_physical_RDATA_wire\,
            RADDR => \b2v_inst2.mem_mem_0_5_physical_RADDR_wire\,
            WADDR => \b2v_inst2.mem_mem_0_5_physical_WADDR_wire\,
            MASK => \b2v_inst2.mem_mem_0_5_physical_MASK_wire\,
            WDATA => \b2v_inst2.mem_mem_0_5_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__34371\,
            RE => \N__37013\,
            WCLKE => \N__21427\,
            WCLK => \N__34372\,
            WE => \N__36938\
        );

    \b2v_inst7.mem_mem_0_5_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \b2v_inst7.mem_mem_0_5_physical_RDATA_wire\,
            RADDR => \b2v_inst7.mem_mem_0_5_physical_RADDR_wire\,
            WADDR => \b2v_inst7.mem_mem_0_5_physical_WADDR_wire\,
            MASK => \b2v_inst7.mem_mem_0_5_physical_MASK_wire\,
            WDATA => \b2v_inst7.mem_mem_0_5_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__34526\,
            RE => \N__37227\,
            WCLKE => \N__21449\,
            WCLK => \N__34527\,
            WE => \N__37284\
        );

    \clk_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__39654\,
            GLOBALBUFFEROUTPUT => clk_c_g
        );

    \clk_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39656\,
            DIN => \N__39655\,
            DOUT => \N__39654\,
            PACKAGEPIN => clk_wire
        );

    \clk_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__39656\,
            PADOUT => \N__39655\,
            PADIN => \N__39654\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \leds_obuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39645\,
            DIN => \N__39644\,
            DOUT => \N__39643\,
            PACKAGEPIN => leds_wire(9)
        );

    \leds_obuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__39645\,
            PADOUT => \N__39644\,
            PADIN => \N__39643\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__26261\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \swit_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39636\,
            DIN => \N__39635\,
            DOUT => \N__39634\,
            PACKAGEPIN => swit_wire(0)
        );

    \swit_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__39636\,
            PADOUT => \N__39635\,
            PADIN => \N__39634\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => swit_c_0,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \leds_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39627\,
            DIN => \N__39626\,
            DOUT => \N__39625\,
            PACKAGEPIN => leds_wire(3)
        );

    \leds_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__39627\,
            PADOUT => \N__39626\,
            PADIN => \N__39625\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__23653\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \swit_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39618\,
            DIN => \N__39617\,
            DOUT => \N__39616\,
            PACKAGEPIN => swit_wire(6)
        );

    \swit_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__39618\,
            PADOUT => \N__39617\,
            PADIN => \N__39616\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => swit_c_6,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \leds_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39609\,
            DIN => \N__39608\,
            DOUT => \N__39607\,
            PACKAGEPIN => leds_wire(5)
        );

    \leds_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__39609\,
            PADOUT => \N__39608\,
            PADIN => \N__39607\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__17156\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \swit_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39600\,
            DIN => \N__39599\,
            DOUT => \N__39598\,
            PACKAGEPIN => swit_wire(8)
        );

    \swit_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__39600\,
            PADOUT => \N__39599\,
            PADIN => \N__39598\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => swit_c_8,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \swit_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39591\,
            DIN => \N__39590\,
            DOUT => \N__39589\,
            PACKAGEPIN => swit_wire(3)
        );

    \swit_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__39591\,
            PADOUT => \N__39590\,
            PADIN => \N__39589\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => swit_c_3,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \leds_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39582\,
            DIN => \N__39581\,
            DOUT => \N__39580\,
            PACKAGEPIN => leds_wire(0)
        );

    \leds_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__39582\,
            PADOUT => \N__39581\,
            PADIN => \N__39580\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__23404\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \leds_obuf_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39573\,
            DIN => \N__39572\,
            DOUT => \N__39571\,
            PACKAGEPIN => leds_wire(11)
        );

    \leds_obuf_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__39573\,
            PADOUT => \N__39572\,
            PADIN => \N__39571\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__17795\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \swit_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39564\,
            DIN => \N__39563\,
            DOUT => \N__39562\,
            PACKAGEPIN => swit_wire(4)
        );

    \swit_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__39564\,
            PADOUT => \N__39563\,
            PADIN => \N__39562\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => swit_c_4,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \leds_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39555\,
            DIN => \N__39554\,
            DOUT => \N__39553\,
            PACKAGEPIN => leds_wire(7)
        );

    \leds_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__39555\,
            PADOUT => \N__39554\,
            PADIN => \N__39553\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__17764\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \swit_ibuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39546\,
            DIN => \N__39545\,
            DOUT => \N__39544\,
            PACKAGEPIN => swit_wire(10)
        );

    \swit_ibuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__39546\,
            PADOUT => \N__39545\,
            PADIN => \N__39544\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => swit_c_10,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \uart_rx_i_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39537\,
            DIN => \N__39536\,
            DOUT => \N__39535\,
            PACKAGEPIN => uart_rx_i_wire
        );

    \uart_rx_i_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__39537\,
            PADOUT => \N__39536\,
            PADIN => \N__39535\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => uart_rx_i_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \leds_obuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39528\,
            DIN => \N__39527\,
            DOUT => \N__39526\,
            PACKAGEPIN => leds_wire(8)
        );

    \leds_obuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__39528\,
            PADOUT => \N__39527\,
            PADIN => \N__39526\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__24977\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \reset_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39519\,
            DIN => \N__39518\,
            DOUT => \N__39517\,
            PACKAGEPIN => reset_wire
        );

    \reset_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__39519\,
            PADOUT => \N__39518\,
            PADIN => \N__39517\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => reset_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \swit_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39510\,
            DIN => \N__39509\,
            DOUT => \N__39508\,
            PACKAGEPIN => swit_wire(1)
        );

    \swit_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__39510\,
            PADOUT => \N__39509\,
            PADIN => \N__39508\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => swit_c_1,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \leds_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39501\,
            DIN => \N__39500\,
            DOUT => \N__39499\,
            PACKAGEPIN => leds_wire(2)
        );

    \leds_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__39501\,
            PADOUT => \N__39500\,
            PADIN => \N__39499\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__23674\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \leds_obuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39492\,
            DIN => \N__39491\,
            DOUT => \N__39490\,
            PACKAGEPIN => leds_wire(13)
        );

    \leds_obuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__39492\,
            PADOUT => \N__39491\,
            PADIN => \N__39490\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__23332\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \swit_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39483\,
            DIN => \N__39482\,
            DOUT => \N__39481\,
            PACKAGEPIN => swit_wire(2)
        );

    \swit_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__39483\,
            PADOUT => \N__39482\,
            PADIN => \N__39481\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => swit_c_2,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \leds_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39474\,
            DIN => \N__39473\,
            DOUT => \N__39472\,
            PACKAGEPIN => leds_wire(1)
        );

    \leds_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__39474\,
            PADOUT => \N__39473\,
            PADIN => \N__39472\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__23372\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \leds_obuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39465\,
            DIN => \N__39464\,
            DOUT => \N__39463\,
            PACKAGEPIN => leds_wire(10)
        );

    \leds_obuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__39465\,
            PADOUT => \N__39464\,
            PADIN => \N__39463\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__17825\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \swit_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39456\,
            DIN => \N__39455\,
            DOUT => \N__39454\,
            PACKAGEPIN => swit_wire(7)
        );

    \swit_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__39456\,
            PADOUT => \N__39455\,
            PADIN => \N__39454\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => swit_c_7,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \leds_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39447\,
            DIN => \N__39446\,
            DOUT => \N__39445\,
            PACKAGEPIN => leds_wire(4)
        );

    \leds_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__39447\,
            PADOUT => \N__39446\,
            PADIN => \N__39445\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__17192\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \swit_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39438\,
            DIN => \N__39437\,
            DOUT => \N__39436\,
            PACKAGEPIN => swit_wire(9)
        );

    \swit_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__39438\,
            PADOUT => \N__39437\,
            PADIN => \N__39436\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => swit_c_9,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \uart_tx_o_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39429\,
            DIN => \N__39428\,
            DOUT => \N__39427\,
            PACKAGEPIN => uart_tx_o_wire
        );

    \uart_tx_o_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__39429\,
            PADOUT => \N__39428\,
            PADIN => \N__39427\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__26099\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \leds_obuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39420\,
            DIN => \N__39419\,
            DOUT => \N__39418\,
            PACKAGEPIN => leds_wire(12)
        );

    \leds_obuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__39420\,
            PADOUT => \N__39419\,
            PADIN => \N__39418\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__18875\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \swit_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39411\,
            DIN => \N__39410\,
            DOUT => \N__39409\,
            PACKAGEPIN => swit_wire(5)
        );

    \swit_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__39411\,
            PADOUT => \N__39410\,
            PADIN => \N__39409\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => swit_c_5,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \leds_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39402\,
            DIN => \N__39401\,
            DOUT => \N__39400\,
            PACKAGEPIN => leds_wire(6)
        );

    \leds_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__39402\,
            PADOUT => \N__39401\,
            PADIN => \N__39400\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__20432\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__9791\ : CascadeMux
    port map (
            O => \N__39383\,
            I => \N__39380\
        );

    \I__9790\ : InMux
    port map (
            O => \N__39380\,
            I => \N__39377\
        );

    \I__9789\ : LocalMux
    port map (
            O => \N__39377\,
            I => \N__39373\
        );

    \I__9788\ : InMux
    port map (
            O => \N__39376\,
            I => \N__39370\
        );

    \I__9787\ : Span4Mux_v
    port map (
            O => \N__39373\,
            I => \N__39366\
        );

    \I__9786\ : LocalMux
    port map (
            O => \N__39370\,
            I => \N__39363\
        );

    \I__9785\ : InMux
    port map (
            O => \N__39369\,
            I => \N__39360\
        );

    \I__9784\ : Span4Mux_h
    port map (
            O => \N__39366\,
            I => \N__39356\
        );

    \I__9783\ : Span4Mux_h
    port map (
            O => \N__39363\,
            I => \N__39351\
        );

    \I__9782\ : LocalMux
    port map (
            O => \N__39360\,
            I => \N__39351\
        );

    \I__9781\ : InMux
    port map (
            O => \N__39359\,
            I => \N__39346\
        );

    \I__9780\ : Span4Mux_h
    port map (
            O => \N__39356\,
            I => \N__39343\
        );

    \I__9779\ : Span4Mux_v
    port map (
            O => \N__39351\,
            I => \N__39340\
        );

    \I__9778\ : InMux
    port map (
            O => \N__39350\,
            I => \N__39337\
        );

    \I__9777\ : InMux
    port map (
            O => \N__39349\,
            I => \N__39334\
        );

    \I__9776\ : LocalMux
    port map (
            O => \N__39346\,
            I => \b2v_inst.dir_energiaZ0Z_0\
        );

    \I__9775\ : Odrv4
    port map (
            O => \N__39343\,
            I => \b2v_inst.dir_energiaZ0Z_0\
        );

    \I__9774\ : Odrv4
    port map (
            O => \N__39340\,
            I => \b2v_inst.dir_energiaZ0Z_0\
        );

    \I__9773\ : LocalMux
    port map (
            O => \N__39337\,
            I => \b2v_inst.dir_energiaZ0Z_0\
        );

    \I__9772\ : LocalMux
    port map (
            O => \N__39334\,
            I => \b2v_inst.dir_energiaZ0Z_0\
        );

    \I__9771\ : InMux
    port map (
            O => \N__39323\,
            I => \N__39319\
        );

    \I__9770\ : InMux
    port map (
            O => \N__39322\,
            I => \N__39313\
        );

    \I__9769\ : LocalMux
    port map (
            O => \N__39319\,
            I => \N__39310\
        );

    \I__9768\ : InMux
    port map (
            O => \N__39318\,
            I => \N__39307\
        );

    \I__9767\ : InMux
    port map (
            O => \N__39317\,
            I => \N__39300\
        );

    \I__9766\ : CascadeMux
    port map (
            O => \N__39316\,
            I => \N__39297\
        );

    \I__9765\ : LocalMux
    port map (
            O => \N__39313\,
            I => \N__39294\
        );

    \I__9764\ : Span4Mux_v
    port map (
            O => \N__39310\,
            I => \N__39289\
        );

    \I__9763\ : LocalMux
    port map (
            O => \N__39307\,
            I => \N__39289\
        );

    \I__9762\ : InMux
    port map (
            O => \N__39306\,
            I => \N__39286\
        );

    \I__9761\ : InMux
    port map (
            O => \N__39305\,
            I => \N__39283\
        );

    \I__9760\ : InMux
    port map (
            O => \N__39304\,
            I => \N__39280\
        );

    \I__9759\ : InMux
    port map (
            O => \N__39303\,
            I => \N__39277\
        );

    \I__9758\ : LocalMux
    port map (
            O => \N__39300\,
            I => \N__39274\
        );

    \I__9757\ : InMux
    port map (
            O => \N__39297\,
            I => \N__39270\
        );

    \I__9756\ : Span4Mux_v
    port map (
            O => \N__39294\,
            I => \N__39267\
        );

    \I__9755\ : Span4Mux_v
    port map (
            O => \N__39289\,
            I => \N__39264\
        );

    \I__9754\ : LocalMux
    port map (
            O => \N__39286\,
            I => \N__39261\
        );

    \I__9753\ : LocalMux
    port map (
            O => \N__39283\,
            I => \N__39258\
        );

    \I__9752\ : LocalMux
    port map (
            O => \N__39280\,
            I => \N__39255\
        );

    \I__9751\ : LocalMux
    port map (
            O => \N__39277\,
            I => \N__39252\
        );

    \I__9750\ : Span4Mux_h
    port map (
            O => \N__39274\,
            I => \N__39249\
        );

    \I__9749\ : InMux
    port map (
            O => \N__39273\,
            I => \N__39246\
        );

    \I__9748\ : LocalMux
    port map (
            O => \N__39270\,
            I => \N__39243\
        );

    \I__9747\ : Span4Mux_h
    port map (
            O => \N__39267\,
            I => \N__39237\
        );

    \I__9746\ : Span4Mux_h
    port map (
            O => \N__39264\,
            I => \N__39237\
        );

    \I__9745\ : Span4Mux_v
    port map (
            O => \N__39261\,
            I => \N__39228\
        );

    \I__9744\ : Span4Mux_v
    port map (
            O => \N__39258\,
            I => \N__39228\
        );

    \I__9743\ : Span4Mux_h
    port map (
            O => \N__39255\,
            I => \N__39228\
        );

    \I__9742\ : Span4Mux_v
    port map (
            O => \N__39252\,
            I => \N__39228\
        );

    \I__9741\ : Sp12to4
    port map (
            O => \N__39249\,
            I => \N__39223\
        );

    \I__9740\ : LocalMux
    port map (
            O => \N__39246\,
            I => \N__39220\
        );

    \I__9739\ : Span4Mux_h
    port map (
            O => \N__39243\,
            I => \N__39217\
        );

    \I__9738\ : InMux
    port map (
            O => \N__39242\,
            I => \N__39214\
        );

    \I__9737\ : Span4Mux_v
    port map (
            O => \N__39237\,
            I => \N__39209\
        );

    \I__9736\ : Span4Mux_h
    port map (
            O => \N__39228\,
            I => \N__39209\
        );

    \I__9735\ : InMux
    port map (
            O => \N__39227\,
            I => \N__39204\
        );

    \I__9734\ : InMux
    port map (
            O => \N__39226\,
            I => \N__39204\
        );

    \I__9733\ : Span12Mux_v
    port map (
            O => \N__39223\,
            I => \N__39199\
        );

    \I__9732\ : Span12Mux_h
    port map (
            O => \N__39220\,
            I => \N__39199\
        );

    \I__9731\ : Odrv4
    port map (
            O => \N__39217\,
            I => \b2v_inst.indiceZ0Z_0\
        );

    \I__9730\ : LocalMux
    port map (
            O => \N__39214\,
            I => \b2v_inst.indiceZ0Z_0\
        );

    \I__9729\ : Odrv4
    port map (
            O => \N__39209\,
            I => \b2v_inst.indiceZ0Z_0\
        );

    \I__9728\ : LocalMux
    port map (
            O => \N__39204\,
            I => \b2v_inst.indiceZ0Z_0\
        );

    \I__9727\ : Odrv12
    port map (
            O => \N__39199\,
            I => \b2v_inst.indiceZ0Z_0\
        );

    \I__9726\ : CascadeMux
    port map (
            O => \N__39188\,
            I => \N__39184\
        );

    \I__9725\ : CascadeMux
    port map (
            O => \N__39187\,
            I => \N__39181\
        );

    \I__9724\ : CascadeBuf
    port map (
            O => \N__39184\,
            I => \N__39178\
        );

    \I__9723\ : CascadeBuf
    port map (
            O => \N__39181\,
            I => \N__39175\
        );

    \I__9722\ : CascadeMux
    port map (
            O => \N__39178\,
            I => \N__39172\
        );

    \I__9721\ : CascadeMux
    port map (
            O => \N__39175\,
            I => \N__39169\
        );

    \I__9720\ : CascadeBuf
    port map (
            O => \N__39172\,
            I => \N__39166\
        );

    \I__9719\ : CascadeBuf
    port map (
            O => \N__39169\,
            I => \N__39163\
        );

    \I__9718\ : CascadeMux
    port map (
            O => \N__39166\,
            I => \N__39160\
        );

    \I__9717\ : CascadeMux
    port map (
            O => \N__39163\,
            I => \N__39157\
        );

    \I__9716\ : InMux
    port map (
            O => \N__39160\,
            I => \N__39154\
        );

    \I__9715\ : InMux
    port map (
            O => \N__39157\,
            I => \N__39151\
        );

    \I__9714\ : LocalMux
    port map (
            O => \N__39154\,
            I => \N_360_i\
        );

    \I__9713\ : LocalMux
    port map (
            O => \N__39151\,
            I => \N_360_i\
        );

    \I__9712\ : InMux
    port map (
            O => \N__39146\,
            I => \N__39143\
        );

    \I__9711\ : LocalMux
    port map (
            O => \N__39143\,
            I => \N__39140\
        );

    \I__9710\ : Span4Mux_h
    port map (
            O => \N__39140\,
            I => \N__39135\
        );

    \I__9709\ : InMux
    port map (
            O => \N__39139\,
            I => \N__39132\
        );

    \I__9708\ : InMux
    port map (
            O => \N__39138\,
            I => \N__39129\
        );

    \I__9707\ : Span4Mux_h
    port map (
            O => \N__39135\,
            I => \N__39124\
        );

    \I__9706\ : LocalMux
    port map (
            O => \N__39132\,
            I => \N__39124\
        );

    \I__9705\ : LocalMux
    port map (
            O => \N__39129\,
            I => \N__39119\
        );

    \I__9704\ : Span4Mux_h
    port map (
            O => \N__39124\,
            I => \N__39116\
        );

    \I__9703\ : InMux
    port map (
            O => \N__39123\,
            I => \N__39113\
        );

    \I__9702\ : InMux
    port map (
            O => \N__39122\,
            I => \N__39110\
        );

    \I__9701\ : Odrv4
    port map (
            O => \N__39119\,
            I => \b2v_inst.dir_energiaZ0Z_8\
        );

    \I__9700\ : Odrv4
    port map (
            O => \N__39116\,
            I => \b2v_inst.dir_energiaZ0Z_8\
        );

    \I__9699\ : LocalMux
    port map (
            O => \N__39113\,
            I => \b2v_inst.dir_energiaZ0Z_8\
        );

    \I__9698\ : LocalMux
    port map (
            O => \N__39110\,
            I => \b2v_inst.dir_energiaZ0Z_8\
        );

    \I__9697\ : CascadeMux
    port map (
            O => \N__39101\,
            I => \N__39097\
        );

    \I__9696\ : CascadeMux
    port map (
            O => \N__39100\,
            I => \N__39094\
        );

    \I__9695\ : InMux
    port map (
            O => \N__39097\,
            I => \N__39091\
        );

    \I__9694\ : InMux
    port map (
            O => \N__39094\,
            I => \N__39088\
        );

    \I__9693\ : LocalMux
    port map (
            O => \N__39091\,
            I => \N__39085\
        );

    \I__9692\ : LocalMux
    port map (
            O => \N__39088\,
            I => \N__39082\
        );

    \I__9691\ : Span4Mux_v
    port map (
            O => \N__39085\,
            I => \N__39076\
        );

    \I__9690\ : Span4Mux_v
    port map (
            O => \N__39082\,
            I => \N__39073\
        );

    \I__9689\ : InMux
    port map (
            O => \N__39081\,
            I => \N__39070\
        );

    \I__9688\ : InMux
    port map (
            O => \N__39080\,
            I => \N__39065\
        );

    \I__9687\ : InMux
    port map (
            O => \N__39079\,
            I => \N__39062\
        );

    \I__9686\ : Span4Mux_v
    port map (
            O => \N__39076\,
            I => \N__39059\
        );

    \I__9685\ : Span4Mux_v
    port map (
            O => \N__39073\,
            I => \N__39053\
        );

    \I__9684\ : LocalMux
    port map (
            O => \N__39070\,
            I => \N__39053\
        );

    \I__9683\ : InMux
    port map (
            O => \N__39069\,
            I => \N__39050\
        );

    \I__9682\ : InMux
    port map (
            O => \N__39068\,
            I => \N__39046\
        );

    \I__9681\ : LocalMux
    port map (
            O => \N__39065\,
            I => \N__39041\
        );

    \I__9680\ : LocalMux
    port map (
            O => \N__39062\,
            I => \N__39041\
        );

    \I__9679\ : Span4Mux_v
    port map (
            O => \N__39059\,
            I => \N__39038\
        );

    \I__9678\ : InMux
    port map (
            O => \N__39058\,
            I => \N__39035\
        );

    \I__9677\ : Span4Mux_v
    port map (
            O => \N__39053\,
            I => \N__39031\
        );

    \I__9676\ : LocalMux
    port map (
            O => \N__39050\,
            I => \N__39028\
        );

    \I__9675\ : InMux
    port map (
            O => \N__39049\,
            I => \N__39023\
        );

    \I__9674\ : LocalMux
    port map (
            O => \N__39046\,
            I => \N__39018\
        );

    \I__9673\ : Span4Mux_v
    port map (
            O => \N__39041\,
            I => \N__39018\
        );

    \I__9672\ : Span4Mux_v
    port map (
            O => \N__39038\,
            I => \N__39013\
        );

    \I__9671\ : LocalMux
    port map (
            O => \N__39035\,
            I => \N__39013\
        );

    \I__9670\ : InMux
    port map (
            O => \N__39034\,
            I => \N__39010\
        );

    \I__9669\ : Span4Mux_h
    port map (
            O => \N__39031\,
            I => \N__39007\
        );

    \I__9668\ : Span4Mux_v
    port map (
            O => \N__39028\,
            I => \N__39004\
        );

    \I__9667\ : InMux
    port map (
            O => \N__39027\,
            I => \N__39001\
        );

    \I__9666\ : InMux
    port map (
            O => \N__39026\,
            I => \N__38998\
        );

    \I__9665\ : LocalMux
    port map (
            O => \N__39023\,
            I => \N__38995\
        );

    \I__9664\ : Span4Mux_h
    port map (
            O => \N__39018\,
            I => \N__38992\
        );

    \I__9663\ : Span4Mux_h
    port map (
            O => \N__39013\,
            I => \N__38987\
        );

    \I__9662\ : LocalMux
    port map (
            O => \N__39010\,
            I => \N__38987\
        );

    \I__9661\ : Span4Mux_h
    port map (
            O => \N__39007\,
            I => \N__38980\
        );

    \I__9660\ : Span4Mux_h
    port map (
            O => \N__39004\,
            I => \N__38980\
        );

    \I__9659\ : LocalMux
    port map (
            O => \N__39001\,
            I => \N__38980\
        );

    \I__9658\ : LocalMux
    port map (
            O => \N__38998\,
            I => \b2v_inst.indiceZ0Z_8\
        );

    \I__9657\ : Odrv4
    port map (
            O => \N__38995\,
            I => \b2v_inst.indiceZ0Z_8\
        );

    \I__9656\ : Odrv4
    port map (
            O => \N__38992\,
            I => \b2v_inst.indiceZ0Z_8\
        );

    \I__9655\ : Odrv4
    port map (
            O => \N__38987\,
            I => \b2v_inst.indiceZ0Z_8\
        );

    \I__9654\ : Odrv4
    port map (
            O => \N__38980\,
            I => \b2v_inst.indiceZ0Z_8\
        );

    \I__9653\ : CascadeMux
    port map (
            O => \N__38969\,
            I => \N__38965\
        );

    \I__9652\ : CascadeMux
    port map (
            O => \N__38968\,
            I => \N__38962\
        );

    \I__9651\ : CascadeBuf
    port map (
            O => \N__38965\,
            I => \N__38959\
        );

    \I__9650\ : CascadeBuf
    port map (
            O => \N__38962\,
            I => \N__38956\
        );

    \I__9649\ : CascadeMux
    port map (
            O => \N__38959\,
            I => \N__38953\
        );

    \I__9648\ : CascadeMux
    port map (
            O => \N__38956\,
            I => \N__38950\
        );

    \I__9647\ : CascadeBuf
    port map (
            O => \N__38953\,
            I => \N__38947\
        );

    \I__9646\ : CascadeBuf
    port map (
            O => \N__38950\,
            I => \N__38944\
        );

    \I__9645\ : CascadeMux
    port map (
            O => \N__38947\,
            I => \N__38941\
        );

    \I__9644\ : CascadeMux
    port map (
            O => \N__38944\,
            I => \N__38938\
        );

    \I__9643\ : InMux
    port map (
            O => \N__38941\,
            I => \N__38935\
        );

    \I__9642\ : InMux
    port map (
            O => \N__38938\,
            I => \N__38932\
        );

    \I__9641\ : LocalMux
    port map (
            O => \N__38935\,
            I => \N_443_i\
        );

    \I__9640\ : LocalMux
    port map (
            O => \N__38932\,
            I => \N_443_i\
        );

    \I__9639\ : CascadeMux
    port map (
            O => \N__38927\,
            I => \N__38924\
        );

    \I__9638\ : InMux
    port map (
            O => \N__38924\,
            I => \N__38921\
        );

    \I__9637\ : LocalMux
    port map (
            O => \N__38921\,
            I => \N__38918\
        );

    \I__9636\ : Span4Mux_v
    port map (
            O => \N__38918\,
            I => \N__38914\
        );

    \I__9635\ : InMux
    port map (
            O => \N__38917\,
            I => \N__38911\
        );

    \I__9634\ : Span4Mux_h
    port map (
            O => \N__38914\,
            I => \N__38906\
        );

    \I__9633\ : LocalMux
    port map (
            O => \N__38911\,
            I => \N__38902\
        );

    \I__9632\ : CascadeMux
    port map (
            O => \N__38910\,
            I => \N__38899\
        );

    \I__9631\ : CascadeMux
    port map (
            O => \N__38909\,
            I => \N__38896\
        );

    \I__9630\ : Span4Mux_h
    port map (
            O => \N__38906\,
            I => \N__38893\
        );

    \I__9629\ : InMux
    port map (
            O => \N__38905\,
            I => \N__38890\
        );

    \I__9628\ : Span4Mux_h
    port map (
            O => \N__38902\,
            I => \N__38887\
        );

    \I__9627\ : InMux
    port map (
            O => \N__38899\,
            I => \N__38884\
        );

    \I__9626\ : InMux
    port map (
            O => \N__38896\,
            I => \N__38881\
        );

    \I__9625\ : Odrv4
    port map (
            O => \N__38893\,
            I => \b2v_inst.dir_energiaZ0Z_7\
        );

    \I__9624\ : LocalMux
    port map (
            O => \N__38890\,
            I => \b2v_inst.dir_energiaZ0Z_7\
        );

    \I__9623\ : Odrv4
    port map (
            O => \N__38887\,
            I => \b2v_inst.dir_energiaZ0Z_7\
        );

    \I__9622\ : LocalMux
    port map (
            O => \N__38884\,
            I => \b2v_inst.dir_energiaZ0Z_7\
        );

    \I__9621\ : LocalMux
    port map (
            O => \N__38881\,
            I => \b2v_inst.dir_energiaZ0Z_7\
        );

    \I__9620\ : InMux
    port map (
            O => \N__38870\,
            I => \N__38867\
        );

    \I__9619\ : LocalMux
    port map (
            O => \N__38867\,
            I => \N__38863\
        );

    \I__9618\ : InMux
    port map (
            O => \N__38866\,
            I => \N__38857\
        );

    \I__9617\ : Span4Mux_v
    port map (
            O => \N__38863\,
            I => \N__38854\
        );

    \I__9616\ : CascadeMux
    port map (
            O => \N__38862\,
            I => \N__38851\
        );

    \I__9615\ : InMux
    port map (
            O => \N__38861\,
            I => \N__38848\
        );

    \I__9614\ : CascadeMux
    port map (
            O => \N__38860\,
            I => \N__38844\
        );

    \I__9613\ : LocalMux
    port map (
            O => \N__38857\,
            I => \N__38840\
        );

    \I__9612\ : Sp12to4
    port map (
            O => \N__38854\,
            I => \N__38837\
        );

    \I__9611\ : InMux
    port map (
            O => \N__38851\,
            I => \N__38833\
        );

    \I__9610\ : LocalMux
    port map (
            O => \N__38848\,
            I => \N__38830\
        );

    \I__9609\ : InMux
    port map (
            O => \N__38847\,
            I => \N__38825\
        );

    \I__9608\ : InMux
    port map (
            O => \N__38844\,
            I => \N__38822\
        );

    \I__9607\ : InMux
    port map (
            O => \N__38843\,
            I => \N__38819\
        );

    \I__9606\ : Span12Mux_h
    port map (
            O => \N__38840\,
            I => \N__38814\
        );

    \I__9605\ : Span12Mux_h
    port map (
            O => \N__38837\,
            I => \N__38814\
        );

    \I__9604\ : InMux
    port map (
            O => \N__38836\,
            I => \N__38811\
        );

    \I__9603\ : LocalMux
    port map (
            O => \N__38833\,
            I => \N__38808\
        );

    \I__9602\ : Span4Mux_v
    port map (
            O => \N__38830\,
            I => \N__38805\
        );

    \I__9601\ : InMux
    port map (
            O => \N__38829\,
            I => \N__38802\
        );

    \I__9600\ : InMux
    port map (
            O => \N__38828\,
            I => \N__38799\
        );

    \I__9599\ : LocalMux
    port map (
            O => \N__38825\,
            I => \N__38794\
        );

    \I__9598\ : LocalMux
    port map (
            O => \N__38822\,
            I => \N__38794\
        );

    \I__9597\ : LocalMux
    port map (
            O => \N__38819\,
            I => \N__38790\
        );

    \I__9596\ : Span12Mux_v
    port map (
            O => \N__38814\,
            I => \N__38785\
        );

    \I__9595\ : LocalMux
    port map (
            O => \N__38811\,
            I => \N__38785\
        );

    \I__9594\ : Span4Mux_v
    port map (
            O => \N__38808\,
            I => \N__38782\
        );

    \I__9593\ : Span4Mux_h
    port map (
            O => \N__38805\,
            I => \N__38779\
        );

    \I__9592\ : LocalMux
    port map (
            O => \N__38802\,
            I => \N__38772\
        );

    \I__9591\ : LocalMux
    port map (
            O => \N__38799\,
            I => \N__38772\
        );

    \I__9590\ : Span4Mux_v
    port map (
            O => \N__38794\,
            I => \N__38772\
        );

    \I__9589\ : InMux
    port map (
            O => \N__38793\,
            I => \N__38769\
        );

    \I__9588\ : Odrv12
    port map (
            O => \N__38790\,
            I => \b2v_inst.indiceZ0Z_7\
        );

    \I__9587\ : Odrv12
    port map (
            O => \N__38785\,
            I => \b2v_inst.indiceZ0Z_7\
        );

    \I__9586\ : Odrv4
    port map (
            O => \N__38782\,
            I => \b2v_inst.indiceZ0Z_7\
        );

    \I__9585\ : Odrv4
    port map (
            O => \N__38779\,
            I => \b2v_inst.indiceZ0Z_7\
        );

    \I__9584\ : Odrv4
    port map (
            O => \N__38772\,
            I => \b2v_inst.indiceZ0Z_7\
        );

    \I__9583\ : LocalMux
    port map (
            O => \N__38769\,
            I => \b2v_inst.indiceZ0Z_7\
        );

    \I__9582\ : CascadeMux
    port map (
            O => \N__38756\,
            I => \N__38752\
        );

    \I__9581\ : CascadeMux
    port map (
            O => \N__38755\,
            I => \N__38749\
        );

    \I__9580\ : CascadeBuf
    port map (
            O => \N__38752\,
            I => \N__38746\
        );

    \I__9579\ : CascadeBuf
    port map (
            O => \N__38749\,
            I => \N__38743\
        );

    \I__9578\ : CascadeMux
    port map (
            O => \N__38746\,
            I => \N__38740\
        );

    \I__9577\ : CascadeMux
    port map (
            O => \N__38743\,
            I => \N__38737\
        );

    \I__9576\ : CascadeBuf
    port map (
            O => \N__38740\,
            I => \N__38734\
        );

    \I__9575\ : CascadeBuf
    port map (
            O => \N__38737\,
            I => \N__38731\
        );

    \I__9574\ : CascadeMux
    port map (
            O => \N__38734\,
            I => \N__38728\
        );

    \I__9573\ : CascadeMux
    port map (
            O => \N__38731\,
            I => \N__38725\
        );

    \I__9572\ : InMux
    port map (
            O => \N__38728\,
            I => \N__38722\
        );

    \I__9571\ : InMux
    port map (
            O => \N__38725\,
            I => \N__38719\
        );

    \I__9570\ : LocalMux
    port map (
            O => \N__38722\,
            I => \N_353_i\
        );

    \I__9569\ : LocalMux
    port map (
            O => \N__38719\,
            I => \N_353_i\
        );

    \I__9568\ : CascadeMux
    port map (
            O => \N__38714\,
            I => \N__38711\
        );

    \I__9567\ : InMux
    port map (
            O => \N__38711\,
            I => \N__38708\
        );

    \I__9566\ : LocalMux
    port map (
            O => \N__38708\,
            I => \N__38704\
        );

    \I__9565\ : InMux
    port map (
            O => \N__38707\,
            I => \N__38701\
        );

    \I__9564\ : Span4Mux_v
    port map (
            O => \N__38704\,
            I => \N__38698\
        );

    \I__9563\ : LocalMux
    port map (
            O => \N__38701\,
            I => \N__38694\
        );

    \I__9562\ : Sp12to4
    port map (
            O => \N__38698\,
            I => \N__38689\
        );

    \I__9561\ : InMux
    port map (
            O => \N__38697\,
            I => \N__38686\
        );

    \I__9560\ : Span4Mux_h
    port map (
            O => \N__38694\,
            I => \N__38683\
        );

    \I__9559\ : InMux
    port map (
            O => \N__38693\,
            I => \N__38680\
        );

    \I__9558\ : InMux
    port map (
            O => \N__38692\,
            I => \N__38677\
        );

    \I__9557\ : Odrv12
    port map (
            O => \N__38689\,
            I => \b2v_inst.dir_energiaZ0Z_1\
        );

    \I__9556\ : LocalMux
    port map (
            O => \N__38686\,
            I => \b2v_inst.dir_energiaZ0Z_1\
        );

    \I__9555\ : Odrv4
    port map (
            O => \N__38683\,
            I => \b2v_inst.dir_energiaZ0Z_1\
        );

    \I__9554\ : LocalMux
    port map (
            O => \N__38680\,
            I => \b2v_inst.dir_energiaZ0Z_1\
        );

    \I__9553\ : LocalMux
    port map (
            O => \N__38677\,
            I => \b2v_inst.dir_energiaZ0Z_1\
        );

    \I__9552\ : InMux
    port map (
            O => \N__38666\,
            I => \N__38661\
        );

    \I__9551\ : InMux
    port map (
            O => \N__38665\,
            I => \N__38657\
        );

    \I__9550\ : CascadeMux
    port map (
            O => \N__38664\,
            I => \N__38653\
        );

    \I__9549\ : LocalMux
    port map (
            O => \N__38661\,
            I => \N__38650\
        );

    \I__9548\ : InMux
    port map (
            O => \N__38660\,
            I => \N__38647\
        );

    \I__9547\ : LocalMux
    port map (
            O => \N__38657\,
            I => \N__38643\
        );

    \I__9546\ : InMux
    port map (
            O => \N__38656\,
            I => \N__38637\
        );

    \I__9545\ : InMux
    port map (
            O => \N__38653\,
            I => \N__38634\
        );

    \I__9544\ : Span4Mux_v
    port map (
            O => \N__38650\,
            I => \N__38629\
        );

    \I__9543\ : LocalMux
    port map (
            O => \N__38647\,
            I => \N__38629\
        );

    \I__9542\ : InMux
    port map (
            O => \N__38646\,
            I => \N__38626\
        );

    \I__9541\ : Span4Mux_v
    port map (
            O => \N__38643\,
            I => \N__38622\
        );

    \I__9540\ : InMux
    port map (
            O => \N__38642\,
            I => \N__38619\
        );

    \I__9539\ : InMux
    port map (
            O => \N__38641\,
            I => \N__38616\
        );

    \I__9538\ : InMux
    port map (
            O => \N__38640\,
            I => \N__38613\
        );

    \I__9537\ : LocalMux
    port map (
            O => \N__38637\,
            I => \N__38610\
        );

    \I__9536\ : LocalMux
    port map (
            O => \N__38634\,
            I => \N__38607\
        );

    \I__9535\ : Span4Mux_v
    port map (
            O => \N__38629\,
            I => \N__38604\
        );

    \I__9534\ : LocalMux
    port map (
            O => \N__38626\,
            I => \N__38600\
        );

    \I__9533\ : InMux
    port map (
            O => \N__38625\,
            I => \N__38597\
        );

    \I__9532\ : Span4Mux_v
    port map (
            O => \N__38622\,
            I => \N__38594\
        );

    \I__9531\ : LocalMux
    port map (
            O => \N__38619\,
            I => \N__38591\
        );

    \I__9530\ : LocalMux
    port map (
            O => \N__38616\,
            I => \N__38588\
        );

    \I__9529\ : LocalMux
    port map (
            O => \N__38613\,
            I => \N__38584\
        );

    \I__9528\ : Span4Mux_v
    port map (
            O => \N__38610\,
            I => \N__38579\
        );

    \I__9527\ : Span4Mux_v
    port map (
            O => \N__38607\,
            I => \N__38579\
        );

    \I__9526\ : Sp12to4
    port map (
            O => \N__38604\,
            I => \N__38576\
        );

    \I__9525\ : CascadeMux
    port map (
            O => \N__38603\,
            I => \N__38570\
        );

    \I__9524\ : Span4Mux_v
    port map (
            O => \N__38600\,
            I => \N__38567\
        );

    \I__9523\ : LocalMux
    port map (
            O => \N__38597\,
            I => \N__38564\
        );

    \I__9522\ : Span4Mux_v
    port map (
            O => \N__38594\,
            I => \N__38559\
        );

    \I__9521\ : Span4Mux_h
    port map (
            O => \N__38591\,
            I => \N__38559\
        );

    \I__9520\ : Span4Mux_v
    port map (
            O => \N__38588\,
            I => \N__38556\
        );

    \I__9519\ : InMux
    port map (
            O => \N__38587\,
            I => \N__38553\
        );

    \I__9518\ : Span4Mux_v
    port map (
            O => \N__38584\,
            I => \N__38548\
        );

    \I__9517\ : Span4Mux_h
    port map (
            O => \N__38579\,
            I => \N__38548\
        );

    \I__9516\ : Span12Mux_h
    port map (
            O => \N__38576\,
            I => \N__38545\
        );

    \I__9515\ : InMux
    port map (
            O => \N__38575\,
            I => \N__38540\
        );

    \I__9514\ : InMux
    port map (
            O => \N__38574\,
            I => \N__38540\
        );

    \I__9513\ : InMux
    port map (
            O => \N__38573\,
            I => \N__38537\
        );

    \I__9512\ : InMux
    port map (
            O => \N__38570\,
            I => \N__38534\
        );

    \I__9511\ : Span4Mux_h
    port map (
            O => \N__38567\,
            I => \N__38523\
        );

    \I__9510\ : Span4Mux_v
    port map (
            O => \N__38564\,
            I => \N__38523\
        );

    \I__9509\ : Span4Mux_v
    port map (
            O => \N__38559\,
            I => \N__38523\
        );

    \I__9508\ : Span4Mux_h
    port map (
            O => \N__38556\,
            I => \N__38523\
        );

    \I__9507\ : LocalMux
    port map (
            O => \N__38553\,
            I => \N__38523\
        );

    \I__9506\ : Odrv4
    port map (
            O => \N__38548\,
            I => \b2v_inst.indiceZ0Z_1\
        );

    \I__9505\ : Odrv12
    port map (
            O => \N__38545\,
            I => \b2v_inst.indiceZ0Z_1\
        );

    \I__9504\ : LocalMux
    port map (
            O => \N__38540\,
            I => \b2v_inst.indiceZ0Z_1\
        );

    \I__9503\ : LocalMux
    port map (
            O => \N__38537\,
            I => \b2v_inst.indiceZ0Z_1\
        );

    \I__9502\ : LocalMux
    port map (
            O => \N__38534\,
            I => \b2v_inst.indiceZ0Z_1\
        );

    \I__9501\ : Odrv4
    port map (
            O => \N__38523\,
            I => \b2v_inst.indiceZ0Z_1\
        );

    \I__9500\ : CascadeMux
    port map (
            O => \N__38510\,
            I => \N__38506\
        );

    \I__9499\ : CascadeMux
    port map (
            O => \N__38509\,
            I => \N__38503\
        );

    \I__9498\ : CascadeBuf
    port map (
            O => \N__38506\,
            I => \N__38500\
        );

    \I__9497\ : CascadeBuf
    port map (
            O => \N__38503\,
            I => \N__38497\
        );

    \I__9496\ : CascadeMux
    port map (
            O => \N__38500\,
            I => \N__38494\
        );

    \I__9495\ : CascadeMux
    port map (
            O => \N__38497\,
            I => \N__38491\
        );

    \I__9494\ : CascadeBuf
    port map (
            O => \N__38494\,
            I => \N__38488\
        );

    \I__9493\ : CascadeBuf
    port map (
            O => \N__38491\,
            I => \N__38485\
        );

    \I__9492\ : CascadeMux
    port map (
            O => \N__38488\,
            I => \N__38482\
        );

    \I__9491\ : CascadeMux
    port map (
            O => \N__38485\,
            I => \N__38479\
        );

    \I__9490\ : InMux
    port map (
            O => \N__38482\,
            I => \N__38476\
        );

    \I__9489\ : InMux
    port map (
            O => \N__38479\,
            I => \N__38473\
        );

    \I__9488\ : LocalMux
    port map (
            O => \N__38476\,
            I => \N_359_i\
        );

    \I__9487\ : LocalMux
    port map (
            O => \N__38473\,
            I => \N_359_i\
        );

    \I__9486\ : InMux
    port map (
            O => \N__38468\,
            I => \N__38447\
        );

    \I__9485\ : InMux
    port map (
            O => \N__38467\,
            I => \N__38447\
        );

    \I__9484\ : InMux
    port map (
            O => \N__38466\,
            I => \N__38447\
        );

    \I__9483\ : InMux
    port map (
            O => \N__38465\,
            I => \N__38447\
        );

    \I__9482\ : InMux
    port map (
            O => \N__38464\,
            I => \N__38447\
        );

    \I__9481\ : InMux
    port map (
            O => \N__38463\,
            I => \N__38434\
        );

    \I__9480\ : InMux
    port map (
            O => \N__38462\,
            I => \N__38434\
        );

    \I__9479\ : InMux
    port map (
            O => \N__38461\,
            I => \N__38434\
        );

    \I__9478\ : InMux
    port map (
            O => \N__38460\,
            I => \N__38434\
        );

    \I__9477\ : InMux
    port map (
            O => \N__38459\,
            I => \N__38434\
        );

    \I__9476\ : InMux
    port map (
            O => \N__38458\,
            I => \N__38434\
        );

    \I__9475\ : LocalMux
    port map (
            O => \N__38447\,
            I => \b2v_inst.N_645\
        );

    \I__9474\ : LocalMux
    port map (
            O => \N__38434\,
            I => \b2v_inst.N_645\
        );

    \I__9473\ : InMux
    port map (
            O => \N__38429\,
            I => \N__38426\
        );

    \I__9472\ : LocalMux
    port map (
            O => \N__38426\,
            I => \N__38423\
        );

    \I__9471\ : Span4Mux_h
    port map (
            O => \N__38423\,
            I => \N__38419\
        );

    \I__9470\ : InMux
    port map (
            O => \N__38422\,
            I => \N__38416\
        );

    \I__9469\ : Span4Mux_h
    port map (
            O => \N__38419\,
            I => \N__38413\
        );

    \I__9468\ : LocalMux
    port map (
            O => \N__38416\,
            I => \N__38409\
        );

    \I__9467\ : Span4Mux_h
    port map (
            O => \N__38413\,
            I => \N__38404\
        );

    \I__9466\ : InMux
    port map (
            O => \N__38412\,
            I => \N__38401\
        );

    \I__9465\ : Span4Mux_h
    port map (
            O => \N__38409\,
            I => \N__38398\
        );

    \I__9464\ : InMux
    port map (
            O => \N__38408\,
            I => \N__38395\
        );

    \I__9463\ : InMux
    port map (
            O => \N__38407\,
            I => \N__38392\
        );

    \I__9462\ : Odrv4
    port map (
            O => \N__38404\,
            I => \b2v_inst.dir_energiaZ0Z_6\
        );

    \I__9461\ : LocalMux
    port map (
            O => \N__38401\,
            I => \b2v_inst.dir_energiaZ0Z_6\
        );

    \I__9460\ : Odrv4
    port map (
            O => \N__38398\,
            I => \b2v_inst.dir_energiaZ0Z_6\
        );

    \I__9459\ : LocalMux
    port map (
            O => \N__38395\,
            I => \b2v_inst.dir_energiaZ0Z_6\
        );

    \I__9458\ : LocalMux
    port map (
            O => \N__38392\,
            I => \b2v_inst.dir_energiaZ0Z_6\
        );

    \I__9457\ : CascadeMux
    port map (
            O => \N__38381\,
            I => \N__38378\
        );

    \I__9456\ : InMux
    port map (
            O => \N__38378\,
            I => \N__38374\
        );

    \I__9455\ : InMux
    port map (
            O => \N__38377\,
            I => \N__38371\
        );

    \I__9454\ : LocalMux
    port map (
            O => \N__38374\,
            I => \N__38366\
        );

    \I__9453\ : LocalMux
    port map (
            O => \N__38371\,
            I => \N__38363\
        );

    \I__9452\ : InMux
    port map (
            O => \N__38370\,
            I => \N__38360\
        );

    \I__9451\ : InMux
    port map (
            O => \N__38369\,
            I => \N__38356\
        );

    \I__9450\ : Span4Mux_h
    port map (
            O => \N__38366\,
            I => \N__38352\
        );

    \I__9449\ : Span4Mux_v
    port map (
            O => \N__38363\,
            I => \N__38349\
        );

    \I__9448\ : LocalMux
    port map (
            O => \N__38360\,
            I => \N__38346\
        );

    \I__9447\ : InMux
    port map (
            O => \N__38359\,
            I => \N__38343\
        );

    \I__9446\ : LocalMux
    port map (
            O => \N__38356\,
            I => \N__38339\
        );

    \I__9445\ : InMux
    port map (
            O => \N__38355\,
            I => \N__38334\
        );

    \I__9444\ : Sp12to4
    port map (
            O => \N__38352\,
            I => \N__38331\
        );

    \I__9443\ : Span4Mux_v
    port map (
            O => \N__38349\,
            I => \N__38328\
        );

    \I__9442\ : Span4Mux_v
    port map (
            O => \N__38346\,
            I => \N__38323\
        );

    \I__9441\ : LocalMux
    port map (
            O => \N__38343\,
            I => \N__38320\
        );

    \I__9440\ : InMux
    port map (
            O => \N__38342\,
            I => \N__38317\
        );

    \I__9439\ : Sp12to4
    port map (
            O => \N__38339\,
            I => \N__38314\
        );

    \I__9438\ : InMux
    port map (
            O => \N__38338\,
            I => \N__38310\
        );

    \I__9437\ : InMux
    port map (
            O => \N__38337\,
            I => \N__38307\
        );

    \I__9436\ : LocalMux
    port map (
            O => \N__38334\,
            I => \N__38300\
        );

    \I__9435\ : Span12Mux_v
    port map (
            O => \N__38331\,
            I => \N__38300\
        );

    \I__9434\ : Sp12to4
    port map (
            O => \N__38328\,
            I => \N__38300\
        );

    \I__9433\ : InMux
    port map (
            O => \N__38327\,
            I => \N__38297\
        );

    \I__9432\ : InMux
    port map (
            O => \N__38326\,
            I => \N__38294\
        );

    \I__9431\ : Span4Mux_h
    port map (
            O => \N__38323\,
            I => \N__38289\
        );

    \I__9430\ : Span4Mux_v
    port map (
            O => \N__38320\,
            I => \N__38289\
        );

    \I__9429\ : LocalMux
    port map (
            O => \N__38317\,
            I => \N__38284\
        );

    \I__9428\ : Span12Mux_v
    port map (
            O => \N__38314\,
            I => \N__38284\
        );

    \I__9427\ : InMux
    port map (
            O => \N__38313\,
            I => \N__38281\
        );

    \I__9426\ : LocalMux
    port map (
            O => \N__38310\,
            I => \b2v_inst.indiceZ0Z_6\
        );

    \I__9425\ : LocalMux
    port map (
            O => \N__38307\,
            I => \b2v_inst.indiceZ0Z_6\
        );

    \I__9424\ : Odrv12
    port map (
            O => \N__38300\,
            I => \b2v_inst.indiceZ0Z_6\
        );

    \I__9423\ : LocalMux
    port map (
            O => \N__38297\,
            I => \b2v_inst.indiceZ0Z_6\
        );

    \I__9422\ : LocalMux
    port map (
            O => \N__38294\,
            I => \b2v_inst.indiceZ0Z_6\
        );

    \I__9421\ : Odrv4
    port map (
            O => \N__38289\,
            I => \b2v_inst.indiceZ0Z_6\
        );

    \I__9420\ : Odrv12
    port map (
            O => \N__38284\,
            I => \b2v_inst.indiceZ0Z_6\
        );

    \I__9419\ : LocalMux
    port map (
            O => \N__38281\,
            I => \b2v_inst.indiceZ0Z_6\
        );

    \I__9418\ : InMux
    port map (
            O => \N__38264\,
            I => \N__38248\
        );

    \I__9417\ : InMux
    port map (
            O => \N__38263\,
            I => \N__38248\
        );

    \I__9416\ : InMux
    port map (
            O => \N__38262\,
            I => \N__38248\
        );

    \I__9415\ : InMux
    port map (
            O => \N__38261\,
            I => \N__38248\
        );

    \I__9414\ : InMux
    port map (
            O => \N__38260\,
            I => \N__38248\
        );

    \I__9413\ : InMux
    port map (
            O => \N__38259\,
            I => \N__38239\
        );

    \I__9412\ : LocalMux
    port map (
            O => \N__38248\,
            I => \N__38236\
        );

    \I__9411\ : InMux
    port map (
            O => \N__38247\,
            I => \N__38231\
        );

    \I__9410\ : InMux
    port map (
            O => \N__38246\,
            I => \N__38231\
        );

    \I__9409\ : InMux
    port map (
            O => \N__38245\,
            I => \N__38222\
        );

    \I__9408\ : InMux
    port map (
            O => \N__38244\,
            I => \N__38222\
        );

    \I__9407\ : InMux
    port map (
            O => \N__38243\,
            I => \N__38222\
        );

    \I__9406\ : InMux
    port map (
            O => \N__38242\,
            I => \N__38222\
        );

    \I__9405\ : LocalMux
    port map (
            O => \N__38239\,
            I => \N__38219\
        );

    \I__9404\ : Span4Mux_v
    port map (
            O => \N__38236\,
            I => \N__38212\
        );

    \I__9403\ : LocalMux
    port map (
            O => \N__38231\,
            I => \N__38212\
        );

    \I__9402\ : LocalMux
    port map (
            O => \N__38222\,
            I => \N__38212\
        );

    \I__9401\ : Span4Mux_h
    port map (
            O => \N__38219\,
            I => \N__38209\
        );

    \I__9400\ : Span4Mux_h
    port map (
            O => \N__38212\,
            I => \N__38206\
        );

    \I__9399\ : Span4Mux_h
    port map (
            O => \N__38209\,
            I => \N__38203\
        );

    \I__9398\ : Odrv4
    port map (
            O => \N__38206\,
            I => \b2v_inst.N_484\
        );

    \I__9397\ : Odrv4
    port map (
            O => \N__38203\,
            I => \b2v_inst.N_484\
        );

    \I__9396\ : CascadeMux
    port map (
            O => \N__38198\,
            I => \N__38194\
        );

    \I__9395\ : CascadeMux
    port map (
            O => \N__38197\,
            I => \N__38191\
        );

    \I__9394\ : CascadeBuf
    port map (
            O => \N__38194\,
            I => \N__38188\
        );

    \I__9393\ : CascadeBuf
    port map (
            O => \N__38191\,
            I => \N__38185\
        );

    \I__9392\ : CascadeMux
    port map (
            O => \N__38188\,
            I => \N__38182\
        );

    \I__9391\ : CascadeMux
    port map (
            O => \N__38185\,
            I => \N__38179\
        );

    \I__9390\ : CascadeBuf
    port map (
            O => \N__38182\,
            I => \N__38176\
        );

    \I__9389\ : CascadeBuf
    port map (
            O => \N__38179\,
            I => \N__38173\
        );

    \I__9388\ : CascadeMux
    port map (
            O => \N__38176\,
            I => \N__38170\
        );

    \I__9387\ : CascadeMux
    port map (
            O => \N__38173\,
            I => \N__38167\
        );

    \I__9386\ : InMux
    port map (
            O => \N__38170\,
            I => \N__38164\
        );

    \I__9385\ : InMux
    port map (
            O => \N__38167\,
            I => \N__38161\
        );

    \I__9384\ : LocalMux
    port map (
            O => \N__38164\,
            I => \N_354_i\
        );

    \I__9383\ : LocalMux
    port map (
            O => \N__38161\,
            I => \N_354_i\
        );

    \I__9382\ : CascadeMux
    port map (
            O => \N__38156\,
            I => \N__38152\
        );

    \I__9381\ : InMux
    port map (
            O => \N__38155\,
            I => \N__38145\
        );

    \I__9380\ : InMux
    port map (
            O => \N__38152\,
            I => \N__38145\
        );

    \I__9379\ : InMux
    port map (
            O => \N__38151\,
            I => \N__38140\
        );

    \I__9378\ : InMux
    port map (
            O => \N__38150\,
            I => \N__38140\
        );

    \I__9377\ : LocalMux
    port map (
            O => \N__38145\,
            I => \N__38125\
        );

    \I__9376\ : LocalMux
    port map (
            O => \N__38140\,
            I => \N__38120\
        );

    \I__9375\ : SRMux
    port map (
            O => \N__38139\,
            I => \N__37847\
        );

    \I__9374\ : SRMux
    port map (
            O => \N__38138\,
            I => \N__37847\
        );

    \I__9373\ : SRMux
    port map (
            O => \N__38137\,
            I => \N__37847\
        );

    \I__9372\ : SRMux
    port map (
            O => \N__38136\,
            I => \N__37847\
        );

    \I__9371\ : SRMux
    port map (
            O => \N__38135\,
            I => \N__37847\
        );

    \I__9370\ : SRMux
    port map (
            O => \N__38134\,
            I => \N__37847\
        );

    \I__9369\ : SRMux
    port map (
            O => \N__38133\,
            I => \N__37847\
        );

    \I__9368\ : SRMux
    port map (
            O => \N__38132\,
            I => \N__37847\
        );

    \I__9367\ : SRMux
    port map (
            O => \N__38131\,
            I => \N__37847\
        );

    \I__9366\ : SRMux
    port map (
            O => \N__38130\,
            I => \N__37847\
        );

    \I__9365\ : SRMux
    port map (
            O => \N__38129\,
            I => \N__37847\
        );

    \I__9364\ : SRMux
    port map (
            O => \N__38128\,
            I => \N__37847\
        );

    \I__9363\ : Glb2LocalMux
    port map (
            O => \N__38125\,
            I => \N__37847\
        );

    \I__9362\ : SRMux
    port map (
            O => \N__38124\,
            I => \N__37847\
        );

    \I__9361\ : SRMux
    port map (
            O => \N__38123\,
            I => \N__37847\
        );

    \I__9360\ : Glb2LocalMux
    port map (
            O => \N__38120\,
            I => \N__37847\
        );

    \I__9359\ : SRMux
    port map (
            O => \N__38119\,
            I => \N__37847\
        );

    \I__9358\ : SRMux
    port map (
            O => \N__38118\,
            I => \N__37847\
        );

    \I__9357\ : SRMux
    port map (
            O => \N__38117\,
            I => \N__37847\
        );

    \I__9356\ : SRMux
    port map (
            O => \N__38116\,
            I => \N__37847\
        );

    \I__9355\ : SRMux
    port map (
            O => \N__38115\,
            I => \N__37847\
        );

    \I__9354\ : SRMux
    port map (
            O => \N__38114\,
            I => \N__37847\
        );

    \I__9353\ : SRMux
    port map (
            O => \N__38113\,
            I => \N__37847\
        );

    \I__9352\ : SRMux
    port map (
            O => \N__38112\,
            I => \N__37847\
        );

    \I__9351\ : SRMux
    port map (
            O => \N__38111\,
            I => \N__37847\
        );

    \I__9350\ : SRMux
    port map (
            O => \N__38110\,
            I => \N__37847\
        );

    \I__9349\ : SRMux
    port map (
            O => \N__38109\,
            I => \N__37847\
        );

    \I__9348\ : SRMux
    port map (
            O => \N__38108\,
            I => \N__37847\
        );

    \I__9347\ : SRMux
    port map (
            O => \N__38107\,
            I => \N__37847\
        );

    \I__9346\ : SRMux
    port map (
            O => \N__38106\,
            I => \N__37847\
        );

    \I__9345\ : SRMux
    port map (
            O => \N__38105\,
            I => \N__37847\
        );

    \I__9344\ : SRMux
    port map (
            O => \N__38104\,
            I => \N__37847\
        );

    \I__9343\ : SRMux
    port map (
            O => \N__38103\,
            I => \N__37847\
        );

    \I__9342\ : SRMux
    port map (
            O => \N__38102\,
            I => \N__37847\
        );

    \I__9341\ : SRMux
    port map (
            O => \N__38101\,
            I => \N__37847\
        );

    \I__9340\ : SRMux
    port map (
            O => \N__38100\,
            I => \N__37847\
        );

    \I__9339\ : SRMux
    port map (
            O => \N__38099\,
            I => \N__37847\
        );

    \I__9338\ : SRMux
    port map (
            O => \N__38098\,
            I => \N__37847\
        );

    \I__9337\ : SRMux
    port map (
            O => \N__38097\,
            I => \N__37847\
        );

    \I__9336\ : SRMux
    port map (
            O => \N__38096\,
            I => \N__37847\
        );

    \I__9335\ : SRMux
    port map (
            O => \N__38095\,
            I => \N__37847\
        );

    \I__9334\ : SRMux
    port map (
            O => \N__38094\,
            I => \N__37847\
        );

    \I__9333\ : SRMux
    port map (
            O => \N__38093\,
            I => \N__37847\
        );

    \I__9332\ : SRMux
    port map (
            O => \N__38092\,
            I => \N__37847\
        );

    \I__9331\ : SRMux
    port map (
            O => \N__38091\,
            I => \N__37847\
        );

    \I__9330\ : SRMux
    port map (
            O => \N__38090\,
            I => \N__37847\
        );

    \I__9329\ : SRMux
    port map (
            O => \N__38089\,
            I => \N__37847\
        );

    \I__9328\ : SRMux
    port map (
            O => \N__38088\,
            I => \N__37847\
        );

    \I__9327\ : SRMux
    port map (
            O => \N__38087\,
            I => \N__37847\
        );

    \I__9326\ : SRMux
    port map (
            O => \N__38086\,
            I => \N__37847\
        );

    \I__9325\ : SRMux
    port map (
            O => \N__38085\,
            I => \N__37847\
        );

    \I__9324\ : SRMux
    port map (
            O => \N__38084\,
            I => \N__37847\
        );

    \I__9323\ : SRMux
    port map (
            O => \N__38083\,
            I => \N__37847\
        );

    \I__9322\ : SRMux
    port map (
            O => \N__38082\,
            I => \N__37847\
        );

    \I__9321\ : SRMux
    port map (
            O => \N__38081\,
            I => \N__37847\
        );

    \I__9320\ : SRMux
    port map (
            O => \N__38080\,
            I => \N__37847\
        );

    \I__9319\ : SRMux
    port map (
            O => \N__38079\,
            I => \N__37847\
        );

    \I__9318\ : SRMux
    port map (
            O => \N__38078\,
            I => \N__37847\
        );

    \I__9317\ : SRMux
    port map (
            O => \N__38077\,
            I => \N__37847\
        );

    \I__9316\ : SRMux
    port map (
            O => \N__38076\,
            I => \N__37847\
        );

    \I__9315\ : SRMux
    port map (
            O => \N__38075\,
            I => \N__37847\
        );

    \I__9314\ : SRMux
    port map (
            O => \N__38074\,
            I => \N__37847\
        );

    \I__9313\ : SRMux
    port map (
            O => \N__38073\,
            I => \N__37847\
        );

    \I__9312\ : SRMux
    port map (
            O => \N__38072\,
            I => \N__37847\
        );

    \I__9311\ : SRMux
    port map (
            O => \N__38071\,
            I => \N__37847\
        );

    \I__9310\ : SRMux
    port map (
            O => \N__38070\,
            I => \N__37847\
        );

    \I__9309\ : SRMux
    port map (
            O => \N__38069\,
            I => \N__37847\
        );

    \I__9308\ : SRMux
    port map (
            O => \N__38068\,
            I => \N__37847\
        );

    \I__9307\ : SRMux
    port map (
            O => \N__38067\,
            I => \N__37847\
        );

    \I__9306\ : SRMux
    port map (
            O => \N__38066\,
            I => \N__37847\
        );

    \I__9305\ : SRMux
    port map (
            O => \N__38065\,
            I => \N__37847\
        );

    \I__9304\ : SRMux
    port map (
            O => \N__38064\,
            I => \N__37847\
        );

    \I__9303\ : SRMux
    port map (
            O => \N__38063\,
            I => \N__37847\
        );

    \I__9302\ : SRMux
    port map (
            O => \N__38062\,
            I => \N__37847\
        );

    \I__9301\ : SRMux
    port map (
            O => \N__38061\,
            I => \N__37847\
        );

    \I__9300\ : SRMux
    port map (
            O => \N__38060\,
            I => \N__37847\
        );

    \I__9299\ : SRMux
    port map (
            O => \N__38059\,
            I => \N__37847\
        );

    \I__9298\ : SRMux
    port map (
            O => \N__38058\,
            I => \N__37847\
        );

    \I__9297\ : SRMux
    port map (
            O => \N__38057\,
            I => \N__37847\
        );

    \I__9296\ : SRMux
    port map (
            O => \N__38056\,
            I => \N__37847\
        );

    \I__9295\ : SRMux
    port map (
            O => \N__38055\,
            I => \N__37847\
        );

    \I__9294\ : SRMux
    port map (
            O => \N__38054\,
            I => \N__37847\
        );

    \I__9293\ : SRMux
    port map (
            O => \N__38053\,
            I => \N__37847\
        );

    \I__9292\ : SRMux
    port map (
            O => \N__38052\,
            I => \N__37847\
        );

    \I__9291\ : SRMux
    port map (
            O => \N__38051\,
            I => \N__37847\
        );

    \I__9290\ : SRMux
    port map (
            O => \N__38050\,
            I => \N__37847\
        );

    \I__9289\ : SRMux
    port map (
            O => \N__38049\,
            I => \N__37847\
        );

    \I__9288\ : SRMux
    port map (
            O => \N__38048\,
            I => \N__37847\
        );

    \I__9287\ : SRMux
    port map (
            O => \N__38047\,
            I => \N__37847\
        );

    \I__9286\ : SRMux
    port map (
            O => \N__38046\,
            I => \N__37847\
        );

    \I__9285\ : SRMux
    port map (
            O => \N__38045\,
            I => \N__37847\
        );

    \I__9284\ : SRMux
    port map (
            O => \N__38044\,
            I => \N__37847\
        );

    \I__9283\ : SRMux
    port map (
            O => \N__38043\,
            I => \N__37847\
        );

    \I__9282\ : SRMux
    port map (
            O => \N__38042\,
            I => \N__37847\
        );

    \I__9281\ : SRMux
    port map (
            O => \N__38041\,
            I => \N__37847\
        );

    \I__9280\ : SRMux
    port map (
            O => \N__38040\,
            I => \N__37847\
        );

    \I__9279\ : GlobalMux
    port map (
            O => \N__37847\,
            I => \N__37844\
        );

    \I__9278\ : gio2CtrlBuf
    port map (
            O => \N__37844\,
            I => reset_c_i_g
        );

    \I__9277\ : InMux
    port map (
            O => \N__37841\,
            I => \N__37837\
        );

    \I__9276\ : CascadeMux
    port map (
            O => \N__37840\,
            I => \N__37832\
        );

    \I__9275\ : LocalMux
    port map (
            O => \N__37837\,
            I => \N__37827\
        );

    \I__9274\ : InMux
    port map (
            O => \N__37836\,
            I => \N__37824\
        );

    \I__9273\ : CascadeMux
    port map (
            O => \N__37835\,
            I => \N__37820\
        );

    \I__9272\ : InMux
    port map (
            O => \N__37832\,
            I => \N__37814\
        );

    \I__9271\ : InMux
    port map (
            O => \N__37831\,
            I => \N__37814\
        );

    \I__9270\ : CascadeMux
    port map (
            O => \N__37830\,
            I => \N__37810\
        );

    \I__9269\ : Span4Mux_v
    port map (
            O => \N__37827\,
            I => \N__37802\
        );

    \I__9268\ : LocalMux
    port map (
            O => \N__37824\,
            I => \N__37802\
        );

    \I__9267\ : InMux
    port map (
            O => \N__37823\,
            I => \N__37799\
        );

    \I__9266\ : InMux
    port map (
            O => \N__37820\,
            I => \N__37794\
        );

    \I__9265\ : InMux
    port map (
            O => \N__37819\,
            I => \N__37794\
        );

    \I__9264\ : LocalMux
    port map (
            O => \N__37814\,
            I => \N__37786\
        );

    \I__9263\ : InMux
    port map (
            O => \N__37813\,
            I => \N__37783\
        );

    \I__9262\ : InMux
    port map (
            O => \N__37810\,
            I => \N__37778\
        );

    \I__9261\ : InMux
    port map (
            O => \N__37809\,
            I => \N__37778\
        );

    \I__9260\ : InMux
    port map (
            O => \N__37808\,
            I => \N__37773\
        );

    \I__9259\ : InMux
    port map (
            O => \N__37807\,
            I => \N__37773\
        );

    \I__9258\ : Span4Mux_v
    port map (
            O => \N__37802\,
            I => \N__37766\
        );

    \I__9257\ : LocalMux
    port map (
            O => \N__37799\,
            I => \N__37766\
        );

    \I__9256\ : LocalMux
    port map (
            O => \N__37794\,
            I => \N__37766\
        );

    \I__9255\ : InMux
    port map (
            O => \N__37793\,
            I => \N__37763\
        );

    \I__9254\ : InMux
    port map (
            O => \N__37792\,
            I => \N__37760\
        );

    \I__9253\ : InMux
    port map (
            O => \N__37791\,
            I => \N__37754\
        );

    \I__9252\ : InMux
    port map (
            O => \N__37790\,
            I => \N__37754\
        );

    \I__9251\ : InMux
    port map (
            O => \N__37789\,
            I => \N__37750\
        );

    \I__9250\ : Span4Mux_h
    port map (
            O => \N__37786\,
            I => \N__37741\
        );

    \I__9249\ : LocalMux
    port map (
            O => \N__37783\,
            I => \N__37741\
        );

    \I__9248\ : LocalMux
    port map (
            O => \N__37778\,
            I => \N__37741\
        );

    \I__9247\ : LocalMux
    port map (
            O => \N__37773\,
            I => \N__37741\
        );

    \I__9246\ : Span4Mux_v
    port map (
            O => \N__37766\,
            I => \N__37734\
        );

    \I__9245\ : LocalMux
    port map (
            O => \N__37763\,
            I => \N__37734\
        );

    \I__9244\ : LocalMux
    port map (
            O => \N__37760\,
            I => \N__37734\
        );

    \I__9243\ : CascadeMux
    port map (
            O => \N__37759\,
            I => \N__37729\
        );

    \I__9242\ : LocalMux
    port map (
            O => \N__37754\,
            I => \N__37725\
        );

    \I__9241\ : InMux
    port map (
            O => \N__37753\,
            I => \N__37722\
        );

    \I__9240\ : LocalMux
    port map (
            O => \N__37750\,
            I => \N__37719\
        );

    \I__9239\ : Span4Mux_v
    port map (
            O => \N__37741\,
            I => \N__37716\
        );

    \I__9238\ : Span4Mux_v
    port map (
            O => \N__37734\,
            I => \N__37713\
        );

    \I__9237\ : InMux
    port map (
            O => \N__37733\,
            I => \N__37710\
        );

    \I__9236\ : InMux
    port map (
            O => \N__37732\,
            I => \N__37706\
        );

    \I__9235\ : InMux
    port map (
            O => \N__37729\,
            I => \N__37701\
        );

    \I__9234\ : InMux
    port map (
            O => \N__37728\,
            I => \N__37701\
        );

    \I__9233\ : Span4Mux_v
    port map (
            O => \N__37725\,
            I => \N__37698\
        );

    \I__9232\ : LocalMux
    port map (
            O => \N__37722\,
            I => \N__37695\
        );

    \I__9231\ : Span4Mux_v
    port map (
            O => \N__37719\,
            I => \N__37692\
        );

    \I__9230\ : Span4Mux_h
    port map (
            O => \N__37716\,
            I => \N__37685\
        );

    \I__9229\ : Span4Mux_h
    port map (
            O => \N__37713\,
            I => \N__37685\
        );

    \I__9228\ : LocalMux
    port map (
            O => \N__37710\,
            I => \N__37685\
        );

    \I__9227\ : CascadeMux
    port map (
            O => \N__37709\,
            I => \N__37682\
        );

    \I__9226\ : LocalMux
    port map (
            O => \N__37706\,
            I => \N__37673\
        );

    \I__9225\ : LocalMux
    port map (
            O => \N__37701\,
            I => \N__37673\
        );

    \I__9224\ : Span4Mux_h
    port map (
            O => \N__37698\,
            I => \N__37664\
        );

    \I__9223\ : Span4Mux_v
    port map (
            O => \N__37695\,
            I => \N__37664\
        );

    \I__9222\ : Span4Mux_h
    port map (
            O => \N__37692\,
            I => \N__37664\
        );

    \I__9221\ : Span4Mux_h
    port map (
            O => \N__37685\,
            I => \N__37664\
        );

    \I__9220\ : InMux
    port map (
            O => \N__37682\,
            I => \N__37661\
        );

    \I__9219\ : InMux
    port map (
            O => \N__37681\,
            I => \N__37658\
        );

    \I__9218\ : InMux
    port map (
            O => \N__37680\,
            I => \N__37653\
        );

    \I__9217\ : InMux
    port map (
            O => \N__37679\,
            I => \N__37653\
        );

    \I__9216\ : InMux
    port map (
            O => \N__37678\,
            I => \N__37650\
        );

    \I__9215\ : Odrv12
    port map (
            O => \N__37673\,
            I => \b2v_inst.N_828\
        );

    \I__9214\ : Odrv4
    port map (
            O => \N__37664\,
            I => \b2v_inst.N_828\
        );

    \I__9213\ : LocalMux
    port map (
            O => \N__37661\,
            I => \b2v_inst.N_828\
        );

    \I__9212\ : LocalMux
    port map (
            O => \N__37658\,
            I => \b2v_inst.N_828\
        );

    \I__9211\ : LocalMux
    port map (
            O => \N__37653\,
            I => \b2v_inst.N_828\
        );

    \I__9210\ : LocalMux
    port map (
            O => \N__37650\,
            I => \b2v_inst.N_828\
        );

    \I__9209\ : InMux
    port map (
            O => \N__37637\,
            I => \N__37634\
        );

    \I__9208\ : LocalMux
    port map (
            O => \N__37634\,
            I => \b2v_inst.un16_data_ram_cantidad_o_cry_4_c_RNIDGFOZ0\
        );

    \I__9207\ : CascadeMux
    port map (
            O => \N__37631\,
            I => \N__37628\
        );

    \I__9206\ : InMux
    port map (
            O => \N__37628\,
            I => \N__37623\
        );

    \I__9205\ : CascadeMux
    port map (
            O => \N__37627\,
            I => \N__37620\
        );

    \I__9204\ : CascadeMux
    port map (
            O => \N__37626\,
            I => \N__37617\
        );

    \I__9203\ : LocalMux
    port map (
            O => \N__37623\,
            I => \N__37614\
        );

    \I__9202\ : InMux
    port map (
            O => \N__37620\,
            I => \N__37611\
        );

    \I__9201\ : InMux
    port map (
            O => \N__37617\,
            I => \N__37608\
        );

    \I__9200\ : Span4Mux_v
    port map (
            O => \N__37614\,
            I => \N__37605\
        );

    \I__9199\ : LocalMux
    port map (
            O => \N__37611\,
            I => \N__37602\
        );

    \I__9198\ : LocalMux
    port map (
            O => \N__37608\,
            I => \N__37599\
        );

    \I__9197\ : Span4Mux_h
    port map (
            O => \N__37605\,
            I => \N__37594\
        );

    \I__9196\ : Span4Mux_h
    port map (
            O => \N__37602\,
            I => \N__37591\
        );

    \I__9195\ : Span4Mux_v
    port map (
            O => \N__37599\,
            I => \N__37588\
        );

    \I__9194\ : InMux
    port map (
            O => \N__37598\,
            I => \N__37585\
        );

    \I__9193\ : InMux
    port map (
            O => \N__37597\,
            I => \N__37582\
        );

    \I__9192\ : Span4Mux_h
    port map (
            O => \N__37594\,
            I => \N__37573\
        );

    \I__9191\ : Span4Mux_v
    port map (
            O => \N__37591\,
            I => \N__37573\
        );

    \I__9190\ : Span4Mux_h
    port map (
            O => \N__37588\,
            I => \N__37573\
        );

    \I__9189\ : LocalMux
    port map (
            O => \N__37585\,
            I => \N__37573\
        );

    \I__9188\ : LocalMux
    port map (
            O => \N__37582\,
            I => \N__37570\
        );

    \I__9187\ : Span4Mux_h
    port map (
            O => \N__37573\,
            I => \N__37567\
        );

    \I__9186\ : Odrv12
    port map (
            O => \N__37570\,
            I => b2v_inst_data_a_escribir_5
        );

    \I__9185\ : Odrv4
    port map (
            O => \N__37567\,
            I => b2v_inst_data_a_escribir_5
        );

    \I__9184\ : InMux
    port map (
            O => \N__37562\,
            I => \N__37557\
        );

    \I__9183\ : InMux
    port map (
            O => \N__37561\,
            I => \N__37554\
        );

    \I__9182\ : CascadeMux
    port map (
            O => \N__37560\,
            I => \N__37551\
        );

    \I__9181\ : LocalMux
    port map (
            O => \N__37557\,
            I => \N__37540\
        );

    \I__9180\ : LocalMux
    port map (
            O => \N__37554\,
            I => \N__37537\
        );

    \I__9179\ : InMux
    port map (
            O => \N__37551\,
            I => \N__37532\
        );

    \I__9178\ : InMux
    port map (
            O => \N__37550\,
            I => \N__37532\
        );

    \I__9177\ : InMux
    port map (
            O => \N__37549\,
            I => \N__37527\
        );

    \I__9176\ : InMux
    port map (
            O => \N__37548\,
            I => \N__37524\
        );

    \I__9175\ : InMux
    port map (
            O => \N__37547\,
            I => \N__37521\
        );

    \I__9174\ : InMux
    port map (
            O => \N__37546\,
            I => \N__37516\
        );

    \I__9173\ : InMux
    port map (
            O => \N__37545\,
            I => \N__37516\
        );

    \I__9172\ : InMux
    port map (
            O => \N__37544\,
            I => \N__37511\
        );

    \I__9171\ : InMux
    port map (
            O => \N__37543\,
            I => \N__37511\
        );

    \I__9170\ : Span4Mux_v
    port map (
            O => \N__37540\,
            I => \N__37504\
        );

    \I__9169\ : Span4Mux_h
    port map (
            O => \N__37537\,
            I => \N__37504\
        );

    \I__9168\ : LocalMux
    port map (
            O => \N__37532\,
            I => \N__37499\
        );

    \I__9167\ : InMux
    port map (
            O => \N__37531\,
            I => \N__37491\
        );

    \I__9166\ : InMux
    port map (
            O => \N__37530\,
            I => \N__37491\
        );

    \I__9165\ : LocalMux
    port map (
            O => \N__37527\,
            I => \N__37480\
        );

    \I__9164\ : LocalMux
    port map (
            O => \N__37524\,
            I => \N__37480\
        );

    \I__9163\ : LocalMux
    port map (
            O => \N__37521\,
            I => \N__37480\
        );

    \I__9162\ : LocalMux
    port map (
            O => \N__37516\,
            I => \N__37480\
        );

    \I__9161\ : LocalMux
    port map (
            O => \N__37511\,
            I => \N__37480\
        );

    \I__9160\ : InMux
    port map (
            O => \N__37510\,
            I => \N__37474\
        );

    \I__9159\ : InMux
    port map (
            O => \N__37509\,
            I => \N__37474\
        );

    \I__9158\ : Span4Mux_h
    port map (
            O => \N__37504\,
            I => \N__37471\
        );

    \I__9157\ : InMux
    port map (
            O => \N__37503\,
            I => \N__37468\
        );

    \I__9156\ : InMux
    port map (
            O => \N__37502\,
            I => \N__37462\
        );

    \I__9155\ : Span4Mux_h
    port map (
            O => \N__37499\,
            I => \N__37456\
        );

    \I__9154\ : InMux
    port map (
            O => \N__37498\,
            I => \N__37453\
        );

    \I__9153\ : InMux
    port map (
            O => \N__37497\,
            I => \N__37450\
        );

    \I__9152\ : InMux
    port map (
            O => \N__37496\,
            I => \N__37446\
        );

    \I__9151\ : LocalMux
    port map (
            O => \N__37491\,
            I => \N__37441\
        );

    \I__9150\ : Span4Mux_v
    port map (
            O => \N__37480\,
            I => \N__37441\
        );

    \I__9149\ : InMux
    port map (
            O => \N__37479\,
            I => \N__37438\
        );

    \I__9148\ : LocalMux
    port map (
            O => \N__37474\,
            I => \N__37431\
        );

    \I__9147\ : Span4Mux_h
    port map (
            O => \N__37471\,
            I => \N__37431\
        );

    \I__9146\ : LocalMux
    port map (
            O => \N__37468\,
            I => \N__37431\
        );

    \I__9145\ : InMux
    port map (
            O => \N__37467\,
            I => \N__37426\
        );

    \I__9144\ : InMux
    port map (
            O => \N__37466\,
            I => \N__37426\
        );

    \I__9143\ : InMux
    port map (
            O => \N__37465\,
            I => \N__37423\
        );

    \I__9142\ : LocalMux
    port map (
            O => \N__37462\,
            I => \N__37420\
        );

    \I__9141\ : InMux
    port map (
            O => \N__37461\,
            I => \N__37415\
        );

    \I__9140\ : InMux
    port map (
            O => \N__37460\,
            I => \N__37415\
        );

    \I__9139\ : InMux
    port map (
            O => \N__37459\,
            I => \N__37412\
        );

    \I__9138\ : Span4Mux_v
    port map (
            O => \N__37456\,
            I => \N__37407\
        );

    \I__9137\ : LocalMux
    port map (
            O => \N__37453\,
            I => \N__37407\
        );

    \I__9136\ : LocalMux
    port map (
            O => \N__37450\,
            I => \N__37401\
        );

    \I__9135\ : InMux
    port map (
            O => \N__37449\,
            I => \N__37398\
        );

    \I__9134\ : LocalMux
    port map (
            O => \N__37446\,
            I => \N__37393\
        );

    \I__9133\ : Span4Mux_h
    port map (
            O => \N__37441\,
            I => \N__37390\
        );

    \I__9132\ : LocalMux
    port map (
            O => \N__37438\,
            I => \N__37385\
        );

    \I__9131\ : Span4Mux_v
    port map (
            O => \N__37431\,
            I => \N__37385\
        );

    \I__9130\ : LocalMux
    port map (
            O => \N__37426\,
            I => \N__37381\
        );

    \I__9129\ : LocalMux
    port map (
            O => \N__37423\,
            I => \N__37370\
        );

    \I__9128\ : Span4Mux_v
    port map (
            O => \N__37420\,
            I => \N__37370\
        );

    \I__9127\ : LocalMux
    port map (
            O => \N__37415\,
            I => \N__37370\
        );

    \I__9126\ : LocalMux
    port map (
            O => \N__37412\,
            I => \N__37370\
        );

    \I__9125\ : Span4Mux_h
    port map (
            O => \N__37407\,
            I => \N__37370\
        );

    \I__9124\ : InMux
    port map (
            O => \N__37406\,
            I => \N__37365\
        );

    \I__9123\ : InMux
    port map (
            O => \N__37405\,
            I => \N__37365\
        );

    \I__9122\ : InMux
    port map (
            O => \N__37404\,
            I => \N__37362\
        );

    \I__9121\ : Span12Mux_h
    port map (
            O => \N__37401\,
            I => \N__37359\
        );

    \I__9120\ : LocalMux
    port map (
            O => \N__37398\,
            I => \N__37356\
        );

    \I__9119\ : InMux
    port map (
            O => \N__37397\,
            I => \N__37351\
        );

    \I__9118\ : InMux
    port map (
            O => \N__37396\,
            I => \N__37351\
        );

    \I__9117\ : Span4Mux_h
    port map (
            O => \N__37393\,
            I => \N__37348\
        );

    \I__9116\ : Span4Mux_h
    port map (
            O => \N__37390\,
            I => \N__37343\
        );

    \I__9115\ : Span4Mux_v
    port map (
            O => \N__37385\,
            I => \N__37343\
        );

    \I__9114\ : InMux
    port map (
            O => \N__37384\,
            I => \N__37340\
        );

    \I__9113\ : Span4Mux_h
    port map (
            O => \N__37381\,
            I => \N__37335\
        );

    \I__9112\ : Span4Mux_h
    port map (
            O => \N__37370\,
            I => \N__37335\
        );

    \I__9111\ : LocalMux
    port map (
            O => \N__37365\,
            I => \b2v_inst.N_514\
        );

    \I__9110\ : LocalMux
    port map (
            O => \N__37362\,
            I => \b2v_inst.N_514\
        );

    \I__9109\ : Odrv12
    port map (
            O => \N__37359\,
            I => \b2v_inst.N_514\
        );

    \I__9108\ : Odrv4
    port map (
            O => \N__37356\,
            I => \b2v_inst.N_514\
        );

    \I__9107\ : LocalMux
    port map (
            O => \N__37351\,
            I => \b2v_inst.N_514\
        );

    \I__9106\ : Odrv4
    port map (
            O => \N__37348\,
            I => \b2v_inst.N_514\
        );

    \I__9105\ : Odrv4
    port map (
            O => \N__37343\,
            I => \b2v_inst.N_514\
        );

    \I__9104\ : LocalMux
    port map (
            O => \N__37340\,
            I => \b2v_inst.N_514\
        );

    \I__9103\ : Odrv4
    port map (
            O => \N__37335\,
            I => \b2v_inst.N_514\
        );

    \I__9102\ : InMux
    port map (
            O => \N__37316\,
            I => \N__37313\
        );

    \I__9101\ : LocalMux
    port map (
            O => \N__37313\,
            I => \N__37310\
        );

    \I__9100\ : Odrv4
    port map (
            O => \N__37310\,
            I => \N_547_i\
        );

    \I__9099\ : CascadeMux
    port map (
            O => \N__37307\,
            I => \N__37304\
        );

    \I__9098\ : InMux
    port map (
            O => \N__37304\,
            I => \N__37293\
        );

    \I__9097\ : CascadeMux
    port map (
            O => \N__37303\,
            I => \N__37289\
        );

    \I__9096\ : InMux
    port map (
            O => \N__37302\,
            I => \N__37273\
        );

    \I__9095\ : InMux
    port map (
            O => \N__37301\,
            I => \N__37273\
        );

    \I__9094\ : InMux
    port map (
            O => \N__37300\,
            I => \N__37273\
        );

    \I__9093\ : InMux
    port map (
            O => \N__37299\,
            I => \N__37273\
        );

    \I__9092\ : InMux
    port map (
            O => \N__37298\,
            I => \N__37266\
        );

    \I__9091\ : InMux
    port map (
            O => \N__37297\,
            I => \N__37266\
        );

    \I__9090\ : InMux
    port map (
            O => \N__37296\,
            I => \N__37266\
        );

    \I__9089\ : LocalMux
    port map (
            O => \N__37293\,
            I => \N__37260\
        );

    \I__9088\ : SRMux
    port map (
            O => \N__37292\,
            I => \N__37257\
        );

    \I__9087\ : InMux
    port map (
            O => \N__37289\,
            I => \N__37253\
        );

    \I__9086\ : CascadeMux
    port map (
            O => \N__37288\,
            I => \N__37250\
        );

    \I__9085\ : SRMux
    port map (
            O => \N__37287\,
            I => \N__37246\
        );

    \I__9084\ : SRMux
    port map (
            O => \N__37286\,
            I => \N__37243\
        );

    \I__9083\ : SRMux
    port map (
            O => \N__37285\,
            I => \N__37239\
        );

    \I__9082\ : SRMux
    port map (
            O => \N__37284\,
            I => \N__37236\
        );

    \I__9081\ : SRMux
    port map (
            O => \N__37283\,
            I => \N__37232\
        );

    \I__9080\ : SRMux
    port map (
            O => \N__37282\,
            I => \N__37228\
        );

    \I__9079\ : LocalMux
    port map (
            O => \N__37273\,
            I => \N__37221\
        );

    \I__9078\ : LocalMux
    port map (
            O => \N__37266\,
            I => \N__37221\
        );

    \I__9077\ : InMux
    port map (
            O => \N__37265\,
            I => \N__37218\
        );

    \I__9076\ : InMux
    port map (
            O => \N__37264\,
            I => \N__37214\
        );

    \I__9075\ : InMux
    port map (
            O => \N__37263\,
            I => \N__37209\
        );

    \I__9074\ : Span4Mux_v
    port map (
            O => \N__37260\,
            I => \N__37206\
        );

    \I__9073\ : LocalMux
    port map (
            O => \N__37257\,
            I => \N__37203\
        );

    \I__9072\ : SRMux
    port map (
            O => \N__37256\,
            I => \N__37200\
        );

    \I__9071\ : LocalMux
    port map (
            O => \N__37253\,
            I => \N__37195\
        );

    \I__9070\ : InMux
    port map (
            O => \N__37250\,
            I => \N__37192\
        );

    \I__9069\ : SRMux
    port map (
            O => \N__37249\,
            I => \N__37189\
        );

    \I__9068\ : LocalMux
    port map (
            O => \N__37246\,
            I => \N__37184\
        );

    \I__9067\ : LocalMux
    port map (
            O => \N__37243\,
            I => \N__37184\
        );

    \I__9066\ : SRMux
    port map (
            O => \N__37242\,
            I => \N__37181\
        );

    \I__9065\ : LocalMux
    port map (
            O => \N__37239\,
            I => \N__37176\
        );

    \I__9064\ : LocalMux
    port map (
            O => \N__37236\,
            I => \N__37176\
        );

    \I__9063\ : SRMux
    port map (
            O => \N__37235\,
            I => \N__37173\
        );

    \I__9062\ : LocalMux
    port map (
            O => \N__37232\,
            I => \N__37170\
        );

    \I__9061\ : SRMux
    port map (
            O => \N__37231\,
            I => \N__37167\
        );

    \I__9060\ : LocalMux
    port map (
            O => \N__37228\,
            I => \N__37164\
        );

    \I__9059\ : SRMux
    port map (
            O => \N__37227\,
            I => \N__37161\
        );

    \I__9058\ : SRMux
    port map (
            O => \N__37226\,
            I => \N__37148\
        );

    \I__9057\ : Span4Mux_h
    port map (
            O => \N__37221\,
            I => \N__37143\
        );

    \I__9056\ : LocalMux
    port map (
            O => \N__37218\,
            I => \N__37143\
        );

    \I__9055\ : InMux
    port map (
            O => \N__37217\,
            I => \N__37140\
        );

    \I__9054\ : LocalMux
    port map (
            O => \N__37214\,
            I => \N__37137\
        );

    \I__9053\ : SRMux
    port map (
            O => \N__37213\,
            I => \N__37134\
        );

    \I__9052\ : SRMux
    port map (
            O => \N__37212\,
            I => \N__37130\
        );

    \I__9051\ : LocalMux
    port map (
            O => \N__37209\,
            I => \N__37126\
        );

    \I__9050\ : Span4Mux_h
    port map (
            O => \N__37206\,
            I => \N__37119\
        );

    \I__9049\ : Span4Mux_v
    port map (
            O => \N__37203\,
            I => \N__37119\
        );

    \I__9048\ : LocalMux
    port map (
            O => \N__37200\,
            I => \N__37119\
        );

    \I__9047\ : SRMux
    port map (
            O => \N__37199\,
            I => \N__37116\
        );

    \I__9046\ : SRMux
    port map (
            O => \N__37198\,
            I => \N__37113\
        );

    \I__9045\ : Span4Mux_h
    port map (
            O => \N__37195\,
            I => \N__37107\
        );

    \I__9044\ : LocalMux
    port map (
            O => \N__37192\,
            I => \N__37107\
        );

    \I__9043\ : LocalMux
    port map (
            O => \N__37189\,
            I => \N__37100\
        );

    \I__9042\ : Span4Mux_v
    port map (
            O => \N__37184\,
            I => \N__37100\
        );

    \I__9041\ : LocalMux
    port map (
            O => \N__37181\,
            I => \N__37100\
        );

    \I__9040\ : Span4Mux_v
    port map (
            O => \N__37176\,
            I => \N__37095\
        );

    \I__9039\ : LocalMux
    port map (
            O => \N__37173\,
            I => \N__37095\
        );

    \I__9038\ : Span4Mux_v
    port map (
            O => \N__37170\,
            I => \N__37090\
        );

    \I__9037\ : LocalMux
    port map (
            O => \N__37167\,
            I => \N__37090\
        );

    \I__9036\ : Span4Mux_v
    port map (
            O => \N__37164\,
            I => \N__37085\
        );

    \I__9035\ : LocalMux
    port map (
            O => \N__37161\,
            I => \N__37085\
        );

    \I__9034\ : SRMux
    port map (
            O => \N__37160\,
            I => \N__37082\
        );

    \I__9033\ : CascadeMux
    port map (
            O => \N__37159\,
            I => \N__37079\
        );

    \I__9032\ : CascadeMux
    port map (
            O => \N__37158\,
            I => \N__37076\
        );

    \I__9031\ : CascadeMux
    port map (
            O => \N__37157\,
            I => \N__37073\
        );

    \I__9030\ : CascadeMux
    port map (
            O => \N__37156\,
            I => \N__37070\
        );

    \I__9029\ : CascadeMux
    port map (
            O => \N__37155\,
            I => \N__37067\
        );

    \I__9028\ : CascadeMux
    port map (
            O => \N__37154\,
            I => \N__37064\
        );

    \I__9027\ : CascadeMux
    port map (
            O => \N__37153\,
            I => \N__37060\
        );

    \I__9026\ : CascadeMux
    port map (
            O => \N__37152\,
            I => \N__37057\
        );

    \I__9025\ : CascadeMux
    port map (
            O => \N__37151\,
            I => \N__37053\
        );

    \I__9024\ : LocalMux
    port map (
            O => \N__37148\,
            I => \N__37050\
        );

    \I__9023\ : Span4Mux_v
    port map (
            O => \N__37143\,
            I => \N__37047\
        );

    \I__9022\ : LocalMux
    port map (
            O => \N__37140\,
            I => \N__37044\
        );

    \I__9021\ : Span4Mux_v
    port map (
            O => \N__37137\,
            I => \N__37039\
        );

    \I__9020\ : LocalMux
    port map (
            O => \N__37134\,
            I => \N__37039\
        );

    \I__9019\ : CascadeMux
    port map (
            O => \N__37133\,
            I => \N__37036\
        );

    \I__9018\ : LocalMux
    port map (
            O => \N__37130\,
            I => \N__37033\
        );

    \I__9017\ : SRMux
    port map (
            O => \N__37129\,
            I => \N__37030\
        );

    \I__9016\ : Span4Mux_v
    port map (
            O => \N__37126\,
            I => \N__37026\
        );

    \I__9015\ : Span4Mux_h
    port map (
            O => \N__37119\,
            I => \N__37019\
        );

    \I__9014\ : LocalMux
    port map (
            O => \N__37116\,
            I => \N__37019\
        );

    \I__9013\ : LocalMux
    port map (
            O => \N__37113\,
            I => \N__37019\
        );

    \I__9012\ : SRMux
    port map (
            O => \N__37112\,
            I => \N__37016\
        );

    \I__9011\ : Span4Mux_v
    port map (
            O => \N__37107\,
            I => \N__37009\
        );

    \I__9010\ : Span4Mux_v
    port map (
            O => \N__37100\,
            I => \N__37004\
        );

    \I__9009\ : Span4Mux_v
    port map (
            O => \N__37095\,
            I => \N__37004\
        );

    \I__9008\ : Span4Mux_v
    port map (
            O => \N__37090\,
            I => \N__36997\
        );

    \I__9007\ : Span4Mux_v
    port map (
            O => \N__37085\,
            I => \N__36997\
        );

    \I__9006\ : LocalMux
    port map (
            O => \N__37082\,
            I => \N__36997\
        );

    \I__9005\ : InMux
    port map (
            O => \N__37079\,
            I => \N__36991\
        );

    \I__9004\ : InMux
    port map (
            O => \N__37076\,
            I => \N__36991\
        );

    \I__9003\ : InMux
    port map (
            O => \N__37073\,
            I => \N__36984\
        );

    \I__9002\ : InMux
    port map (
            O => \N__37070\,
            I => \N__36984\
        );

    \I__9001\ : InMux
    port map (
            O => \N__37067\,
            I => \N__36984\
        );

    \I__9000\ : InMux
    port map (
            O => \N__37064\,
            I => \N__36975\
        );

    \I__8999\ : InMux
    port map (
            O => \N__37063\,
            I => \N__36975\
        );

    \I__8998\ : InMux
    port map (
            O => \N__37060\,
            I => \N__36975\
        );

    \I__8997\ : InMux
    port map (
            O => \N__37057\,
            I => \N__36975\
        );

    \I__8996\ : InMux
    port map (
            O => \N__37056\,
            I => \N__36970\
        );

    \I__8995\ : InMux
    port map (
            O => \N__37053\,
            I => \N__36970\
        );

    \I__8994\ : Span4Mux_h
    port map (
            O => \N__37050\,
            I => \N__36967\
        );

    \I__8993\ : Span4Mux_h
    port map (
            O => \N__37047\,
            I => \N__36960\
        );

    \I__8992\ : Span4Mux_v
    port map (
            O => \N__37044\,
            I => \N__36960\
        );

    \I__8991\ : Span4Mux_h
    port map (
            O => \N__37039\,
            I => \N__36960\
        );

    \I__8990\ : InMux
    port map (
            O => \N__37036\,
            I => \N__36957\
        );

    \I__8989\ : Span4Mux_v
    port map (
            O => \N__37033\,
            I => \N__36952\
        );

    \I__8988\ : LocalMux
    port map (
            O => \N__37030\,
            I => \N__36952\
        );

    \I__8987\ : SRMux
    port map (
            O => \N__37029\,
            I => \N__36949\
        );

    \I__8986\ : Span4Mux_h
    port map (
            O => \N__37026\,
            I => \N__36942\
        );

    \I__8985\ : Span4Mux_v
    port map (
            O => \N__37019\,
            I => \N__36942\
        );

    \I__8984\ : LocalMux
    port map (
            O => \N__37016\,
            I => \N__36942\
        );

    \I__8983\ : SRMux
    port map (
            O => \N__37015\,
            I => \N__36939\
        );

    \I__8982\ : SRMux
    port map (
            O => \N__37014\,
            I => \N__36935\
        );

    \I__8981\ : SRMux
    port map (
            O => \N__37013\,
            I => \N__36932\
        );

    \I__8980\ : SRMux
    port map (
            O => \N__37012\,
            I => \N__36929\
        );

    \I__8979\ : Span4Mux_v
    port map (
            O => \N__37009\,
            I => \N__36922\
        );

    \I__8978\ : Span4Mux_h
    port map (
            O => \N__37004\,
            I => \N__36922\
        );

    \I__8977\ : Span4Mux_h
    port map (
            O => \N__36997\,
            I => \N__36922\
        );

    \I__8976\ : SRMux
    port map (
            O => \N__36996\,
            I => \N__36918\
        );

    \I__8975\ : LocalMux
    port map (
            O => \N__36991\,
            I => \N__36915\
        );

    \I__8974\ : LocalMux
    port map (
            O => \N__36984\,
            I => \N__36908\
        );

    \I__8973\ : LocalMux
    port map (
            O => \N__36975\,
            I => \N__36908\
        );

    \I__8972\ : LocalMux
    port map (
            O => \N__36970\,
            I => \N__36908\
        );

    \I__8971\ : Span4Mux_h
    port map (
            O => \N__36967\,
            I => \N__36905\
        );

    \I__8970\ : Span4Mux_h
    port map (
            O => \N__36960\,
            I => \N__36900\
        );

    \I__8969\ : LocalMux
    port map (
            O => \N__36957\,
            I => \N__36900\
        );

    \I__8968\ : Span4Mux_v
    port map (
            O => \N__36952\,
            I => \N__36891\
        );

    \I__8967\ : LocalMux
    port map (
            O => \N__36949\,
            I => \N__36891\
        );

    \I__8966\ : Span4Mux_h
    port map (
            O => \N__36942\,
            I => \N__36891\
        );

    \I__8965\ : LocalMux
    port map (
            O => \N__36939\,
            I => \N__36891\
        );

    \I__8964\ : SRMux
    port map (
            O => \N__36938\,
            I => \N__36888\
        );

    \I__8963\ : LocalMux
    port map (
            O => \N__36935\,
            I => \N__36883\
        );

    \I__8962\ : LocalMux
    port map (
            O => \N__36932\,
            I => \N__36883\
        );

    \I__8961\ : LocalMux
    port map (
            O => \N__36929\,
            I => \N__36880\
        );

    \I__8960\ : Span4Mux_h
    port map (
            O => \N__36922\,
            I => \N__36877\
        );

    \I__8959\ : SRMux
    port map (
            O => \N__36921\,
            I => \N__36874\
        );

    \I__8958\ : LocalMux
    port map (
            O => \N__36918\,
            I => \N__36871\
        );

    \I__8957\ : Span12Mux_v
    port map (
            O => \N__36915\,
            I => \N__36868\
        );

    \I__8956\ : Span12Mux_v
    port map (
            O => \N__36908\,
            I => \N__36865\
        );

    \I__8955\ : Sp12to4
    port map (
            O => \N__36905\,
            I => \N__36862\
        );

    \I__8954\ : Span4Mux_v
    port map (
            O => \N__36900\,
            I => \N__36859\
        );

    \I__8953\ : Span4Mux_v
    port map (
            O => \N__36891\,
            I => \N__36854\
        );

    \I__8952\ : LocalMux
    port map (
            O => \N__36888\,
            I => \N__36854\
        );

    \I__8951\ : Span4Mux_v
    port map (
            O => \N__36883\,
            I => \N__36851\
        );

    \I__8950\ : Span4Mux_v
    port map (
            O => \N__36880\,
            I => \N__36848\
        );

    \I__8949\ : Span4Mux_h
    port map (
            O => \N__36877\,
            I => \N__36844\
        );

    \I__8948\ : LocalMux
    port map (
            O => \N__36874\,
            I => \N__36841\
        );

    \I__8947\ : Span4Mux_h
    port map (
            O => \N__36871\,
            I => \N__36838\
        );

    \I__8946\ : Span12Mux_h
    port map (
            O => \N__36868\,
            I => \N__36831\
        );

    \I__8945\ : Span12Mux_h
    port map (
            O => \N__36865\,
            I => \N__36831\
        );

    \I__8944\ : Span12Mux_s11_v
    port map (
            O => \N__36862\,
            I => \N__36826\
        );

    \I__8943\ : Sp12to4
    port map (
            O => \N__36859\,
            I => \N__36826\
        );

    \I__8942\ : Span4Mux_v
    port map (
            O => \N__36854\,
            I => \N__36819\
        );

    \I__8941\ : Span4Mux_v
    port map (
            O => \N__36851\,
            I => \N__36819\
        );

    \I__8940\ : Span4Mux_h
    port map (
            O => \N__36848\,
            I => \N__36819\
        );

    \I__8939\ : SRMux
    port map (
            O => \N__36847\,
            I => \N__36816\
        );

    \I__8938\ : Span4Mux_h
    port map (
            O => \N__36844\,
            I => \N__36809\
        );

    \I__8937\ : Span4Mux_h
    port map (
            O => \N__36841\,
            I => \N__36809\
        );

    \I__8936\ : Span4Mux_v
    port map (
            O => \N__36838\,
            I => \N__36809\
        );

    \I__8935\ : SRMux
    port map (
            O => \N__36837\,
            I => \N__36806\
        );

    \I__8934\ : SRMux
    port map (
            O => \N__36836\,
            I => \N__36803\
        );

    \I__8933\ : Odrv12
    port map (
            O => \N__36831\,
            I => \CONSTANT_ONE_NET\
        );

    \I__8932\ : Odrv12
    port map (
            O => \N__36826\,
            I => \CONSTANT_ONE_NET\
        );

    \I__8931\ : Odrv4
    port map (
            O => \N__36819\,
            I => \CONSTANT_ONE_NET\
        );

    \I__8930\ : LocalMux
    port map (
            O => \N__36816\,
            I => \CONSTANT_ONE_NET\
        );

    \I__8929\ : Odrv4
    port map (
            O => \N__36809\,
            I => \CONSTANT_ONE_NET\
        );

    \I__8928\ : LocalMux
    port map (
            O => \N__36806\,
            I => \CONSTANT_ONE_NET\
        );

    \I__8927\ : LocalMux
    port map (
            O => \N__36803\,
            I => \CONSTANT_ONE_NET\
        );

    \I__8926\ : InMux
    port map (
            O => \N__36788\,
            I => \N__36784\
        );

    \I__8925\ : InMux
    port map (
            O => \N__36787\,
            I => \N__36781\
        );

    \I__8924\ : LocalMux
    port map (
            O => \N__36784\,
            I => \N__36777\
        );

    \I__8923\ : LocalMux
    port map (
            O => \N__36781\,
            I => \N__36773\
        );

    \I__8922\ : InMux
    port map (
            O => \N__36780\,
            I => \N__36770\
        );

    \I__8921\ : Span12Mux_h
    port map (
            O => \N__36777\,
            I => \N__36767\
        );

    \I__8920\ : InMux
    port map (
            O => \N__36776\,
            I => \N__36764\
        );

    \I__8919\ : Span4Mux_v
    port map (
            O => \N__36773\,
            I => \N__36759\
        );

    \I__8918\ : LocalMux
    port map (
            O => \N__36770\,
            I => \N__36759\
        );

    \I__8917\ : Odrv12
    port map (
            O => \N__36767\,
            I => \b2v_inst.dir_energiaZ0Z_10\
        );

    \I__8916\ : LocalMux
    port map (
            O => \N__36764\,
            I => \b2v_inst.dir_energiaZ0Z_10\
        );

    \I__8915\ : Odrv4
    port map (
            O => \N__36759\,
            I => \b2v_inst.dir_energiaZ0Z_10\
        );

    \I__8914\ : CascadeMux
    port map (
            O => \N__36752\,
            I => \N__36748\
        );

    \I__8913\ : InMux
    port map (
            O => \N__36751\,
            I => \N__36742\
        );

    \I__8912\ : InMux
    port map (
            O => \N__36748\,
            I => \N__36739\
        );

    \I__8911\ : InMux
    port map (
            O => \N__36747\,
            I => \N__36735\
        );

    \I__8910\ : CascadeMux
    port map (
            O => \N__36746\,
            I => \N__36732\
        );

    \I__8909\ : InMux
    port map (
            O => \N__36745\,
            I => \N__36729\
        );

    \I__8908\ : LocalMux
    port map (
            O => \N__36742\,
            I => \N__36723\
        );

    \I__8907\ : LocalMux
    port map (
            O => \N__36739\,
            I => \N__36720\
        );

    \I__8906\ : CascadeMux
    port map (
            O => \N__36738\,
            I => \N__36717\
        );

    \I__8905\ : LocalMux
    port map (
            O => \N__36735\,
            I => \N__36714\
        );

    \I__8904\ : InMux
    port map (
            O => \N__36732\,
            I => \N__36711\
        );

    \I__8903\ : LocalMux
    port map (
            O => \N__36729\,
            I => \N__36707\
        );

    \I__8902\ : InMux
    port map (
            O => \N__36728\,
            I => \N__36704\
        );

    \I__8901\ : InMux
    port map (
            O => \N__36727\,
            I => \N__36701\
        );

    \I__8900\ : CascadeMux
    port map (
            O => \N__36726\,
            I => \N__36698\
        );

    \I__8899\ : Span4Mux_v
    port map (
            O => \N__36723\,
            I => \N__36692\
        );

    \I__8898\ : Span4Mux_v
    port map (
            O => \N__36720\,
            I => \N__36692\
        );

    \I__8897\ : InMux
    port map (
            O => \N__36717\,
            I => \N__36689\
        );

    \I__8896\ : Span4Mux_v
    port map (
            O => \N__36714\,
            I => \N__36684\
        );

    \I__8895\ : LocalMux
    port map (
            O => \N__36711\,
            I => \N__36684\
        );

    \I__8894\ : InMux
    port map (
            O => \N__36710\,
            I => \N__36681\
        );

    \I__8893\ : Span4Mux_v
    port map (
            O => \N__36707\,
            I => \N__36674\
        );

    \I__8892\ : LocalMux
    port map (
            O => \N__36704\,
            I => \N__36674\
        );

    \I__8891\ : LocalMux
    port map (
            O => \N__36701\,
            I => \N__36674\
        );

    \I__8890\ : InMux
    port map (
            O => \N__36698\,
            I => \N__36671\
        );

    \I__8889\ : InMux
    port map (
            O => \N__36697\,
            I => \N__36668\
        );

    \I__8888\ : Sp12to4
    port map (
            O => \N__36692\,
            I => \N__36665\
        );

    \I__8887\ : LocalMux
    port map (
            O => \N__36689\,
            I => \N__36662\
        );

    \I__8886\ : Sp12to4
    port map (
            O => \N__36684\,
            I => \N__36657\
        );

    \I__8885\ : LocalMux
    port map (
            O => \N__36681\,
            I => \N__36657\
        );

    \I__8884\ : Span4Mux_h
    port map (
            O => \N__36674\,
            I => \N__36652\
        );

    \I__8883\ : LocalMux
    port map (
            O => \N__36671\,
            I => \N__36652\
        );

    \I__8882\ : LocalMux
    port map (
            O => \N__36668\,
            I => \N__36649\
        );

    \I__8881\ : Span12Mux_h
    port map (
            O => \N__36665\,
            I => \N__36644\
        );

    \I__8880\ : Sp12to4
    port map (
            O => \N__36662\,
            I => \N__36644\
        );

    \I__8879\ : Span12Mux_v
    port map (
            O => \N__36657\,
            I => \N__36641\
        );

    \I__8878\ : Span4Mux_h
    port map (
            O => \N__36652\,
            I => \N__36638\
        );

    \I__8877\ : Odrv4
    port map (
            O => \N__36649\,
            I => \b2v_inst.indiceZ0Z_10\
        );

    \I__8876\ : Odrv12
    port map (
            O => \N__36644\,
            I => \b2v_inst.indiceZ0Z_10\
        );

    \I__8875\ : Odrv12
    port map (
            O => \N__36641\,
            I => \b2v_inst.indiceZ0Z_10\
        );

    \I__8874\ : Odrv4
    port map (
            O => \N__36638\,
            I => \b2v_inst.indiceZ0Z_10\
        );

    \I__8873\ : CascadeMux
    port map (
            O => \N__36629\,
            I => \N__36626\
        );

    \I__8872\ : CascadeBuf
    port map (
            O => \N__36626\,
            I => \N__36622\
        );

    \I__8871\ : CascadeMux
    port map (
            O => \N__36625\,
            I => \N__36619\
        );

    \I__8870\ : CascadeMux
    port map (
            O => \N__36622\,
            I => \N__36616\
        );

    \I__8869\ : CascadeBuf
    port map (
            O => \N__36619\,
            I => \N__36613\
        );

    \I__8868\ : CascadeBuf
    port map (
            O => \N__36616\,
            I => \N__36610\
        );

    \I__8867\ : CascadeMux
    port map (
            O => \N__36613\,
            I => \N__36607\
        );

    \I__8866\ : CascadeMux
    port map (
            O => \N__36610\,
            I => \N__36604\
        );

    \I__8865\ : CascadeBuf
    port map (
            O => \N__36607\,
            I => \N__36601\
        );

    \I__8864\ : InMux
    port map (
            O => \N__36604\,
            I => \N__36598\
        );

    \I__8863\ : CascadeMux
    port map (
            O => \N__36601\,
            I => \N__36595\
        );

    \I__8862\ : LocalMux
    port map (
            O => \N__36598\,
            I => \N__36592\
        );

    \I__8861\ : InMux
    port map (
            O => \N__36595\,
            I => \N__36589\
        );

    \I__8860\ : Span4Mux_h
    port map (
            O => \N__36592\,
            I => \N__36586\
        );

    \I__8859\ : LocalMux
    port map (
            O => \N__36589\,
            I => \N_445_i\
        );

    \I__8858\ : Odrv4
    port map (
            O => \N__36586\,
            I => \N_445_i\
        );

    \I__8857\ : InMux
    port map (
            O => \N__36581\,
            I => \N__36577\
        );

    \I__8856\ : InMux
    port map (
            O => \N__36580\,
            I => \N__36574\
        );

    \I__8855\ : LocalMux
    port map (
            O => \N__36577\,
            I => \N__36566\
        );

    \I__8854\ : LocalMux
    port map (
            O => \N__36574\,
            I => \N__36562\
        );

    \I__8853\ : InMux
    port map (
            O => \N__36573\,
            I => \N__36559\
        );

    \I__8852\ : InMux
    port map (
            O => \N__36572\,
            I => \N__36556\
        );

    \I__8851\ : InMux
    port map (
            O => \N__36571\,
            I => \N__36553\
        );

    \I__8850\ : InMux
    port map (
            O => \N__36570\,
            I => \N__36550\
        );

    \I__8849\ : InMux
    port map (
            O => \N__36569\,
            I => \N__36547\
        );

    \I__8848\ : Sp12to4
    port map (
            O => \N__36566\,
            I => \N__36544\
        );

    \I__8847\ : InMux
    port map (
            O => \N__36565\,
            I => \N__36541\
        );

    \I__8846\ : Span4Mux_v
    port map (
            O => \N__36562\,
            I => \N__36536\
        );

    \I__8845\ : LocalMux
    port map (
            O => \N__36559\,
            I => \N__36536\
        );

    \I__8844\ : LocalMux
    port map (
            O => \N__36556\,
            I => \N__36531\
        );

    \I__8843\ : LocalMux
    port map (
            O => \N__36553\,
            I => \N__36531\
        );

    \I__8842\ : LocalMux
    port map (
            O => \N__36550\,
            I => \N__36528\
        );

    \I__8841\ : LocalMux
    port map (
            O => \N__36547\,
            I => \N__36524\
        );

    \I__8840\ : Span12Mux_v
    port map (
            O => \N__36544\,
            I => \N__36520\
        );

    \I__8839\ : LocalMux
    port map (
            O => \N__36541\,
            I => \N__36513\
        );

    \I__8838\ : Span4Mux_v
    port map (
            O => \N__36536\,
            I => \N__36513\
        );

    \I__8837\ : Span4Mux_h
    port map (
            O => \N__36531\,
            I => \N__36513\
        );

    \I__8836\ : Span4Mux_h
    port map (
            O => \N__36528\,
            I => \N__36509\
        );

    \I__8835\ : InMux
    port map (
            O => \N__36527\,
            I => \N__36506\
        );

    \I__8834\ : Span4Mux_v
    port map (
            O => \N__36524\,
            I => \N__36503\
        );

    \I__8833\ : InMux
    port map (
            O => \N__36523\,
            I => \N__36500\
        );

    \I__8832\ : Span12Mux_h
    port map (
            O => \N__36520\,
            I => \N__36496\
        );

    \I__8831\ : Span4Mux_h
    port map (
            O => \N__36513\,
            I => \N__36493\
        );

    \I__8830\ : InMux
    port map (
            O => \N__36512\,
            I => \N__36490\
        );

    \I__8829\ : Span4Mux_v
    port map (
            O => \N__36509\,
            I => \N__36481\
        );

    \I__8828\ : LocalMux
    port map (
            O => \N__36506\,
            I => \N__36481\
        );

    \I__8827\ : Span4Mux_h
    port map (
            O => \N__36503\,
            I => \N__36481\
        );

    \I__8826\ : LocalMux
    port map (
            O => \N__36500\,
            I => \N__36481\
        );

    \I__8825\ : InMux
    port map (
            O => \N__36499\,
            I => \N__36478\
        );

    \I__8824\ : Odrv12
    port map (
            O => \N__36496\,
            I => \b2v_inst.indiceZ0Z_3\
        );

    \I__8823\ : Odrv4
    port map (
            O => \N__36493\,
            I => \b2v_inst.indiceZ0Z_3\
        );

    \I__8822\ : LocalMux
    port map (
            O => \N__36490\,
            I => \b2v_inst.indiceZ0Z_3\
        );

    \I__8821\ : Odrv4
    port map (
            O => \N__36481\,
            I => \b2v_inst.indiceZ0Z_3\
        );

    \I__8820\ : LocalMux
    port map (
            O => \N__36478\,
            I => \b2v_inst.indiceZ0Z_3\
        );

    \I__8819\ : CascadeMux
    port map (
            O => \N__36467\,
            I => \N__36464\
        );

    \I__8818\ : InMux
    port map (
            O => \N__36464\,
            I => \N__36460\
        );

    \I__8817\ : InMux
    port map (
            O => \N__36463\,
            I => \N__36457\
        );

    \I__8816\ : LocalMux
    port map (
            O => \N__36460\,
            I => \N__36454\
        );

    \I__8815\ : LocalMux
    port map (
            O => \N__36457\,
            I => \N__36450\
        );

    \I__8814\ : Span12Mux_v
    port map (
            O => \N__36454\,
            I => \N__36445\
        );

    \I__8813\ : InMux
    port map (
            O => \N__36453\,
            I => \N__36442\
        );

    \I__8812\ : Span4Mux_v
    port map (
            O => \N__36450\,
            I => \N__36439\
        );

    \I__8811\ : InMux
    port map (
            O => \N__36449\,
            I => \N__36436\
        );

    \I__8810\ : InMux
    port map (
            O => \N__36448\,
            I => \N__36433\
        );

    \I__8809\ : Odrv12
    port map (
            O => \N__36445\,
            I => \b2v_inst.dir_energiaZ0Z_3\
        );

    \I__8808\ : LocalMux
    port map (
            O => \N__36442\,
            I => \b2v_inst.dir_energiaZ0Z_3\
        );

    \I__8807\ : Odrv4
    port map (
            O => \N__36439\,
            I => \b2v_inst.dir_energiaZ0Z_3\
        );

    \I__8806\ : LocalMux
    port map (
            O => \N__36436\,
            I => \b2v_inst.dir_energiaZ0Z_3\
        );

    \I__8805\ : LocalMux
    port map (
            O => \N__36433\,
            I => \b2v_inst.dir_energiaZ0Z_3\
        );

    \I__8804\ : CascadeMux
    port map (
            O => \N__36422\,
            I => \N__36418\
        );

    \I__8803\ : CascadeMux
    port map (
            O => \N__36421\,
            I => \N__36415\
        );

    \I__8802\ : CascadeBuf
    port map (
            O => \N__36418\,
            I => \N__36412\
        );

    \I__8801\ : CascadeBuf
    port map (
            O => \N__36415\,
            I => \N__36409\
        );

    \I__8800\ : CascadeMux
    port map (
            O => \N__36412\,
            I => \N__36406\
        );

    \I__8799\ : CascadeMux
    port map (
            O => \N__36409\,
            I => \N__36403\
        );

    \I__8798\ : CascadeBuf
    port map (
            O => \N__36406\,
            I => \N__36400\
        );

    \I__8797\ : CascadeBuf
    port map (
            O => \N__36403\,
            I => \N__36397\
        );

    \I__8796\ : CascadeMux
    port map (
            O => \N__36400\,
            I => \N__36394\
        );

    \I__8795\ : CascadeMux
    port map (
            O => \N__36397\,
            I => \N__36391\
        );

    \I__8794\ : InMux
    port map (
            O => \N__36394\,
            I => \N__36388\
        );

    \I__8793\ : InMux
    port map (
            O => \N__36391\,
            I => \N__36385\
        );

    \I__8792\ : LocalMux
    port map (
            O => \N__36388\,
            I => \N__36382\
        );

    \I__8791\ : LocalMux
    port map (
            O => \N__36385\,
            I => \N_357_i\
        );

    \I__8790\ : Odrv4
    port map (
            O => \N__36382\,
            I => \N_357_i\
        );

    \I__8789\ : InMux
    port map (
            O => \N__36377\,
            I => \N__36372\
        );

    \I__8788\ : InMux
    port map (
            O => \N__36376\,
            I => \N__36369\
        );

    \I__8787\ : CascadeMux
    port map (
            O => \N__36375\,
            I => \N__36364\
        );

    \I__8786\ : LocalMux
    port map (
            O => \N__36372\,
            I => \N__36360\
        );

    \I__8785\ : LocalMux
    port map (
            O => \N__36369\,
            I => \N__36354\
        );

    \I__8784\ : InMux
    port map (
            O => \N__36368\,
            I => \N__36351\
        );

    \I__8783\ : InMux
    port map (
            O => \N__36367\,
            I => \N__36348\
        );

    \I__8782\ : InMux
    port map (
            O => \N__36364\,
            I => \N__36344\
        );

    \I__8781\ : InMux
    port map (
            O => \N__36363\,
            I => \N__36341\
        );

    \I__8780\ : Span4Mux_v
    port map (
            O => \N__36360\,
            I => \N__36338\
        );

    \I__8779\ : InMux
    port map (
            O => \N__36359\,
            I => \N__36334\
        );

    \I__8778\ : InMux
    port map (
            O => \N__36358\,
            I => \N__36331\
        );

    \I__8777\ : InMux
    port map (
            O => \N__36357\,
            I => \N__36328\
        );

    \I__8776\ : Sp12to4
    port map (
            O => \N__36354\,
            I => \N__36325\
        );

    \I__8775\ : LocalMux
    port map (
            O => \N__36351\,
            I => \N__36322\
        );

    \I__8774\ : LocalMux
    port map (
            O => \N__36348\,
            I => \N__36319\
        );

    \I__8773\ : InMux
    port map (
            O => \N__36347\,
            I => \N__36316\
        );

    \I__8772\ : LocalMux
    port map (
            O => \N__36344\,
            I => \N__36313\
        );

    \I__8771\ : LocalMux
    port map (
            O => \N__36341\,
            I => \N__36310\
        );

    \I__8770\ : Span4Mux_v
    port map (
            O => \N__36338\,
            I => \N__36306\
        );

    \I__8769\ : InMux
    port map (
            O => \N__36337\,
            I => \N__36303\
        );

    \I__8768\ : LocalMux
    port map (
            O => \N__36334\,
            I => \N__36296\
        );

    \I__8767\ : LocalMux
    port map (
            O => \N__36331\,
            I => \N__36296\
        );

    \I__8766\ : LocalMux
    port map (
            O => \N__36328\,
            I => \N__36296\
        );

    \I__8765\ : Span12Mux_v
    port map (
            O => \N__36325\,
            I => \N__36293\
        );

    \I__8764\ : Span4Mux_v
    port map (
            O => \N__36322\,
            I => \N__36286\
        );

    \I__8763\ : Span4Mux_v
    port map (
            O => \N__36319\,
            I => \N__36286\
        );

    \I__8762\ : LocalMux
    port map (
            O => \N__36316\,
            I => \N__36286\
        );

    \I__8761\ : Span4Mux_v
    port map (
            O => \N__36313\,
            I => \N__36283\
        );

    \I__8760\ : Span4Mux_v
    port map (
            O => \N__36310\,
            I => \N__36280\
        );

    \I__8759\ : InMux
    port map (
            O => \N__36309\,
            I => \N__36277\
        );

    \I__8758\ : Span4Mux_v
    port map (
            O => \N__36306\,
            I => \N__36270\
        );

    \I__8757\ : LocalMux
    port map (
            O => \N__36303\,
            I => \N__36270\
        );

    \I__8756\ : Span4Mux_v
    port map (
            O => \N__36296\,
            I => \N__36270\
        );

    \I__8755\ : Odrv12
    port map (
            O => \N__36293\,
            I => \b2v_inst.indiceZ0Z_4\
        );

    \I__8754\ : Odrv4
    port map (
            O => \N__36286\,
            I => \b2v_inst.indiceZ0Z_4\
        );

    \I__8753\ : Odrv4
    port map (
            O => \N__36283\,
            I => \b2v_inst.indiceZ0Z_4\
        );

    \I__8752\ : Odrv4
    port map (
            O => \N__36280\,
            I => \b2v_inst.indiceZ0Z_4\
        );

    \I__8751\ : LocalMux
    port map (
            O => \N__36277\,
            I => \b2v_inst.indiceZ0Z_4\
        );

    \I__8750\ : Odrv4
    port map (
            O => \N__36270\,
            I => \b2v_inst.indiceZ0Z_4\
        );

    \I__8749\ : CascadeMux
    port map (
            O => \N__36257\,
            I => \N__36254\
        );

    \I__8748\ : InMux
    port map (
            O => \N__36254\,
            I => \N__36251\
        );

    \I__8747\ : LocalMux
    port map (
            O => \N__36251\,
            I => \N__36248\
        );

    \I__8746\ : Span4Mux_v
    port map (
            O => \N__36248\,
            I => \N__36243\
        );

    \I__8745\ : InMux
    port map (
            O => \N__36247\,
            I => \N__36240\
        );

    \I__8744\ : InMux
    port map (
            O => \N__36246\,
            I => \N__36237\
        );

    \I__8743\ : Span4Mux_h
    port map (
            O => \N__36243\,
            I => \N__36233\
        );

    \I__8742\ : LocalMux
    port map (
            O => \N__36240\,
            I => \N__36230\
        );

    \I__8741\ : LocalMux
    port map (
            O => \N__36237\,
            I => \N__36227\
        );

    \I__8740\ : InMux
    port map (
            O => \N__36236\,
            I => \N__36224\
        );

    \I__8739\ : Span4Mux_h
    port map (
            O => \N__36233\,
            I => \N__36219\
        );

    \I__8738\ : Span4Mux_v
    port map (
            O => \N__36230\,
            I => \N__36219\
        );

    \I__8737\ : Span4Mux_v
    port map (
            O => \N__36227\,
            I => \N__36214\
        );

    \I__8736\ : LocalMux
    port map (
            O => \N__36224\,
            I => \N__36214\
        );

    \I__8735\ : Odrv4
    port map (
            O => \N__36219\,
            I => \b2v_inst.dir_energiaZ0Z_4\
        );

    \I__8734\ : Odrv4
    port map (
            O => \N__36214\,
            I => \b2v_inst.dir_energiaZ0Z_4\
        );

    \I__8733\ : CascadeMux
    port map (
            O => \N__36209\,
            I => \N__36205\
        );

    \I__8732\ : CascadeMux
    port map (
            O => \N__36208\,
            I => \N__36202\
        );

    \I__8731\ : CascadeBuf
    port map (
            O => \N__36205\,
            I => \N__36199\
        );

    \I__8730\ : CascadeBuf
    port map (
            O => \N__36202\,
            I => \N__36196\
        );

    \I__8729\ : CascadeMux
    port map (
            O => \N__36199\,
            I => \N__36193\
        );

    \I__8728\ : CascadeMux
    port map (
            O => \N__36196\,
            I => \N__36190\
        );

    \I__8727\ : CascadeBuf
    port map (
            O => \N__36193\,
            I => \N__36187\
        );

    \I__8726\ : CascadeBuf
    port map (
            O => \N__36190\,
            I => \N__36184\
        );

    \I__8725\ : CascadeMux
    port map (
            O => \N__36187\,
            I => \N__36181\
        );

    \I__8724\ : CascadeMux
    port map (
            O => \N__36184\,
            I => \N__36178\
        );

    \I__8723\ : InMux
    port map (
            O => \N__36181\,
            I => \N__36175\
        );

    \I__8722\ : InMux
    port map (
            O => \N__36178\,
            I => \N__36172\
        );

    \I__8721\ : LocalMux
    port map (
            O => \N__36175\,
            I => \N__36169\
        );

    \I__8720\ : LocalMux
    port map (
            O => \N__36172\,
            I => \N_356_i\
        );

    \I__8719\ : Odrv4
    port map (
            O => \N__36169\,
            I => \N_356_i\
        );

    \I__8718\ : CascadeMux
    port map (
            O => \N__36164\,
            I => \N__36161\
        );

    \I__8717\ : InMux
    port map (
            O => \N__36161\,
            I => \N__36158\
        );

    \I__8716\ : LocalMux
    port map (
            O => \N__36158\,
            I => \N__36155\
        );

    \I__8715\ : Span4Mux_v
    port map (
            O => \N__36155\,
            I => \N__36151\
        );

    \I__8714\ : InMux
    port map (
            O => \N__36154\,
            I => \N__36148\
        );

    \I__8713\ : Span4Mux_h
    port map (
            O => \N__36151\,
            I => \N__36143\
        );

    \I__8712\ : LocalMux
    port map (
            O => \N__36148\,
            I => \N__36140\
        );

    \I__8711\ : InMux
    port map (
            O => \N__36147\,
            I => \N__36137\
        );

    \I__8710\ : InMux
    port map (
            O => \N__36146\,
            I => \N__36134\
        );

    \I__8709\ : Span4Mux_h
    port map (
            O => \N__36143\,
            I => \N__36127\
        );

    \I__8708\ : Span4Mux_v
    port map (
            O => \N__36140\,
            I => \N__36127\
        );

    \I__8707\ : LocalMux
    port map (
            O => \N__36137\,
            I => \N__36127\
        );

    \I__8706\ : LocalMux
    port map (
            O => \N__36134\,
            I => \b2v_inst.dir_energiaZ0Z_2\
        );

    \I__8705\ : Odrv4
    port map (
            O => \N__36127\,
            I => \b2v_inst.dir_energiaZ0Z_2\
        );

    \I__8704\ : InMux
    port map (
            O => \N__36122\,
            I => \N__36118\
        );

    \I__8703\ : InMux
    port map (
            O => \N__36121\,
            I => \N__36115\
        );

    \I__8702\ : LocalMux
    port map (
            O => \N__36118\,
            I => \N__36110\
        );

    \I__8701\ : LocalMux
    port map (
            O => \N__36115\,
            I => \N__36107\
        );

    \I__8700\ : InMux
    port map (
            O => \N__36114\,
            I => \N__36104\
        );

    \I__8699\ : CascadeMux
    port map (
            O => \N__36113\,
            I => \N__36100\
        );

    \I__8698\ : Span4Mux_h
    port map (
            O => \N__36110\,
            I => \N__36097\
        );

    \I__8697\ : Span4Mux_h
    port map (
            O => \N__36107\,
            I => \N__36093\
        );

    \I__8696\ : LocalMux
    port map (
            O => \N__36104\,
            I => \N__36089\
        );

    \I__8695\ : InMux
    port map (
            O => \N__36103\,
            I => \N__36086\
        );

    \I__8694\ : InMux
    port map (
            O => \N__36100\,
            I => \N__36083\
        );

    \I__8693\ : Span4Mux_h
    port map (
            O => \N__36097\,
            I => \N__36080\
        );

    \I__8692\ : InMux
    port map (
            O => \N__36096\,
            I => \N__36077\
        );

    \I__8691\ : Span4Mux_h
    port map (
            O => \N__36093\,
            I => \N__36073\
        );

    \I__8690\ : InMux
    port map (
            O => \N__36092\,
            I => \N__36070\
        );

    \I__8689\ : Span4Mux_v
    port map (
            O => \N__36089\,
            I => \N__36067\
        );

    \I__8688\ : LocalMux
    port map (
            O => \N__36086\,
            I => \N__36064\
        );

    \I__8687\ : LocalMux
    port map (
            O => \N__36083\,
            I => \N__36057\
        );

    \I__8686\ : Span4Mux_v
    port map (
            O => \N__36080\,
            I => \N__36057\
        );

    \I__8685\ : LocalMux
    port map (
            O => \N__36077\,
            I => \N__36057\
        );

    \I__8684\ : CascadeMux
    port map (
            O => \N__36076\,
            I => \N__36054\
        );

    \I__8683\ : Sp12to4
    port map (
            O => \N__36073\,
            I => \N__36051\
        );

    \I__8682\ : LocalMux
    port map (
            O => \N__36070\,
            I => \N__36045\
        );

    \I__8681\ : Span4Mux_h
    port map (
            O => \N__36067\,
            I => \N__36045\
        );

    \I__8680\ : Span4Mux_h
    port map (
            O => \N__36064\,
            I => \N__36040\
        );

    \I__8679\ : Span4Mux_v
    port map (
            O => \N__36057\,
            I => \N__36037\
        );

    \I__8678\ : InMux
    port map (
            O => \N__36054\,
            I => \N__36034\
        );

    \I__8677\ : Span12Mux_v
    port map (
            O => \N__36051\,
            I => \N__36031\
        );

    \I__8676\ : InMux
    port map (
            O => \N__36050\,
            I => \N__36028\
        );

    \I__8675\ : Span4Mux_v
    port map (
            O => \N__36045\,
            I => \N__36025\
        );

    \I__8674\ : InMux
    port map (
            O => \N__36044\,
            I => \N__36022\
        );

    \I__8673\ : InMux
    port map (
            O => \N__36043\,
            I => \N__36019\
        );

    \I__8672\ : Span4Mux_v
    port map (
            O => \N__36040\,
            I => \N__36012\
        );

    \I__8671\ : Span4Mux_h
    port map (
            O => \N__36037\,
            I => \N__36012\
        );

    \I__8670\ : LocalMux
    port map (
            O => \N__36034\,
            I => \N__36012\
        );

    \I__8669\ : Odrv12
    port map (
            O => \N__36031\,
            I => \b2v_inst.indiceZ0Z_2\
        );

    \I__8668\ : LocalMux
    port map (
            O => \N__36028\,
            I => \b2v_inst.indiceZ0Z_2\
        );

    \I__8667\ : Odrv4
    port map (
            O => \N__36025\,
            I => \b2v_inst.indiceZ0Z_2\
        );

    \I__8666\ : LocalMux
    port map (
            O => \N__36022\,
            I => \b2v_inst.indiceZ0Z_2\
        );

    \I__8665\ : LocalMux
    port map (
            O => \N__36019\,
            I => \b2v_inst.indiceZ0Z_2\
        );

    \I__8664\ : Odrv4
    port map (
            O => \N__36012\,
            I => \b2v_inst.indiceZ0Z_2\
        );

    \I__8663\ : CascadeMux
    port map (
            O => \N__35999\,
            I => \N__35995\
        );

    \I__8662\ : CascadeMux
    port map (
            O => \N__35998\,
            I => \N__35992\
        );

    \I__8661\ : CascadeBuf
    port map (
            O => \N__35995\,
            I => \N__35989\
        );

    \I__8660\ : CascadeBuf
    port map (
            O => \N__35992\,
            I => \N__35986\
        );

    \I__8659\ : CascadeMux
    port map (
            O => \N__35989\,
            I => \N__35983\
        );

    \I__8658\ : CascadeMux
    port map (
            O => \N__35986\,
            I => \N__35980\
        );

    \I__8657\ : CascadeBuf
    port map (
            O => \N__35983\,
            I => \N__35977\
        );

    \I__8656\ : CascadeBuf
    port map (
            O => \N__35980\,
            I => \N__35974\
        );

    \I__8655\ : CascadeMux
    port map (
            O => \N__35977\,
            I => \N__35971\
        );

    \I__8654\ : CascadeMux
    port map (
            O => \N__35974\,
            I => \N__35968\
        );

    \I__8653\ : InMux
    port map (
            O => \N__35971\,
            I => \N__35965\
        );

    \I__8652\ : InMux
    port map (
            O => \N__35968\,
            I => \N__35962\
        );

    \I__8651\ : LocalMux
    port map (
            O => \N__35965\,
            I => \N__35959\
        );

    \I__8650\ : LocalMux
    port map (
            O => \N__35962\,
            I => \N_358_i\
        );

    \I__8649\ : Odrv4
    port map (
            O => \N__35959\,
            I => \N_358_i\
        );

    \I__8648\ : CascadeMux
    port map (
            O => \N__35954\,
            I => \N__35949\
        );

    \I__8647\ : InMux
    port map (
            O => \N__35953\,
            I => \N__35946\
        );

    \I__8646\ : CascadeMux
    port map (
            O => \N__35952\,
            I => \N__35943\
        );

    \I__8645\ : InMux
    port map (
            O => \N__35949\,
            I => \N__35940\
        );

    \I__8644\ : LocalMux
    port map (
            O => \N__35946\,
            I => \N__35934\
        );

    \I__8643\ : InMux
    port map (
            O => \N__35943\,
            I => \N__35930\
        );

    \I__8642\ : LocalMux
    port map (
            O => \N__35940\,
            I => \N__35927\
        );

    \I__8641\ : InMux
    port map (
            O => \N__35939\,
            I => \N__35924\
        );

    \I__8640\ : InMux
    port map (
            O => \N__35938\,
            I => \N__35921\
        );

    \I__8639\ : InMux
    port map (
            O => \N__35937\,
            I => \N__35916\
        );

    \I__8638\ : Span4Mux_v
    port map (
            O => \N__35934\,
            I => \N__35912\
        );

    \I__8637\ : InMux
    port map (
            O => \N__35933\,
            I => \N__35907\
        );

    \I__8636\ : LocalMux
    port map (
            O => \N__35930\,
            I => \N__35904\
        );

    \I__8635\ : Span4Mux_h
    port map (
            O => \N__35927\,
            I => \N__35897\
        );

    \I__8634\ : LocalMux
    port map (
            O => \N__35924\,
            I => \N__35897\
        );

    \I__8633\ : LocalMux
    port map (
            O => \N__35921\,
            I => \N__35897\
        );

    \I__8632\ : InMux
    port map (
            O => \N__35920\,
            I => \N__35892\
        );

    \I__8631\ : InMux
    port map (
            O => \N__35919\,
            I => \N__35892\
        );

    \I__8630\ : LocalMux
    port map (
            O => \N__35916\,
            I => \N__35889\
        );

    \I__8629\ : InMux
    port map (
            O => \N__35915\,
            I => \N__35886\
        );

    \I__8628\ : Span4Mux_h
    port map (
            O => \N__35912\,
            I => \N__35883\
        );

    \I__8627\ : InMux
    port map (
            O => \N__35911\,
            I => \N__35880\
        );

    \I__8626\ : InMux
    port map (
            O => \N__35910\,
            I => \N__35877\
        );

    \I__8625\ : LocalMux
    port map (
            O => \N__35907\,
            I => \N__35874\
        );

    \I__8624\ : Span4Mux_h
    port map (
            O => \N__35904\,
            I => \N__35871\
        );

    \I__8623\ : Span4Mux_v
    port map (
            O => \N__35897\,
            I => \N__35866\
        );

    \I__8622\ : LocalMux
    port map (
            O => \N__35892\,
            I => \N__35866\
        );

    \I__8621\ : Span4Mux_v
    port map (
            O => \N__35889\,
            I => \N__35863\
        );

    \I__8620\ : LocalMux
    port map (
            O => \N__35886\,
            I => \N__35860\
        );

    \I__8619\ : Span4Mux_h
    port map (
            O => \N__35883\,
            I => \N__35857\
        );

    \I__8618\ : LocalMux
    port map (
            O => \N__35880\,
            I => \N__35854\
        );

    \I__8617\ : LocalMux
    port map (
            O => \N__35877\,
            I => \N__35847\
        );

    \I__8616\ : Span12Mux_h
    port map (
            O => \N__35874\,
            I => \N__35847\
        );

    \I__8615\ : Sp12to4
    port map (
            O => \N__35871\,
            I => \N__35847\
        );

    \I__8614\ : Span4Mux_h
    port map (
            O => \N__35866\,
            I => \N__35844\
        );

    \I__8613\ : Odrv4
    port map (
            O => \N__35863\,
            I => \b2v_inst.indiceZ0Z_9\
        );

    \I__8612\ : Odrv12
    port map (
            O => \N__35860\,
            I => \b2v_inst.indiceZ0Z_9\
        );

    \I__8611\ : Odrv4
    port map (
            O => \N__35857\,
            I => \b2v_inst.indiceZ0Z_9\
        );

    \I__8610\ : Odrv4
    port map (
            O => \N__35854\,
            I => \b2v_inst.indiceZ0Z_9\
        );

    \I__8609\ : Odrv12
    port map (
            O => \N__35847\,
            I => \b2v_inst.indiceZ0Z_9\
        );

    \I__8608\ : Odrv4
    port map (
            O => \N__35844\,
            I => \b2v_inst.indiceZ0Z_9\
        );

    \I__8607\ : CascadeMux
    port map (
            O => \N__35831\,
            I => \N__35828\
        );

    \I__8606\ : InMux
    port map (
            O => \N__35828\,
            I => \N__35824\
        );

    \I__8605\ : CascadeMux
    port map (
            O => \N__35827\,
            I => \N__35820\
        );

    \I__8604\ : LocalMux
    port map (
            O => \N__35824\,
            I => \N__35816\
        );

    \I__8603\ : InMux
    port map (
            O => \N__35823\,
            I => \N__35813\
        );

    \I__8602\ : InMux
    port map (
            O => \N__35820\,
            I => \N__35809\
        );

    \I__8601\ : InMux
    port map (
            O => \N__35819\,
            I => \N__35806\
        );

    \I__8600\ : Span4Mux_v
    port map (
            O => \N__35816\,
            I => \N__35803\
        );

    \I__8599\ : LocalMux
    port map (
            O => \N__35813\,
            I => \N__35800\
        );

    \I__8598\ : CascadeMux
    port map (
            O => \N__35812\,
            I => \N__35797\
        );

    \I__8597\ : LocalMux
    port map (
            O => \N__35809\,
            I => \N__35792\
        );

    \I__8596\ : LocalMux
    port map (
            O => \N__35806\,
            I => \N__35792\
        );

    \I__8595\ : Sp12to4
    port map (
            O => \N__35803\,
            I => \N__35789\
        );

    \I__8594\ : Span4Mux_h
    port map (
            O => \N__35800\,
            I => \N__35786\
        );

    \I__8593\ : InMux
    port map (
            O => \N__35797\,
            I => \N__35783\
        );

    \I__8592\ : Span4Mux_h
    port map (
            O => \N__35792\,
            I => \N__35780\
        );

    \I__8591\ : Odrv12
    port map (
            O => \N__35789\,
            I => \b2v_inst.dir_energiaZ0Z_9\
        );

    \I__8590\ : Odrv4
    port map (
            O => \N__35786\,
            I => \b2v_inst.dir_energiaZ0Z_9\
        );

    \I__8589\ : LocalMux
    port map (
            O => \N__35783\,
            I => \b2v_inst.dir_energiaZ0Z_9\
        );

    \I__8588\ : Odrv4
    port map (
            O => \N__35780\,
            I => \b2v_inst.dir_energiaZ0Z_9\
        );

    \I__8587\ : CascadeMux
    port map (
            O => \N__35771\,
            I => \N__35767\
        );

    \I__8586\ : CascadeMux
    port map (
            O => \N__35770\,
            I => \N__35764\
        );

    \I__8585\ : CascadeBuf
    port map (
            O => \N__35767\,
            I => \N__35761\
        );

    \I__8584\ : CascadeBuf
    port map (
            O => \N__35764\,
            I => \N__35758\
        );

    \I__8583\ : CascadeMux
    port map (
            O => \N__35761\,
            I => \N__35755\
        );

    \I__8582\ : CascadeMux
    port map (
            O => \N__35758\,
            I => \N__35752\
        );

    \I__8581\ : CascadeBuf
    port map (
            O => \N__35755\,
            I => \N__35749\
        );

    \I__8580\ : CascadeBuf
    port map (
            O => \N__35752\,
            I => \N__35746\
        );

    \I__8579\ : CascadeMux
    port map (
            O => \N__35749\,
            I => \N__35743\
        );

    \I__8578\ : CascadeMux
    port map (
            O => \N__35746\,
            I => \N__35740\
        );

    \I__8577\ : InMux
    port map (
            O => \N__35743\,
            I => \N__35737\
        );

    \I__8576\ : InMux
    port map (
            O => \N__35740\,
            I => \N__35734\
        );

    \I__8575\ : LocalMux
    port map (
            O => \N__35737\,
            I => \N__35731\
        );

    \I__8574\ : LocalMux
    port map (
            O => \N__35734\,
            I => \N_444_i\
        );

    \I__8573\ : Odrv4
    port map (
            O => \N__35731\,
            I => \N_444_i\
        );

    \I__8572\ : InMux
    port map (
            O => \N__35726\,
            I => \N__35723\
        );

    \I__8571\ : LocalMux
    port map (
            O => \N__35723\,
            I => \N__35719\
        );

    \I__8570\ : InMux
    port map (
            O => \N__35722\,
            I => \N__35716\
        );

    \I__8569\ : Span4Mux_h
    port map (
            O => \N__35719\,
            I => \N__35712\
        );

    \I__8568\ : LocalMux
    port map (
            O => \N__35716\,
            I => \N__35707\
        );

    \I__8567\ : CascadeMux
    port map (
            O => \N__35715\,
            I => \N__35702\
        );

    \I__8566\ : Span4Mux_h
    port map (
            O => \N__35712\,
            I => \N__35697\
        );

    \I__8565\ : InMux
    port map (
            O => \N__35711\,
            I => \N__35694\
        );

    \I__8564\ : InMux
    port map (
            O => \N__35710\,
            I => \N__35691\
        );

    \I__8563\ : Span4Mux_v
    port map (
            O => \N__35707\,
            I => \N__35687\
        );

    \I__8562\ : InMux
    port map (
            O => \N__35706\,
            I => \N__35684\
        );

    \I__8561\ : InMux
    port map (
            O => \N__35705\,
            I => \N__35679\
        );

    \I__8560\ : InMux
    port map (
            O => \N__35702\,
            I => \N__35676\
        );

    \I__8559\ : InMux
    port map (
            O => \N__35701\,
            I => \N__35673\
        );

    \I__8558\ : InMux
    port map (
            O => \N__35700\,
            I => \N__35670\
        );

    \I__8557\ : Span4Mux_v
    port map (
            O => \N__35697\,
            I => \N__35664\
        );

    \I__8556\ : LocalMux
    port map (
            O => \N__35694\,
            I => \N__35664\
        );

    \I__8555\ : LocalMux
    port map (
            O => \N__35691\,
            I => \N__35661\
        );

    \I__8554\ : InMux
    port map (
            O => \N__35690\,
            I => \N__35658\
        );

    \I__8553\ : Sp12to4
    port map (
            O => \N__35687\,
            I => \N__35655\
        );

    \I__8552\ : LocalMux
    port map (
            O => \N__35684\,
            I => \N__35652\
        );

    \I__8551\ : InMux
    port map (
            O => \N__35683\,
            I => \N__35649\
        );

    \I__8550\ : InMux
    port map (
            O => \N__35682\,
            I => \N__35646\
        );

    \I__8549\ : LocalMux
    port map (
            O => \N__35679\,
            I => \N__35641\
        );

    \I__8548\ : LocalMux
    port map (
            O => \N__35676\,
            I => \N__35641\
        );

    \I__8547\ : LocalMux
    port map (
            O => \N__35673\,
            I => \N__35636\
        );

    \I__8546\ : LocalMux
    port map (
            O => \N__35670\,
            I => \N__35636\
        );

    \I__8545\ : InMux
    port map (
            O => \N__35669\,
            I => \N__35633\
        );

    \I__8544\ : Span4Mux_h
    port map (
            O => \N__35664\,
            I => \N__35626\
        );

    \I__8543\ : Span4Mux_h
    port map (
            O => \N__35661\,
            I => \N__35626\
        );

    \I__8542\ : LocalMux
    port map (
            O => \N__35658\,
            I => \N__35626\
        );

    \I__8541\ : Span12Mux_h
    port map (
            O => \N__35655\,
            I => \N__35621\
        );

    \I__8540\ : Sp12to4
    port map (
            O => \N__35652\,
            I => \N__35621\
        );

    \I__8539\ : LocalMux
    port map (
            O => \N__35649\,
            I => \N__35618\
        );

    \I__8538\ : LocalMux
    port map (
            O => \N__35646\,
            I => \N__35615\
        );

    \I__8537\ : Span4Mux_v
    port map (
            O => \N__35641\,
            I => \N__35608\
        );

    \I__8536\ : Span4Mux_h
    port map (
            O => \N__35636\,
            I => \N__35608\
        );

    \I__8535\ : LocalMux
    port map (
            O => \N__35633\,
            I => \N__35608\
        );

    \I__8534\ : Span4Mux_h
    port map (
            O => \N__35626\,
            I => \N__35605\
        );

    \I__8533\ : Odrv12
    port map (
            O => \N__35621\,
            I => \b2v_inst.indiceZ0Z_5\
        );

    \I__8532\ : Odrv4
    port map (
            O => \N__35618\,
            I => \b2v_inst.indiceZ0Z_5\
        );

    \I__8531\ : Odrv4
    port map (
            O => \N__35615\,
            I => \b2v_inst.indiceZ0Z_5\
        );

    \I__8530\ : Odrv4
    port map (
            O => \N__35608\,
            I => \b2v_inst.indiceZ0Z_5\
        );

    \I__8529\ : Odrv4
    port map (
            O => \N__35605\,
            I => \b2v_inst.indiceZ0Z_5\
        );

    \I__8528\ : CascadeMux
    port map (
            O => \N__35594\,
            I => \N__35591\
        );

    \I__8527\ : InMux
    port map (
            O => \N__35591\,
            I => \N__35588\
        );

    \I__8526\ : LocalMux
    port map (
            O => \N__35588\,
            I => \N__35585\
        );

    \I__8525\ : Span4Mux_h
    port map (
            O => \N__35585\,
            I => \N__35581\
        );

    \I__8524\ : InMux
    port map (
            O => \N__35584\,
            I => \N__35578\
        );

    \I__8523\ : Span4Mux_h
    port map (
            O => \N__35581\,
            I => \N__35572\
        );

    \I__8522\ : LocalMux
    port map (
            O => \N__35578\,
            I => \N__35572\
        );

    \I__8521\ : InMux
    port map (
            O => \N__35577\,
            I => \N__35567\
        );

    \I__8520\ : Span4Mux_h
    port map (
            O => \N__35572\,
            I => \N__35564\
        );

    \I__8519\ : InMux
    port map (
            O => \N__35571\,
            I => \N__35561\
        );

    \I__8518\ : InMux
    port map (
            O => \N__35570\,
            I => \N__35558\
        );

    \I__8517\ : LocalMux
    port map (
            O => \N__35567\,
            I => \b2v_inst.dir_energiaZ0Z_5\
        );

    \I__8516\ : Odrv4
    port map (
            O => \N__35564\,
            I => \b2v_inst.dir_energiaZ0Z_5\
        );

    \I__8515\ : LocalMux
    port map (
            O => \N__35561\,
            I => \b2v_inst.dir_energiaZ0Z_5\
        );

    \I__8514\ : LocalMux
    port map (
            O => \N__35558\,
            I => \b2v_inst.dir_energiaZ0Z_5\
        );

    \I__8513\ : CascadeMux
    port map (
            O => \N__35549\,
            I => \N__35545\
        );

    \I__8512\ : CascadeMux
    port map (
            O => \N__35548\,
            I => \N__35542\
        );

    \I__8511\ : CascadeBuf
    port map (
            O => \N__35545\,
            I => \N__35539\
        );

    \I__8510\ : CascadeBuf
    port map (
            O => \N__35542\,
            I => \N__35536\
        );

    \I__8509\ : CascadeMux
    port map (
            O => \N__35539\,
            I => \N__35533\
        );

    \I__8508\ : CascadeMux
    port map (
            O => \N__35536\,
            I => \N__35530\
        );

    \I__8507\ : CascadeBuf
    port map (
            O => \N__35533\,
            I => \N__35527\
        );

    \I__8506\ : CascadeBuf
    port map (
            O => \N__35530\,
            I => \N__35524\
        );

    \I__8505\ : CascadeMux
    port map (
            O => \N__35527\,
            I => \N__35521\
        );

    \I__8504\ : CascadeMux
    port map (
            O => \N__35524\,
            I => \N__35518\
        );

    \I__8503\ : InMux
    port map (
            O => \N__35521\,
            I => \N__35515\
        );

    \I__8502\ : InMux
    port map (
            O => \N__35518\,
            I => \N__35512\
        );

    \I__8501\ : LocalMux
    port map (
            O => \N__35515\,
            I => \N__35509\
        );

    \I__8500\ : LocalMux
    port map (
            O => \N__35512\,
            I => \N_355_i\
        );

    \I__8499\ : Odrv4
    port map (
            O => \N__35509\,
            I => \N_355_i\
        );

    \I__8498\ : InMux
    port map (
            O => \N__35504\,
            I => \N__35501\
        );

    \I__8497\ : LocalMux
    port map (
            O => \N__35501\,
            I => \N__35497\
        );

    \I__8496\ : InMux
    port map (
            O => \N__35500\,
            I => \N__35494\
        );

    \I__8495\ : Span4Mux_h
    port map (
            O => \N__35497\,
            I => \N__35488\
        );

    \I__8494\ : LocalMux
    port map (
            O => \N__35494\,
            I => \N__35488\
        );

    \I__8493\ : InMux
    port map (
            O => \N__35493\,
            I => \N__35485\
        );

    \I__8492\ : Span4Mux_v
    port map (
            O => \N__35488\,
            I => \N__35479\
        );

    \I__8491\ : LocalMux
    port map (
            O => \N__35485\,
            I => \N__35479\
        );

    \I__8490\ : InMux
    port map (
            O => \N__35484\,
            I => \N__35476\
        );

    \I__8489\ : Span4Mux_h
    port map (
            O => \N__35479\,
            I => \N__35473\
        );

    \I__8488\ : LocalMux
    port map (
            O => \N__35476\,
            I => \N__35470\
        );

    \I__8487\ : Span4Mux_h
    port map (
            O => \N__35473\,
            I => \N__35467\
        );

    \I__8486\ : Odrv12
    port map (
            O => \N__35470\,
            I => b2v_inst_data_a_escribir_7
        );

    \I__8485\ : Odrv4
    port map (
            O => \N__35467\,
            I => b2v_inst_data_a_escribir_7
        );

    \I__8484\ : InMux
    port map (
            O => \N__35462\,
            I => \N__35459\
        );

    \I__8483\ : LocalMux
    port map (
            O => \N__35459\,
            I => \N__35456\
        );

    \I__8482\ : Span4Mux_v
    port map (
            O => \N__35456\,
            I => \N__35453\
        );

    \I__8481\ : Odrv4
    port map (
            O => \N__35453\,
            I => \N_113_i\
        );

    \I__8480\ : InMux
    port map (
            O => \N__35450\,
            I => \N__35447\
        );

    \I__8479\ : LocalMux
    port map (
            O => \N__35447\,
            I => \N__35444\
        );

    \I__8478\ : Span4Mux_h
    port map (
            O => \N__35444\,
            I => \N__35441\
        );

    \I__8477\ : Span4Mux_v
    port map (
            O => \N__35441\,
            I => \N__35438\
        );

    \I__8476\ : Span4Mux_h
    port map (
            O => \N__35438\,
            I => \N__35435\
        );

    \I__8475\ : Odrv4
    port map (
            O => \N__35435\,
            I => \b2v_inst.addr_ram_iv_i_0_0_1\
        );

    \I__8474\ : CascadeMux
    port map (
            O => \N__35432\,
            I => \N__35429\
        );

    \I__8473\ : InMux
    port map (
            O => \N__35429\,
            I => \N__35426\
        );

    \I__8472\ : LocalMux
    port map (
            O => \N__35426\,
            I => \N__35423\
        );

    \I__8471\ : Span4Mux_h
    port map (
            O => \N__35423\,
            I => \N__35420\
        );

    \I__8470\ : Span4Mux_h
    port map (
            O => \N__35420\,
            I => \N__35417\
        );

    \I__8469\ : Span4Mux_v
    port map (
            O => \N__35417\,
            I => \N__35414\
        );

    \I__8468\ : Odrv4
    port map (
            O => \N__35414\,
            I => \b2v_inst.addr_ram_iv_i_0_1_1\
        );

    \I__8467\ : CascadeMux
    port map (
            O => \N__35411\,
            I => \N__35407\
        );

    \I__8466\ : CascadeMux
    port map (
            O => \N__35410\,
            I => \N__35404\
        );

    \I__8465\ : CascadeBuf
    port map (
            O => \N__35407\,
            I => \N__35401\
        );

    \I__8464\ : CascadeBuf
    port map (
            O => \N__35404\,
            I => \N__35398\
        );

    \I__8463\ : CascadeMux
    port map (
            O => \N__35401\,
            I => \N__35395\
        );

    \I__8462\ : CascadeMux
    port map (
            O => \N__35398\,
            I => \N__35392\
        );

    \I__8461\ : CascadeBuf
    port map (
            O => \N__35395\,
            I => \N__35389\
        );

    \I__8460\ : CascadeBuf
    port map (
            O => \N__35392\,
            I => \N__35386\
        );

    \I__8459\ : CascadeMux
    port map (
            O => \N__35389\,
            I => \N__35383\
        );

    \I__8458\ : CascadeMux
    port map (
            O => \N__35386\,
            I => \N__35380\
        );

    \I__8457\ : CascadeBuf
    port map (
            O => \N__35383\,
            I => \N__35377\
        );

    \I__8456\ : CascadeBuf
    port map (
            O => \N__35380\,
            I => \N__35374\
        );

    \I__8455\ : CascadeMux
    port map (
            O => \N__35377\,
            I => \N__35371\
        );

    \I__8454\ : CascadeMux
    port map (
            O => \N__35374\,
            I => \N__35368\
        );

    \I__8453\ : CascadeBuf
    port map (
            O => \N__35371\,
            I => \N__35365\
        );

    \I__8452\ : CascadeBuf
    port map (
            O => \N__35368\,
            I => \N__35362\
        );

    \I__8451\ : CascadeMux
    port map (
            O => \N__35365\,
            I => \N__35359\
        );

    \I__8450\ : CascadeMux
    port map (
            O => \N__35362\,
            I => \N__35356\
        );

    \I__8449\ : CascadeBuf
    port map (
            O => \N__35359\,
            I => \N__35353\
        );

    \I__8448\ : CascadeBuf
    port map (
            O => \N__35356\,
            I => \N__35350\
        );

    \I__8447\ : CascadeMux
    port map (
            O => \N__35353\,
            I => \N__35347\
        );

    \I__8446\ : CascadeMux
    port map (
            O => \N__35350\,
            I => \N__35344\
        );

    \I__8445\ : InMux
    port map (
            O => \N__35347\,
            I => \N__35341\
        );

    \I__8444\ : InMux
    port map (
            O => \N__35344\,
            I => \N__35338\
        );

    \I__8443\ : LocalMux
    port map (
            O => \N__35341\,
            I => \N__35335\
        );

    \I__8442\ : LocalMux
    port map (
            O => \N__35338\,
            I => \indice_RNI8K233_1\
        );

    \I__8441\ : Odrv4
    port map (
            O => \N__35335\,
            I => \indice_RNI8K233_1\
        );

    \I__8440\ : CascadeMux
    port map (
            O => \N__35330\,
            I => \N__35327\
        );

    \I__8439\ : InMux
    port map (
            O => \N__35327\,
            I => \N__35323\
        );

    \I__8438\ : InMux
    port map (
            O => \N__35326\,
            I => \N__35319\
        );

    \I__8437\ : LocalMux
    port map (
            O => \N__35323\,
            I => \N__35316\
        );

    \I__8436\ : CascadeMux
    port map (
            O => \N__35322\,
            I => \N__35312\
        );

    \I__8435\ : LocalMux
    port map (
            O => \N__35319\,
            I => \N__35309\
        );

    \I__8434\ : Span4Mux_v
    port map (
            O => \N__35316\,
            I => \N__35306\
        );

    \I__8433\ : InMux
    port map (
            O => \N__35315\,
            I => \N__35303\
        );

    \I__8432\ : InMux
    port map (
            O => \N__35312\,
            I => \N__35300\
        );

    \I__8431\ : Span4Mux_h
    port map (
            O => \N__35309\,
            I => \N__35297\
        );

    \I__8430\ : Span4Mux_h
    port map (
            O => \N__35306\,
            I => \N__35294\
        );

    \I__8429\ : LocalMux
    port map (
            O => \N__35303\,
            I => \N__35291\
        );

    \I__8428\ : LocalMux
    port map (
            O => \N__35300\,
            I => \N__35288\
        );

    \I__8427\ : Span4Mux_h
    port map (
            O => \N__35297\,
            I => \N__35285\
        );

    \I__8426\ : Span4Mux_h
    port map (
            O => \N__35294\,
            I => \N__35280\
        );

    \I__8425\ : Span4Mux_h
    port map (
            O => \N__35291\,
            I => \N__35280\
        );

    \I__8424\ : Span12Mux_v
    port map (
            O => \N__35288\,
            I => \N__35277\
        );

    \I__8423\ : Odrv4
    port map (
            O => \N__35285\,
            I => b2v_inst_data_a_escribir_6
        );

    \I__8422\ : Odrv4
    port map (
            O => \N__35280\,
            I => b2v_inst_data_a_escribir_6
        );

    \I__8421\ : Odrv12
    port map (
            O => \N__35277\,
            I => b2v_inst_data_a_escribir_6
        );

    \I__8420\ : InMux
    port map (
            O => \N__35270\,
            I => \N__35267\
        );

    \I__8419\ : LocalMux
    port map (
            O => \N__35267\,
            I => \N__35264\
        );

    \I__8418\ : Span4Mux_v
    port map (
            O => \N__35264\,
            I => \N__35261\
        );

    \I__8417\ : Odrv4
    port map (
            O => \N__35261\,
            I => \N_114_i\
        );

    \I__8416\ : InMux
    port map (
            O => \N__35258\,
            I => \N__35255\
        );

    \I__8415\ : LocalMux
    port map (
            O => \N__35255\,
            I => \N__35252\
        );

    \I__8414\ : Span4Mux_v
    port map (
            O => \N__35252\,
            I => \N__35249\
        );

    \I__8413\ : Span4Mux_h
    port map (
            O => \N__35249\,
            I => \N__35246\
        );

    \I__8412\ : Odrv4
    port map (
            O => \N__35246\,
            I => \b2v_inst.addr_ram_iv_i_0_2\
        );

    \I__8411\ : InMux
    port map (
            O => \N__35243\,
            I => \N__35228\
        );

    \I__8410\ : InMux
    port map (
            O => \N__35242\,
            I => \N__35228\
        );

    \I__8409\ : InMux
    port map (
            O => \N__35241\,
            I => \N__35228\
        );

    \I__8408\ : InMux
    port map (
            O => \N__35240\,
            I => \N__35228\
        );

    \I__8407\ : InMux
    port map (
            O => \N__35239\,
            I => \N__35223\
        );

    \I__8406\ : InMux
    port map (
            O => \N__35238\,
            I => \N__35223\
        );

    \I__8405\ : InMux
    port map (
            O => \N__35237\,
            I => \N__35220\
        );

    \I__8404\ : LocalMux
    port map (
            O => \N__35228\,
            I => \N__35210\
        );

    \I__8403\ : LocalMux
    port map (
            O => \N__35223\,
            I => \N__35210\
        );

    \I__8402\ : LocalMux
    port map (
            O => \N__35220\,
            I => \N__35204\
        );

    \I__8401\ : InMux
    port map (
            O => \N__35219\,
            I => \N__35197\
        );

    \I__8400\ : InMux
    port map (
            O => \N__35218\,
            I => \N__35197\
        );

    \I__8399\ : InMux
    port map (
            O => \N__35217\,
            I => \N__35197\
        );

    \I__8398\ : InMux
    port map (
            O => \N__35216\,
            I => \N__35193\
        );

    \I__8397\ : InMux
    port map (
            O => \N__35215\,
            I => \N__35190\
        );

    \I__8396\ : Span4Mux_v
    port map (
            O => \N__35210\,
            I => \N__35182\
        );

    \I__8395\ : InMux
    port map (
            O => \N__35209\,
            I => \N__35179\
        );

    \I__8394\ : InMux
    port map (
            O => \N__35208\,
            I => \N__35176\
        );

    \I__8393\ : InMux
    port map (
            O => \N__35207\,
            I => \N__35173\
        );

    \I__8392\ : Span4Mux_v
    port map (
            O => \N__35204\,
            I => \N__35167\
        );

    \I__8391\ : LocalMux
    port map (
            O => \N__35197\,
            I => \N__35167\
        );

    \I__8390\ : InMux
    port map (
            O => \N__35196\,
            I => \N__35163\
        );

    \I__8389\ : LocalMux
    port map (
            O => \N__35193\,
            I => \N__35160\
        );

    \I__8388\ : LocalMux
    port map (
            O => \N__35190\,
            I => \N__35157\
        );

    \I__8387\ : InMux
    port map (
            O => \N__35189\,
            I => \N__35148\
        );

    \I__8386\ : InMux
    port map (
            O => \N__35188\,
            I => \N__35148\
        );

    \I__8385\ : InMux
    port map (
            O => \N__35187\,
            I => \N__35148\
        );

    \I__8384\ : InMux
    port map (
            O => \N__35186\,
            I => \N__35148\
        );

    \I__8383\ : InMux
    port map (
            O => \N__35185\,
            I => \N__35145\
        );

    \I__8382\ : Sp12to4
    port map (
            O => \N__35182\,
            I => \N__35140\
        );

    \I__8381\ : LocalMux
    port map (
            O => \N__35179\,
            I => \N__35140\
        );

    \I__8380\ : LocalMux
    port map (
            O => \N__35176\,
            I => \N__35137\
        );

    \I__8379\ : LocalMux
    port map (
            O => \N__35173\,
            I => \N__35134\
        );

    \I__8378\ : InMux
    port map (
            O => \N__35172\,
            I => \N__35131\
        );

    \I__8377\ : Span4Mux_v
    port map (
            O => \N__35167\,
            I => \N__35128\
        );

    \I__8376\ : InMux
    port map (
            O => \N__35166\,
            I => \N__35125\
        );

    \I__8375\ : LocalMux
    port map (
            O => \N__35163\,
            I => \N__35122\
        );

    \I__8374\ : Span4Mux_v
    port map (
            O => \N__35160\,
            I => \N__35119\
        );

    \I__8373\ : Span4Mux_v
    port map (
            O => \N__35157\,
            I => \N__35116\
        );

    \I__8372\ : LocalMux
    port map (
            O => \N__35148\,
            I => \N__35113\
        );

    \I__8371\ : LocalMux
    port map (
            O => \N__35145\,
            I => \N__35108\
        );

    \I__8370\ : Span12Mux_h
    port map (
            O => \N__35140\,
            I => \N__35108\
        );

    \I__8369\ : Span12Mux_h
    port map (
            O => \N__35137\,
            I => \N__35105\
        );

    \I__8368\ : Span4Mux_v
    port map (
            O => \N__35134\,
            I => \N__35100\
        );

    \I__8367\ : LocalMux
    port map (
            O => \N__35131\,
            I => \N__35100\
        );

    \I__8366\ : Span4Mux_h
    port map (
            O => \N__35128\,
            I => \N__35095\
        );

    \I__8365\ : LocalMux
    port map (
            O => \N__35125\,
            I => \N__35095\
        );

    \I__8364\ : Span12Mux_h
    port map (
            O => \N__35122\,
            I => \N__35092\
        );

    \I__8363\ : Odrv4
    port map (
            O => \N__35119\,
            I => \b2v_inst.N_480\
        );

    \I__8362\ : Odrv4
    port map (
            O => \N__35116\,
            I => \b2v_inst.N_480\
        );

    \I__8361\ : Odrv4
    port map (
            O => \N__35113\,
            I => \b2v_inst.N_480\
        );

    \I__8360\ : Odrv12
    port map (
            O => \N__35108\,
            I => \b2v_inst.N_480\
        );

    \I__8359\ : Odrv12
    port map (
            O => \N__35105\,
            I => \b2v_inst.N_480\
        );

    \I__8358\ : Odrv4
    port map (
            O => \N__35100\,
            I => \b2v_inst.N_480\
        );

    \I__8357\ : Odrv4
    port map (
            O => \N__35095\,
            I => \b2v_inst.N_480\
        );

    \I__8356\ : Odrv12
    port map (
            O => \N__35092\,
            I => \b2v_inst.N_480\
        );

    \I__8355\ : CascadeMux
    port map (
            O => \N__35075\,
            I => \N__35072\
        );

    \I__8354\ : InMux
    port map (
            O => \N__35072\,
            I => \N__35069\
        );

    \I__8353\ : LocalMux
    port map (
            O => \N__35069\,
            I => \N__35066\
        );

    \I__8352\ : Span4Mux_v
    port map (
            O => \N__35066\,
            I => \N__35063\
        );

    \I__8351\ : Span4Mux_h
    port map (
            O => \N__35063\,
            I => \N__35060\
        );

    \I__8350\ : Odrv4
    port map (
            O => \N__35060\,
            I => \b2v_inst.addr_ram_iv_i_1_2\
        );

    \I__8349\ : CascadeMux
    port map (
            O => \N__35057\,
            I => \N__35053\
        );

    \I__8348\ : CascadeMux
    port map (
            O => \N__35056\,
            I => \N__35050\
        );

    \I__8347\ : CascadeBuf
    port map (
            O => \N__35053\,
            I => \N__35047\
        );

    \I__8346\ : CascadeBuf
    port map (
            O => \N__35050\,
            I => \N__35044\
        );

    \I__8345\ : CascadeMux
    port map (
            O => \N__35047\,
            I => \N__35041\
        );

    \I__8344\ : CascadeMux
    port map (
            O => \N__35044\,
            I => \N__35038\
        );

    \I__8343\ : CascadeBuf
    port map (
            O => \N__35041\,
            I => \N__35035\
        );

    \I__8342\ : CascadeBuf
    port map (
            O => \N__35038\,
            I => \N__35032\
        );

    \I__8341\ : CascadeMux
    port map (
            O => \N__35035\,
            I => \N__35029\
        );

    \I__8340\ : CascadeMux
    port map (
            O => \N__35032\,
            I => \N__35026\
        );

    \I__8339\ : CascadeBuf
    port map (
            O => \N__35029\,
            I => \N__35023\
        );

    \I__8338\ : CascadeBuf
    port map (
            O => \N__35026\,
            I => \N__35020\
        );

    \I__8337\ : CascadeMux
    port map (
            O => \N__35023\,
            I => \N__35017\
        );

    \I__8336\ : CascadeMux
    port map (
            O => \N__35020\,
            I => \N__35014\
        );

    \I__8335\ : CascadeBuf
    port map (
            O => \N__35017\,
            I => \N__35011\
        );

    \I__8334\ : CascadeBuf
    port map (
            O => \N__35014\,
            I => \N__35008\
        );

    \I__8333\ : CascadeMux
    port map (
            O => \N__35011\,
            I => \N__35005\
        );

    \I__8332\ : CascadeMux
    port map (
            O => \N__35008\,
            I => \N__35002\
        );

    \I__8331\ : CascadeBuf
    port map (
            O => \N__35005\,
            I => \N__34999\
        );

    \I__8330\ : CascadeBuf
    port map (
            O => \N__35002\,
            I => \N__34996\
        );

    \I__8329\ : CascadeMux
    port map (
            O => \N__34999\,
            I => \N__34993\
        );

    \I__8328\ : CascadeMux
    port map (
            O => \N__34996\,
            I => \N__34990\
        );

    \I__8327\ : InMux
    port map (
            O => \N__34993\,
            I => \N__34987\
        );

    \I__8326\ : InMux
    port map (
            O => \N__34990\,
            I => \N__34984\
        );

    \I__8325\ : LocalMux
    port map (
            O => \N__34987\,
            I => \N__34979\
        );

    \I__8324\ : LocalMux
    port map (
            O => \N__34984\,
            I => \N__34979\
        );

    \I__8323\ : Odrv4
    port map (
            O => \N__34979\,
            I => \indice_RNIDP233_2\
        );

    \I__8322\ : InMux
    port map (
            O => \N__34976\,
            I => \N__34970\
        );

    \I__8321\ : InMux
    port map (
            O => \N__34975\,
            I => \N__34967\
        );

    \I__8320\ : InMux
    port map (
            O => \N__34974\,
            I => \N__34963\
        );

    \I__8319\ : InMux
    port map (
            O => \N__34973\,
            I => \N__34960\
        );

    \I__8318\ : LocalMux
    port map (
            O => \N__34970\,
            I => \N__34957\
        );

    \I__8317\ : LocalMux
    port map (
            O => \N__34967\,
            I => \N__34954\
        );

    \I__8316\ : CascadeMux
    port map (
            O => \N__34966\,
            I => \N__34951\
        );

    \I__8315\ : LocalMux
    port map (
            O => \N__34963\,
            I => \N__34948\
        );

    \I__8314\ : LocalMux
    port map (
            O => \N__34960\,
            I => \N__34945\
        );

    \I__8313\ : Span4Mux_h
    port map (
            O => \N__34957\,
            I => \N__34942\
        );

    \I__8312\ : Span4Mux_v
    port map (
            O => \N__34954\,
            I => \N__34939\
        );

    \I__8311\ : InMux
    port map (
            O => \N__34951\,
            I => \N__34936\
        );

    \I__8310\ : Span4Mux_v
    port map (
            O => \N__34948\,
            I => \N__34931\
        );

    \I__8309\ : Span4Mux_v
    port map (
            O => \N__34945\,
            I => \N__34931\
        );

    \I__8308\ : Span4Mux_v
    port map (
            O => \N__34942\,
            I => \N__34928\
        );

    \I__8307\ : Sp12to4
    port map (
            O => \N__34939\,
            I => \N__34921\
        );

    \I__8306\ : LocalMux
    port map (
            O => \N__34936\,
            I => \N__34921\
        );

    \I__8305\ : Sp12to4
    port map (
            O => \N__34931\,
            I => \N__34921\
        );

    \I__8304\ : Odrv4
    port map (
            O => \N__34928\,
            I => b2v_inst_data_a_escribir_0
        );

    \I__8303\ : Odrv12
    port map (
            O => \N__34921\,
            I => b2v_inst_data_a_escribir_0
        );

    \I__8302\ : InMux
    port map (
            O => \N__34916\,
            I => \N__34913\
        );

    \I__8301\ : LocalMux
    port map (
            O => \N__34913\,
            I => \N_557_i\
        );

    \I__8300\ : InMux
    port map (
            O => \N__34910\,
            I => \N__34904\
        );

    \I__8299\ : CascadeMux
    port map (
            O => \N__34909\,
            I => \N__34900\
        );

    \I__8298\ : InMux
    port map (
            O => \N__34908\,
            I => \N__34897\
        );

    \I__8297\ : InMux
    port map (
            O => \N__34907\,
            I => \N__34894\
        );

    \I__8296\ : LocalMux
    port map (
            O => \N__34904\,
            I => \N__34891\
        );

    \I__8295\ : InMux
    port map (
            O => \N__34903\,
            I => \N__34888\
        );

    \I__8294\ : InMux
    port map (
            O => \N__34900\,
            I => \N__34885\
        );

    \I__8293\ : LocalMux
    port map (
            O => \N__34897\,
            I => b2v_inst_cantidad_temp_0
        );

    \I__8292\ : LocalMux
    port map (
            O => \N__34894\,
            I => b2v_inst_cantidad_temp_0
        );

    \I__8291\ : Odrv12
    port map (
            O => \N__34891\,
            I => b2v_inst_cantidad_temp_0
        );

    \I__8290\ : LocalMux
    port map (
            O => \N__34888\,
            I => b2v_inst_cantidad_temp_0
        );

    \I__8289\ : LocalMux
    port map (
            O => \N__34885\,
            I => b2v_inst_cantidad_temp_0
        );

    \I__8288\ : InMux
    port map (
            O => \N__34874\,
            I => \N__34871\
        );

    \I__8287\ : LocalMux
    port map (
            O => \N__34871\,
            I => \N__34867\
        );

    \I__8286\ : InMux
    port map (
            O => \N__34870\,
            I => \N__34862\
        );

    \I__8285\ : Span4Mux_h
    port map (
            O => \N__34867\,
            I => \N__34859\
        );

    \I__8284\ : InMux
    port map (
            O => \N__34866\,
            I => \N__34856\
        );

    \I__8283\ : InMux
    port map (
            O => \N__34865\,
            I => \N__34853\
        );

    \I__8282\ : LocalMux
    port map (
            O => \N__34862\,
            I => b2v_inst_cantidad_temp_1
        );

    \I__8281\ : Odrv4
    port map (
            O => \N__34859\,
            I => b2v_inst_cantidad_temp_1
        );

    \I__8280\ : LocalMux
    port map (
            O => \N__34856\,
            I => b2v_inst_cantidad_temp_1
        );

    \I__8279\ : LocalMux
    port map (
            O => \N__34853\,
            I => b2v_inst_cantidad_temp_1
        );

    \I__8278\ : CascadeMux
    port map (
            O => \N__34844\,
            I => \N__34841\
        );

    \I__8277\ : InMux
    port map (
            O => \N__34841\,
            I => \N__34835\
        );

    \I__8276\ : InMux
    port map (
            O => \N__34840\,
            I => \N__34832\
        );

    \I__8275\ : CascadeMux
    port map (
            O => \N__34839\,
            I => \N__34829\
        );

    \I__8274\ : InMux
    port map (
            O => \N__34838\,
            I => \N__34826\
        );

    \I__8273\ : LocalMux
    port map (
            O => \N__34835\,
            I => \N__34822\
        );

    \I__8272\ : LocalMux
    port map (
            O => \N__34832\,
            I => \N__34819\
        );

    \I__8271\ : InMux
    port map (
            O => \N__34829\,
            I => \N__34816\
        );

    \I__8270\ : LocalMux
    port map (
            O => \N__34826\,
            I => \N__34813\
        );

    \I__8269\ : InMux
    port map (
            O => \N__34825\,
            I => \N__34810\
        );

    \I__8268\ : Span4Mux_h
    port map (
            O => \N__34822\,
            I => \N__34807\
        );

    \I__8267\ : Span4Mux_v
    port map (
            O => \N__34819\,
            I => \N__34804\
        );

    \I__8266\ : LocalMux
    port map (
            O => \N__34816\,
            I => \N__34801\
        );

    \I__8265\ : Span4Mux_v
    port map (
            O => \N__34813\,
            I => \N__34798\
        );

    \I__8264\ : LocalMux
    port map (
            O => \N__34810\,
            I => \N__34795\
        );

    \I__8263\ : Span4Mux_v
    port map (
            O => \N__34807\,
            I => \N__34792\
        );

    \I__8262\ : Span4Mux_h
    port map (
            O => \N__34804\,
            I => \N__34787\
        );

    \I__8261\ : Span4Mux_h
    port map (
            O => \N__34801\,
            I => \N__34787\
        );

    \I__8260\ : Span4Mux_h
    port map (
            O => \N__34798\,
            I => \N__34782\
        );

    \I__8259\ : Span4Mux_h
    port map (
            O => \N__34795\,
            I => \N__34782\
        );

    \I__8258\ : Odrv4
    port map (
            O => \N__34792\,
            I => b2v_inst_data_a_escribir_1
        );

    \I__8257\ : Odrv4
    port map (
            O => \N__34787\,
            I => b2v_inst_data_a_escribir_1
        );

    \I__8256\ : Odrv4
    port map (
            O => \N__34782\,
            I => b2v_inst_data_a_escribir_1
        );

    \I__8255\ : CascadeMux
    port map (
            O => \N__34775\,
            I => \b2v_inst.cantidad_temp_RNILL3KZ0Z_1_cascade_\
        );

    \I__8254\ : InMux
    port map (
            O => \N__34772\,
            I => \N__34769\
        );

    \I__8253\ : LocalMux
    port map (
            O => \N__34769\,
            I => \N_555_i\
        );

    \I__8252\ : InMux
    port map (
            O => \N__34766\,
            I => \N__34758\
        );

    \I__8251\ : InMux
    port map (
            O => \N__34765\,
            I => \N__34755\
        );

    \I__8250\ : InMux
    port map (
            O => \N__34764\,
            I => \N__34752\
        );

    \I__8249\ : InMux
    port map (
            O => \N__34763\,
            I => \N__34747\
        );

    \I__8248\ : InMux
    port map (
            O => \N__34762\,
            I => \N__34747\
        );

    \I__8247\ : InMux
    port map (
            O => \N__34761\,
            I => \N__34742\
        );

    \I__8246\ : LocalMux
    port map (
            O => \N__34758\,
            I => \N__34738\
        );

    \I__8245\ : LocalMux
    port map (
            O => \N__34755\,
            I => \N__34731\
        );

    \I__8244\ : LocalMux
    port map (
            O => \N__34752\,
            I => \N__34731\
        );

    \I__8243\ : LocalMux
    port map (
            O => \N__34747\,
            I => \N__34731\
        );

    \I__8242\ : CascadeMux
    port map (
            O => \N__34746\,
            I => \N__34728\
        );

    \I__8241\ : InMux
    port map (
            O => \N__34745\,
            I => \N__34722\
        );

    \I__8240\ : LocalMux
    port map (
            O => \N__34742\,
            I => \N__34719\
        );

    \I__8239\ : InMux
    port map (
            O => \N__34741\,
            I => \N__34716\
        );

    \I__8238\ : Span4Mux_v
    port map (
            O => \N__34738\,
            I => \N__34713\
        );

    \I__8237\ : Span4Mux_v
    port map (
            O => \N__34731\,
            I => \N__34710\
        );

    \I__8236\ : InMux
    port map (
            O => \N__34728\,
            I => \N__34707\
        );

    \I__8235\ : CascadeMux
    port map (
            O => \N__34727\,
            I => \N__34703\
        );

    \I__8234\ : InMux
    port map (
            O => \N__34726\,
            I => \N__34698\
        );

    \I__8233\ : InMux
    port map (
            O => \N__34725\,
            I => \N__34698\
        );

    \I__8232\ : LocalMux
    port map (
            O => \N__34722\,
            I => \N__34695\
        );

    \I__8231\ : Span4Mux_h
    port map (
            O => \N__34719\,
            I => \N__34691\
        );

    \I__8230\ : LocalMux
    port map (
            O => \N__34716\,
            I => \N__34688\
        );

    \I__8229\ : Sp12to4
    port map (
            O => \N__34713\,
            I => \N__34681\
        );

    \I__8228\ : Sp12to4
    port map (
            O => \N__34710\,
            I => \N__34681\
        );

    \I__8227\ : LocalMux
    port map (
            O => \N__34707\,
            I => \N__34681\
        );

    \I__8226\ : InMux
    port map (
            O => \N__34706\,
            I => \N__34676\
        );

    \I__8225\ : InMux
    port map (
            O => \N__34703\,
            I => \N__34676\
        );

    \I__8224\ : LocalMux
    port map (
            O => \N__34698\,
            I => \N__34673\
        );

    \I__8223\ : Span4Mux_h
    port map (
            O => \N__34695\,
            I => \N__34670\
        );

    \I__8222\ : InMux
    port map (
            O => \N__34694\,
            I => \N__34667\
        );

    \I__8221\ : Odrv4
    port map (
            O => \N__34691\,
            I => \b2v_inst.stateZ0Z_18\
        );

    \I__8220\ : Odrv12
    port map (
            O => \N__34688\,
            I => \b2v_inst.stateZ0Z_18\
        );

    \I__8219\ : Odrv12
    port map (
            O => \N__34681\,
            I => \b2v_inst.stateZ0Z_18\
        );

    \I__8218\ : LocalMux
    port map (
            O => \N__34676\,
            I => \b2v_inst.stateZ0Z_18\
        );

    \I__8217\ : Odrv4
    port map (
            O => \N__34673\,
            I => \b2v_inst.stateZ0Z_18\
        );

    \I__8216\ : Odrv4
    port map (
            O => \N__34670\,
            I => \b2v_inst.stateZ0Z_18\
        );

    \I__8215\ : LocalMux
    port map (
            O => \N__34667\,
            I => \b2v_inst.stateZ0Z_18\
        );

    \I__8214\ : CascadeMux
    port map (
            O => \N__34652\,
            I => \N__34649\
        );

    \I__8213\ : InMux
    port map (
            O => \N__34649\,
            I => \N__34646\
        );

    \I__8212\ : LocalMux
    port map (
            O => \N__34646\,
            I => \SYNTHESIZED_WIRE_1_3\
        );

    \I__8211\ : InMux
    port map (
            O => \N__34643\,
            I => \N__34639\
        );

    \I__8210\ : InMux
    port map (
            O => \N__34642\,
            I => \N__34636\
        );

    \I__8209\ : LocalMux
    port map (
            O => \N__34639\,
            I => \N__34633\
        );

    \I__8208\ : LocalMux
    port map (
            O => \N__34636\,
            I => \N__34630\
        );

    \I__8207\ : Span4Mux_v
    port map (
            O => \N__34633\,
            I => \N__34620\
        );

    \I__8206\ : Span4Mux_v
    port map (
            O => \N__34630\,
            I => \N__34617\
        );

    \I__8205\ : InMux
    port map (
            O => \N__34629\,
            I => \N__34610\
        );

    \I__8204\ : InMux
    port map (
            O => \N__34628\,
            I => \N__34610\
        );

    \I__8203\ : InMux
    port map (
            O => \N__34627\,
            I => \N__34610\
        );

    \I__8202\ : InMux
    port map (
            O => \N__34626\,
            I => \N__34607\
        );

    \I__8201\ : InMux
    port map (
            O => \N__34625\,
            I => \N__34604\
        );

    \I__8200\ : InMux
    port map (
            O => \N__34624\,
            I => \N__34599\
        );

    \I__8199\ : InMux
    port map (
            O => \N__34623\,
            I => \N__34599\
        );

    \I__8198\ : Sp12to4
    port map (
            O => \N__34620\,
            I => \N__34592\
        );

    \I__8197\ : Sp12to4
    port map (
            O => \N__34617\,
            I => \N__34592\
        );

    \I__8196\ : LocalMux
    port map (
            O => \N__34610\,
            I => \N__34592\
        );

    \I__8195\ : LocalMux
    port map (
            O => \N__34607\,
            I => \N__34589\
        );

    \I__8194\ : LocalMux
    port map (
            O => \N__34604\,
            I => \N__34583\
        );

    \I__8193\ : LocalMux
    port map (
            O => \N__34599\,
            I => \N__34583\
        );

    \I__8192\ : Span12Mux_h
    port map (
            O => \N__34592\,
            I => \N__34579\
        );

    \I__8191\ : Span4Mux_h
    port map (
            O => \N__34589\,
            I => \N__34576\
        );

    \I__8190\ : InMux
    port map (
            O => \N__34588\,
            I => \N__34573\
        );

    \I__8189\ : Span4Mux_h
    port map (
            O => \N__34583\,
            I => \N__34570\
        );

    \I__8188\ : InMux
    port map (
            O => \N__34582\,
            I => \N__34567\
        );

    \I__8187\ : Odrv12
    port map (
            O => \N__34579\,
            I => \b2v_inst.stateZ0Z_9\
        );

    \I__8186\ : Odrv4
    port map (
            O => \N__34576\,
            I => \b2v_inst.stateZ0Z_9\
        );

    \I__8185\ : LocalMux
    port map (
            O => \N__34573\,
            I => \b2v_inst.stateZ0Z_9\
        );

    \I__8184\ : Odrv4
    port map (
            O => \N__34570\,
            I => \b2v_inst.stateZ0Z_9\
        );

    \I__8183\ : LocalMux
    port map (
            O => \N__34567\,
            I => \b2v_inst.stateZ0Z_9\
        );

    \I__8182\ : InMux
    port map (
            O => \N__34556\,
            I => \N__34553\
        );

    \I__8181\ : LocalMux
    port map (
            O => \N__34553\,
            I => \N__34550\
        );

    \I__8180\ : Span4Mux_h
    port map (
            O => \N__34550\,
            I => \N__34546\
        );

    \I__8179\ : InMux
    port map (
            O => \N__34549\,
            I => \N__34542\
        );

    \I__8178\ : Span4Mux_h
    port map (
            O => \N__34546\,
            I => \N__34539\
        );

    \I__8177\ : InMux
    port map (
            O => \N__34545\,
            I => \N__34536\
        );

    \I__8176\ : LocalMux
    port map (
            O => \N__34542\,
            I => b2v_inst_cantidad_temp_3
        );

    \I__8175\ : Odrv4
    port map (
            O => \N__34539\,
            I => b2v_inst_cantidad_temp_3
        );

    \I__8174\ : LocalMux
    port map (
            O => \N__34536\,
            I => b2v_inst_cantidad_temp_3
        );

    \I__8173\ : ClkMux
    port map (
            O => \N__34529\,
            I => \N__34052\
        );

    \I__8172\ : ClkMux
    port map (
            O => \N__34528\,
            I => \N__34052\
        );

    \I__8171\ : ClkMux
    port map (
            O => \N__34527\,
            I => \N__34052\
        );

    \I__8170\ : ClkMux
    port map (
            O => \N__34526\,
            I => \N__34052\
        );

    \I__8169\ : ClkMux
    port map (
            O => \N__34525\,
            I => \N__34052\
        );

    \I__8168\ : ClkMux
    port map (
            O => \N__34524\,
            I => \N__34052\
        );

    \I__8167\ : ClkMux
    port map (
            O => \N__34523\,
            I => \N__34052\
        );

    \I__8166\ : ClkMux
    port map (
            O => \N__34522\,
            I => \N__34052\
        );

    \I__8165\ : ClkMux
    port map (
            O => \N__34521\,
            I => \N__34052\
        );

    \I__8164\ : ClkMux
    port map (
            O => \N__34520\,
            I => \N__34052\
        );

    \I__8163\ : ClkMux
    port map (
            O => \N__34519\,
            I => \N__34052\
        );

    \I__8162\ : ClkMux
    port map (
            O => \N__34518\,
            I => \N__34052\
        );

    \I__8161\ : ClkMux
    port map (
            O => \N__34517\,
            I => \N__34052\
        );

    \I__8160\ : ClkMux
    port map (
            O => \N__34516\,
            I => \N__34052\
        );

    \I__8159\ : ClkMux
    port map (
            O => \N__34515\,
            I => \N__34052\
        );

    \I__8158\ : ClkMux
    port map (
            O => \N__34514\,
            I => \N__34052\
        );

    \I__8157\ : ClkMux
    port map (
            O => \N__34513\,
            I => \N__34052\
        );

    \I__8156\ : ClkMux
    port map (
            O => \N__34512\,
            I => \N__34052\
        );

    \I__8155\ : ClkMux
    port map (
            O => \N__34511\,
            I => \N__34052\
        );

    \I__8154\ : ClkMux
    port map (
            O => \N__34510\,
            I => \N__34052\
        );

    \I__8153\ : ClkMux
    port map (
            O => \N__34509\,
            I => \N__34052\
        );

    \I__8152\ : ClkMux
    port map (
            O => \N__34508\,
            I => \N__34052\
        );

    \I__8151\ : ClkMux
    port map (
            O => \N__34507\,
            I => \N__34052\
        );

    \I__8150\ : ClkMux
    port map (
            O => \N__34506\,
            I => \N__34052\
        );

    \I__8149\ : ClkMux
    port map (
            O => \N__34505\,
            I => \N__34052\
        );

    \I__8148\ : ClkMux
    port map (
            O => \N__34504\,
            I => \N__34052\
        );

    \I__8147\ : ClkMux
    port map (
            O => \N__34503\,
            I => \N__34052\
        );

    \I__8146\ : ClkMux
    port map (
            O => \N__34502\,
            I => \N__34052\
        );

    \I__8145\ : ClkMux
    port map (
            O => \N__34501\,
            I => \N__34052\
        );

    \I__8144\ : ClkMux
    port map (
            O => \N__34500\,
            I => \N__34052\
        );

    \I__8143\ : ClkMux
    port map (
            O => \N__34499\,
            I => \N__34052\
        );

    \I__8142\ : ClkMux
    port map (
            O => \N__34498\,
            I => \N__34052\
        );

    \I__8141\ : ClkMux
    port map (
            O => \N__34497\,
            I => \N__34052\
        );

    \I__8140\ : ClkMux
    port map (
            O => \N__34496\,
            I => \N__34052\
        );

    \I__8139\ : ClkMux
    port map (
            O => \N__34495\,
            I => \N__34052\
        );

    \I__8138\ : ClkMux
    port map (
            O => \N__34494\,
            I => \N__34052\
        );

    \I__8137\ : ClkMux
    port map (
            O => \N__34493\,
            I => \N__34052\
        );

    \I__8136\ : ClkMux
    port map (
            O => \N__34492\,
            I => \N__34052\
        );

    \I__8135\ : ClkMux
    port map (
            O => \N__34491\,
            I => \N__34052\
        );

    \I__8134\ : ClkMux
    port map (
            O => \N__34490\,
            I => \N__34052\
        );

    \I__8133\ : ClkMux
    port map (
            O => \N__34489\,
            I => \N__34052\
        );

    \I__8132\ : ClkMux
    port map (
            O => \N__34488\,
            I => \N__34052\
        );

    \I__8131\ : ClkMux
    port map (
            O => \N__34487\,
            I => \N__34052\
        );

    \I__8130\ : ClkMux
    port map (
            O => \N__34486\,
            I => \N__34052\
        );

    \I__8129\ : ClkMux
    port map (
            O => \N__34485\,
            I => \N__34052\
        );

    \I__8128\ : ClkMux
    port map (
            O => \N__34484\,
            I => \N__34052\
        );

    \I__8127\ : ClkMux
    port map (
            O => \N__34483\,
            I => \N__34052\
        );

    \I__8126\ : ClkMux
    port map (
            O => \N__34482\,
            I => \N__34052\
        );

    \I__8125\ : ClkMux
    port map (
            O => \N__34481\,
            I => \N__34052\
        );

    \I__8124\ : ClkMux
    port map (
            O => \N__34480\,
            I => \N__34052\
        );

    \I__8123\ : ClkMux
    port map (
            O => \N__34479\,
            I => \N__34052\
        );

    \I__8122\ : ClkMux
    port map (
            O => \N__34478\,
            I => \N__34052\
        );

    \I__8121\ : ClkMux
    port map (
            O => \N__34477\,
            I => \N__34052\
        );

    \I__8120\ : ClkMux
    port map (
            O => \N__34476\,
            I => \N__34052\
        );

    \I__8119\ : ClkMux
    port map (
            O => \N__34475\,
            I => \N__34052\
        );

    \I__8118\ : ClkMux
    port map (
            O => \N__34474\,
            I => \N__34052\
        );

    \I__8117\ : ClkMux
    port map (
            O => \N__34473\,
            I => \N__34052\
        );

    \I__8116\ : ClkMux
    port map (
            O => \N__34472\,
            I => \N__34052\
        );

    \I__8115\ : ClkMux
    port map (
            O => \N__34471\,
            I => \N__34052\
        );

    \I__8114\ : ClkMux
    port map (
            O => \N__34470\,
            I => \N__34052\
        );

    \I__8113\ : ClkMux
    port map (
            O => \N__34469\,
            I => \N__34052\
        );

    \I__8112\ : ClkMux
    port map (
            O => \N__34468\,
            I => \N__34052\
        );

    \I__8111\ : ClkMux
    port map (
            O => \N__34467\,
            I => \N__34052\
        );

    \I__8110\ : ClkMux
    port map (
            O => \N__34466\,
            I => \N__34052\
        );

    \I__8109\ : ClkMux
    port map (
            O => \N__34465\,
            I => \N__34052\
        );

    \I__8108\ : ClkMux
    port map (
            O => \N__34464\,
            I => \N__34052\
        );

    \I__8107\ : ClkMux
    port map (
            O => \N__34463\,
            I => \N__34052\
        );

    \I__8106\ : ClkMux
    port map (
            O => \N__34462\,
            I => \N__34052\
        );

    \I__8105\ : ClkMux
    port map (
            O => \N__34461\,
            I => \N__34052\
        );

    \I__8104\ : ClkMux
    port map (
            O => \N__34460\,
            I => \N__34052\
        );

    \I__8103\ : ClkMux
    port map (
            O => \N__34459\,
            I => \N__34052\
        );

    \I__8102\ : ClkMux
    port map (
            O => \N__34458\,
            I => \N__34052\
        );

    \I__8101\ : ClkMux
    port map (
            O => \N__34457\,
            I => \N__34052\
        );

    \I__8100\ : ClkMux
    port map (
            O => \N__34456\,
            I => \N__34052\
        );

    \I__8099\ : ClkMux
    port map (
            O => \N__34455\,
            I => \N__34052\
        );

    \I__8098\ : ClkMux
    port map (
            O => \N__34454\,
            I => \N__34052\
        );

    \I__8097\ : ClkMux
    port map (
            O => \N__34453\,
            I => \N__34052\
        );

    \I__8096\ : ClkMux
    port map (
            O => \N__34452\,
            I => \N__34052\
        );

    \I__8095\ : ClkMux
    port map (
            O => \N__34451\,
            I => \N__34052\
        );

    \I__8094\ : ClkMux
    port map (
            O => \N__34450\,
            I => \N__34052\
        );

    \I__8093\ : ClkMux
    port map (
            O => \N__34449\,
            I => \N__34052\
        );

    \I__8092\ : ClkMux
    port map (
            O => \N__34448\,
            I => \N__34052\
        );

    \I__8091\ : ClkMux
    port map (
            O => \N__34447\,
            I => \N__34052\
        );

    \I__8090\ : ClkMux
    port map (
            O => \N__34446\,
            I => \N__34052\
        );

    \I__8089\ : ClkMux
    port map (
            O => \N__34445\,
            I => \N__34052\
        );

    \I__8088\ : ClkMux
    port map (
            O => \N__34444\,
            I => \N__34052\
        );

    \I__8087\ : ClkMux
    port map (
            O => \N__34443\,
            I => \N__34052\
        );

    \I__8086\ : ClkMux
    port map (
            O => \N__34442\,
            I => \N__34052\
        );

    \I__8085\ : ClkMux
    port map (
            O => \N__34441\,
            I => \N__34052\
        );

    \I__8084\ : ClkMux
    port map (
            O => \N__34440\,
            I => \N__34052\
        );

    \I__8083\ : ClkMux
    port map (
            O => \N__34439\,
            I => \N__34052\
        );

    \I__8082\ : ClkMux
    port map (
            O => \N__34438\,
            I => \N__34052\
        );

    \I__8081\ : ClkMux
    port map (
            O => \N__34437\,
            I => \N__34052\
        );

    \I__8080\ : ClkMux
    port map (
            O => \N__34436\,
            I => \N__34052\
        );

    \I__8079\ : ClkMux
    port map (
            O => \N__34435\,
            I => \N__34052\
        );

    \I__8078\ : ClkMux
    port map (
            O => \N__34434\,
            I => \N__34052\
        );

    \I__8077\ : ClkMux
    port map (
            O => \N__34433\,
            I => \N__34052\
        );

    \I__8076\ : ClkMux
    port map (
            O => \N__34432\,
            I => \N__34052\
        );

    \I__8075\ : ClkMux
    port map (
            O => \N__34431\,
            I => \N__34052\
        );

    \I__8074\ : ClkMux
    port map (
            O => \N__34430\,
            I => \N__34052\
        );

    \I__8073\ : ClkMux
    port map (
            O => \N__34429\,
            I => \N__34052\
        );

    \I__8072\ : ClkMux
    port map (
            O => \N__34428\,
            I => \N__34052\
        );

    \I__8071\ : ClkMux
    port map (
            O => \N__34427\,
            I => \N__34052\
        );

    \I__8070\ : ClkMux
    port map (
            O => \N__34426\,
            I => \N__34052\
        );

    \I__8069\ : ClkMux
    port map (
            O => \N__34425\,
            I => \N__34052\
        );

    \I__8068\ : ClkMux
    port map (
            O => \N__34424\,
            I => \N__34052\
        );

    \I__8067\ : ClkMux
    port map (
            O => \N__34423\,
            I => \N__34052\
        );

    \I__8066\ : ClkMux
    port map (
            O => \N__34422\,
            I => \N__34052\
        );

    \I__8065\ : ClkMux
    port map (
            O => \N__34421\,
            I => \N__34052\
        );

    \I__8064\ : ClkMux
    port map (
            O => \N__34420\,
            I => \N__34052\
        );

    \I__8063\ : ClkMux
    port map (
            O => \N__34419\,
            I => \N__34052\
        );

    \I__8062\ : ClkMux
    port map (
            O => \N__34418\,
            I => \N__34052\
        );

    \I__8061\ : ClkMux
    port map (
            O => \N__34417\,
            I => \N__34052\
        );

    \I__8060\ : ClkMux
    port map (
            O => \N__34416\,
            I => \N__34052\
        );

    \I__8059\ : ClkMux
    port map (
            O => \N__34415\,
            I => \N__34052\
        );

    \I__8058\ : ClkMux
    port map (
            O => \N__34414\,
            I => \N__34052\
        );

    \I__8057\ : ClkMux
    port map (
            O => \N__34413\,
            I => \N__34052\
        );

    \I__8056\ : ClkMux
    port map (
            O => \N__34412\,
            I => \N__34052\
        );

    \I__8055\ : ClkMux
    port map (
            O => \N__34411\,
            I => \N__34052\
        );

    \I__8054\ : ClkMux
    port map (
            O => \N__34410\,
            I => \N__34052\
        );

    \I__8053\ : ClkMux
    port map (
            O => \N__34409\,
            I => \N__34052\
        );

    \I__8052\ : ClkMux
    port map (
            O => \N__34408\,
            I => \N__34052\
        );

    \I__8051\ : ClkMux
    port map (
            O => \N__34407\,
            I => \N__34052\
        );

    \I__8050\ : ClkMux
    port map (
            O => \N__34406\,
            I => \N__34052\
        );

    \I__8049\ : ClkMux
    port map (
            O => \N__34405\,
            I => \N__34052\
        );

    \I__8048\ : ClkMux
    port map (
            O => \N__34404\,
            I => \N__34052\
        );

    \I__8047\ : ClkMux
    port map (
            O => \N__34403\,
            I => \N__34052\
        );

    \I__8046\ : ClkMux
    port map (
            O => \N__34402\,
            I => \N__34052\
        );

    \I__8045\ : ClkMux
    port map (
            O => \N__34401\,
            I => \N__34052\
        );

    \I__8044\ : ClkMux
    port map (
            O => \N__34400\,
            I => \N__34052\
        );

    \I__8043\ : ClkMux
    port map (
            O => \N__34399\,
            I => \N__34052\
        );

    \I__8042\ : ClkMux
    port map (
            O => \N__34398\,
            I => \N__34052\
        );

    \I__8041\ : ClkMux
    port map (
            O => \N__34397\,
            I => \N__34052\
        );

    \I__8040\ : ClkMux
    port map (
            O => \N__34396\,
            I => \N__34052\
        );

    \I__8039\ : ClkMux
    port map (
            O => \N__34395\,
            I => \N__34052\
        );

    \I__8038\ : ClkMux
    port map (
            O => \N__34394\,
            I => \N__34052\
        );

    \I__8037\ : ClkMux
    port map (
            O => \N__34393\,
            I => \N__34052\
        );

    \I__8036\ : ClkMux
    port map (
            O => \N__34392\,
            I => \N__34052\
        );

    \I__8035\ : ClkMux
    port map (
            O => \N__34391\,
            I => \N__34052\
        );

    \I__8034\ : ClkMux
    port map (
            O => \N__34390\,
            I => \N__34052\
        );

    \I__8033\ : ClkMux
    port map (
            O => \N__34389\,
            I => \N__34052\
        );

    \I__8032\ : ClkMux
    port map (
            O => \N__34388\,
            I => \N__34052\
        );

    \I__8031\ : ClkMux
    port map (
            O => \N__34387\,
            I => \N__34052\
        );

    \I__8030\ : ClkMux
    port map (
            O => \N__34386\,
            I => \N__34052\
        );

    \I__8029\ : ClkMux
    port map (
            O => \N__34385\,
            I => \N__34052\
        );

    \I__8028\ : ClkMux
    port map (
            O => \N__34384\,
            I => \N__34052\
        );

    \I__8027\ : ClkMux
    port map (
            O => \N__34383\,
            I => \N__34052\
        );

    \I__8026\ : ClkMux
    port map (
            O => \N__34382\,
            I => \N__34052\
        );

    \I__8025\ : ClkMux
    port map (
            O => \N__34381\,
            I => \N__34052\
        );

    \I__8024\ : ClkMux
    port map (
            O => \N__34380\,
            I => \N__34052\
        );

    \I__8023\ : ClkMux
    port map (
            O => \N__34379\,
            I => \N__34052\
        );

    \I__8022\ : ClkMux
    port map (
            O => \N__34378\,
            I => \N__34052\
        );

    \I__8021\ : ClkMux
    port map (
            O => \N__34377\,
            I => \N__34052\
        );

    \I__8020\ : ClkMux
    port map (
            O => \N__34376\,
            I => \N__34052\
        );

    \I__8019\ : ClkMux
    port map (
            O => \N__34375\,
            I => \N__34052\
        );

    \I__8018\ : ClkMux
    port map (
            O => \N__34374\,
            I => \N__34052\
        );

    \I__8017\ : ClkMux
    port map (
            O => \N__34373\,
            I => \N__34052\
        );

    \I__8016\ : ClkMux
    port map (
            O => \N__34372\,
            I => \N__34052\
        );

    \I__8015\ : ClkMux
    port map (
            O => \N__34371\,
            I => \N__34052\
        );

    \I__8014\ : GlobalMux
    port map (
            O => \N__34052\,
            I => \N__34049\
        );

    \I__8013\ : gio2CtrlBuf
    port map (
            O => \N__34049\,
            I => clk_c_g
        );

    \I__8012\ : InMux
    port map (
            O => \N__34046\,
            I => \N__34043\
        );

    \I__8011\ : LocalMux
    port map (
            O => \N__34043\,
            I => \N__34040\
        );

    \I__8010\ : Span4Mux_h
    port map (
            O => \N__34040\,
            I => \N__34037\
        );

    \I__8009\ : Span4Mux_h
    port map (
            O => \N__34037\,
            I => \N__34034\
        );

    \I__8008\ : Odrv4
    port map (
            O => \N__34034\,
            I => \b2v_inst.addr_ram_iv_i_0_5\
        );

    \I__8007\ : CascadeMux
    port map (
            O => \N__34031\,
            I => \N__34028\
        );

    \I__8006\ : InMux
    port map (
            O => \N__34028\,
            I => \N__34025\
        );

    \I__8005\ : LocalMux
    port map (
            O => \N__34025\,
            I => \N__34022\
        );

    \I__8004\ : Span4Mux_v
    port map (
            O => \N__34022\,
            I => \N__34019\
        );

    \I__8003\ : Span4Mux_h
    port map (
            O => \N__34019\,
            I => \N__34016\
        );

    \I__8002\ : Span4Mux_h
    port map (
            O => \N__34016\,
            I => \N__34013\
        );

    \I__8001\ : Odrv4
    port map (
            O => \N__34013\,
            I => \b2v_inst.addr_ram_iv_i_1_5\
        );

    \I__8000\ : CascadeMux
    port map (
            O => \N__34010\,
            I => \N__34006\
        );

    \I__7999\ : CascadeMux
    port map (
            O => \N__34009\,
            I => \N__34003\
        );

    \I__7998\ : CascadeBuf
    port map (
            O => \N__34006\,
            I => \N__34000\
        );

    \I__7997\ : CascadeBuf
    port map (
            O => \N__34003\,
            I => \N__33997\
        );

    \I__7996\ : CascadeMux
    port map (
            O => \N__34000\,
            I => \N__33994\
        );

    \I__7995\ : CascadeMux
    port map (
            O => \N__33997\,
            I => \N__33991\
        );

    \I__7994\ : CascadeBuf
    port map (
            O => \N__33994\,
            I => \N__33988\
        );

    \I__7993\ : CascadeBuf
    port map (
            O => \N__33991\,
            I => \N__33985\
        );

    \I__7992\ : CascadeMux
    port map (
            O => \N__33988\,
            I => \N__33982\
        );

    \I__7991\ : CascadeMux
    port map (
            O => \N__33985\,
            I => \N__33979\
        );

    \I__7990\ : CascadeBuf
    port map (
            O => \N__33982\,
            I => \N__33976\
        );

    \I__7989\ : CascadeBuf
    port map (
            O => \N__33979\,
            I => \N__33973\
        );

    \I__7988\ : CascadeMux
    port map (
            O => \N__33976\,
            I => \N__33970\
        );

    \I__7987\ : CascadeMux
    port map (
            O => \N__33973\,
            I => \N__33967\
        );

    \I__7986\ : CascadeBuf
    port map (
            O => \N__33970\,
            I => \N__33964\
        );

    \I__7985\ : CascadeBuf
    port map (
            O => \N__33967\,
            I => \N__33961\
        );

    \I__7984\ : CascadeMux
    port map (
            O => \N__33964\,
            I => \N__33958\
        );

    \I__7983\ : CascadeMux
    port map (
            O => \N__33961\,
            I => \N__33955\
        );

    \I__7982\ : CascadeBuf
    port map (
            O => \N__33958\,
            I => \N__33952\
        );

    \I__7981\ : CascadeBuf
    port map (
            O => \N__33955\,
            I => \N__33949\
        );

    \I__7980\ : CascadeMux
    port map (
            O => \N__33952\,
            I => \N__33946\
        );

    \I__7979\ : CascadeMux
    port map (
            O => \N__33949\,
            I => \N__33943\
        );

    \I__7978\ : InMux
    port map (
            O => \N__33946\,
            I => \N__33940\
        );

    \I__7977\ : InMux
    port map (
            O => \N__33943\,
            I => \N__33937\
        );

    \I__7976\ : LocalMux
    port map (
            O => \N__33940\,
            I => \N__33934\
        );

    \I__7975\ : LocalMux
    port map (
            O => \N__33937\,
            I => \indice_RNIS8333_5\
        );

    \I__7974\ : Odrv4
    port map (
            O => \N__33934\,
            I => \indice_RNIS8333_5\
        );

    \I__7973\ : InMux
    port map (
            O => \N__33929\,
            I => \N__33926\
        );

    \I__7972\ : LocalMux
    port map (
            O => \N__33926\,
            I => \N__33923\
        );

    \I__7971\ : Span4Mux_h
    port map (
            O => \N__33923\,
            I => \N__33920\
        );

    \I__7970\ : Span4Mux_h
    port map (
            O => \N__33920\,
            I => \N__33917\
        );

    \I__7969\ : Span4Mux_h
    port map (
            O => \N__33917\,
            I => \N__33914\
        );

    \I__7968\ : Odrv4
    port map (
            O => \N__33914\,
            I => \b2v_inst.addr_ram_iv_i_0_8\
        );

    \I__7967\ : CascadeMux
    port map (
            O => \N__33911\,
            I => \N__33908\
        );

    \I__7966\ : InMux
    port map (
            O => \N__33908\,
            I => \N__33905\
        );

    \I__7965\ : LocalMux
    port map (
            O => \N__33905\,
            I => \N__33902\
        );

    \I__7964\ : Span4Mux_v
    port map (
            O => \N__33902\,
            I => \N__33899\
        );

    \I__7963\ : Sp12to4
    port map (
            O => \N__33899\,
            I => \N__33896\
        );

    \I__7962\ : Odrv12
    port map (
            O => \N__33896\,
            I => \b2v_inst.addr_ram_iv_i_1_8\
        );

    \I__7961\ : CascadeMux
    port map (
            O => \N__33893\,
            I => \N__33889\
        );

    \I__7960\ : CascadeMux
    port map (
            O => \N__33892\,
            I => \N__33886\
        );

    \I__7959\ : CascadeBuf
    port map (
            O => \N__33889\,
            I => \N__33883\
        );

    \I__7958\ : CascadeBuf
    port map (
            O => \N__33886\,
            I => \N__33880\
        );

    \I__7957\ : CascadeMux
    port map (
            O => \N__33883\,
            I => \N__33877\
        );

    \I__7956\ : CascadeMux
    port map (
            O => \N__33880\,
            I => \N__33874\
        );

    \I__7955\ : CascadeBuf
    port map (
            O => \N__33877\,
            I => \N__33871\
        );

    \I__7954\ : CascadeBuf
    port map (
            O => \N__33874\,
            I => \N__33868\
        );

    \I__7953\ : CascadeMux
    port map (
            O => \N__33871\,
            I => \N__33865\
        );

    \I__7952\ : CascadeMux
    port map (
            O => \N__33868\,
            I => \N__33862\
        );

    \I__7951\ : CascadeBuf
    port map (
            O => \N__33865\,
            I => \N__33859\
        );

    \I__7950\ : CascadeBuf
    port map (
            O => \N__33862\,
            I => \N__33856\
        );

    \I__7949\ : CascadeMux
    port map (
            O => \N__33859\,
            I => \N__33853\
        );

    \I__7948\ : CascadeMux
    port map (
            O => \N__33856\,
            I => \N__33850\
        );

    \I__7947\ : CascadeBuf
    port map (
            O => \N__33853\,
            I => \N__33847\
        );

    \I__7946\ : CascadeBuf
    port map (
            O => \N__33850\,
            I => \N__33844\
        );

    \I__7945\ : CascadeMux
    port map (
            O => \N__33847\,
            I => \N__33841\
        );

    \I__7944\ : CascadeMux
    port map (
            O => \N__33844\,
            I => \N__33838\
        );

    \I__7943\ : CascadeBuf
    port map (
            O => \N__33841\,
            I => \N__33835\
        );

    \I__7942\ : CascadeBuf
    port map (
            O => \N__33838\,
            I => \N__33832\
        );

    \I__7941\ : CascadeMux
    port map (
            O => \N__33835\,
            I => \N__33829\
        );

    \I__7940\ : CascadeMux
    port map (
            O => \N__33832\,
            I => \N__33826\
        );

    \I__7939\ : InMux
    port map (
            O => \N__33829\,
            I => \N__33823\
        );

    \I__7938\ : InMux
    port map (
            O => \N__33826\,
            I => \N__33820\
        );

    \I__7937\ : LocalMux
    port map (
            O => \N__33823\,
            I => \N__33817\
        );

    \I__7936\ : LocalMux
    port map (
            O => \N__33820\,
            I => \indice_RNIBO333_8\
        );

    \I__7935\ : Odrv4
    port map (
            O => \N__33817\,
            I => \indice_RNIBO333_8\
        );

    \I__7934\ : InMux
    port map (
            O => \N__33812\,
            I => \N__33809\
        );

    \I__7933\ : LocalMux
    port map (
            O => \N__33809\,
            I => \N__33806\
        );

    \I__7932\ : Span4Mux_v
    port map (
            O => \N__33806\,
            I => \N__33803\
        );

    \I__7931\ : Span4Mux_h
    port map (
            O => \N__33803\,
            I => \N__33800\
        );

    \I__7930\ : Odrv4
    port map (
            O => \N__33800\,
            I => \b2v_inst.addr_ram_iv_i_0_9\
        );

    \I__7929\ : CascadeMux
    port map (
            O => \N__33797\,
            I => \N__33794\
        );

    \I__7928\ : InMux
    port map (
            O => \N__33794\,
            I => \N__33791\
        );

    \I__7927\ : LocalMux
    port map (
            O => \N__33791\,
            I => \N__33788\
        );

    \I__7926\ : Span4Mux_h
    port map (
            O => \N__33788\,
            I => \N__33785\
        );

    \I__7925\ : Span4Mux_h
    port map (
            O => \N__33785\,
            I => \N__33782\
        );

    \I__7924\ : Odrv4
    port map (
            O => \N__33782\,
            I => \b2v_inst.addr_ram_iv_i_1_9\
        );

    \I__7923\ : CascadeMux
    port map (
            O => \N__33779\,
            I => \N__33775\
        );

    \I__7922\ : CascadeMux
    port map (
            O => \N__33778\,
            I => \N__33772\
        );

    \I__7921\ : CascadeBuf
    port map (
            O => \N__33775\,
            I => \N__33769\
        );

    \I__7920\ : CascadeBuf
    port map (
            O => \N__33772\,
            I => \N__33766\
        );

    \I__7919\ : CascadeMux
    port map (
            O => \N__33769\,
            I => \N__33763\
        );

    \I__7918\ : CascadeMux
    port map (
            O => \N__33766\,
            I => \N__33760\
        );

    \I__7917\ : CascadeBuf
    port map (
            O => \N__33763\,
            I => \N__33757\
        );

    \I__7916\ : CascadeBuf
    port map (
            O => \N__33760\,
            I => \N__33754\
        );

    \I__7915\ : CascadeMux
    port map (
            O => \N__33757\,
            I => \N__33751\
        );

    \I__7914\ : CascadeMux
    port map (
            O => \N__33754\,
            I => \N__33748\
        );

    \I__7913\ : CascadeBuf
    port map (
            O => \N__33751\,
            I => \N__33745\
        );

    \I__7912\ : CascadeBuf
    port map (
            O => \N__33748\,
            I => \N__33742\
        );

    \I__7911\ : CascadeMux
    port map (
            O => \N__33745\,
            I => \N__33739\
        );

    \I__7910\ : CascadeMux
    port map (
            O => \N__33742\,
            I => \N__33736\
        );

    \I__7909\ : CascadeBuf
    port map (
            O => \N__33739\,
            I => \N__33733\
        );

    \I__7908\ : CascadeBuf
    port map (
            O => \N__33736\,
            I => \N__33730\
        );

    \I__7907\ : CascadeMux
    port map (
            O => \N__33733\,
            I => \N__33727\
        );

    \I__7906\ : CascadeMux
    port map (
            O => \N__33730\,
            I => \N__33724\
        );

    \I__7905\ : CascadeBuf
    port map (
            O => \N__33727\,
            I => \N__33721\
        );

    \I__7904\ : CascadeBuf
    port map (
            O => \N__33724\,
            I => \N__33718\
        );

    \I__7903\ : CascadeMux
    port map (
            O => \N__33721\,
            I => \N__33715\
        );

    \I__7902\ : CascadeMux
    port map (
            O => \N__33718\,
            I => \N__33712\
        );

    \I__7901\ : InMux
    port map (
            O => \N__33715\,
            I => \N__33709\
        );

    \I__7900\ : InMux
    port map (
            O => \N__33712\,
            I => \N__33706\
        );

    \I__7899\ : LocalMux
    port map (
            O => \N__33709\,
            I => \N__33703\
        );

    \I__7898\ : LocalMux
    port map (
            O => \N__33706\,
            I => \indice_RNIGT333_9\
        );

    \I__7897\ : Odrv4
    port map (
            O => \N__33703\,
            I => \indice_RNIGT333_9\
        );

    \I__7896\ : InMux
    port map (
            O => \N__33698\,
            I => \N__33695\
        );

    \I__7895\ : LocalMux
    port map (
            O => \N__33695\,
            I => \N__33692\
        );

    \I__7894\ : Span4Mux_v
    port map (
            O => \N__33692\,
            I => \N__33689\
        );

    \I__7893\ : Odrv4
    port map (
            O => \N__33689\,
            I => \N_115_i\
        );

    \I__7892\ : CascadeMux
    port map (
            O => \N__33686\,
            I => \N__33683\
        );

    \I__7891\ : InMux
    port map (
            O => \N__33683\,
            I => \N__33679\
        );

    \I__7890\ : CascadeMux
    port map (
            O => \N__33682\,
            I => \N__33676\
        );

    \I__7889\ : LocalMux
    port map (
            O => \N__33679\,
            I => \N__33673\
        );

    \I__7888\ : InMux
    port map (
            O => \N__33676\,
            I => \N__33670\
        );

    \I__7887\ : Span4Mux_v
    port map (
            O => \N__33673\,
            I => \N__33664\
        );

    \I__7886\ : LocalMux
    port map (
            O => \N__33670\,
            I => \N__33664\
        );

    \I__7885\ : InMux
    port map (
            O => \N__33669\,
            I => \N__33661\
        );

    \I__7884\ : Span4Mux_h
    port map (
            O => \N__33664\,
            I => \N__33658\
        );

    \I__7883\ : LocalMux
    port map (
            O => \N__33661\,
            I => \N__33655\
        );

    \I__7882\ : Span4Mux_v
    port map (
            O => \N__33658\,
            I => \N__33652\
        );

    \I__7881\ : Span4Mux_h
    port map (
            O => \N__33655\,
            I => \N__33649\
        );

    \I__7880\ : Sp12to4
    port map (
            O => \N__33652\,
            I => \N__33645\
        );

    \I__7879\ : Span4Mux_h
    port map (
            O => \N__33649\,
            I => \N__33642\
        );

    \I__7878\ : InMux
    port map (
            O => \N__33648\,
            I => \N__33639\
        );

    \I__7877\ : Odrv12
    port map (
            O => \N__33645\,
            I => b2v_inst_data_a_escribir_10
        );

    \I__7876\ : Odrv4
    port map (
            O => \N__33642\,
            I => b2v_inst_data_a_escribir_10
        );

    \I__7875\ : LocalMux
    port map (
            O => \N__33639\,
            I => b2v_inst_data_a_escribir_10
        );

    \I__7874\ : InMux
    port map (
            O => \N__33632\,
            I => \N__33629\
        );

    \I__7873\ : LocalMux
    port map (
            O => \N__33629\,
            I => \N__33626\
        );

    \I__7872\ : Span4Mux_v
    port map (
            O => \N__33626\,
            I => \N__33623\
        );

    \I__7871\ : Odrv4
    port map (
            O => \N__33623\,
            I => \N_110_i\
        );

    \I__7870\ : InMux
    port map (
            O => \N__33620\,
            I => \N__33617\
        );

    \I__7869\ : LocalMux
    port map (
            O => \N__33617\,
            I => \N__33614\
        );

    \I__7868\ : Span4Mux_h
    port map (
            O => \N__33614\,
            I => \N__33611\
        );

    \I__7867\ : Span4Mux_h
    port map (
            O => \N__33611\,
            I => \N__33608\
        );

    \I__7866\ : Odrv4
    port map (
            O => \N__33608\,
            I => \b2v_inst.addr_ram_iv_i_0_0\
        );

    \I__7865\ : CascadeMux
    port map (
            O => \N__33605\,
            I => \N__33602\
        );

    \I__7864\ : InMux
    port map (
            O => \N__33602\,
            I => \N__33599\
        );

    \I__7863\ : LocalMux
    port map (
            O => \N__33599\,
            I => \N__33596\
        );

    \I__7862\ : Span12Mux_s9_h
    port map (
            O => \N__33596\,
            I => \N__33593\
        );

    \I__7861\ : Odrv12
    port map (
            O => \N__33593\,
            I => \b2v_inst.addr_ram_iv_i_1_0\
        );

    \I__7860\ : CascadeMux
    port map (
            O => \N__33590\,
            I => \N__33586\
        );

    \I__7859\ : CascadeMux
    port map (
            O => \N__33589\,
            I => \N__33583\
        );

    \I__7858\ : CascadeBuf
    port map (
            O => \N__33586\,
            I => \N__33580\
        );

    \I__7857\ : CascadeBuf
    port map (
            O => \N__33583\,
            I => \N__33577\
        );

    \I__7856\ : CascadeMux
    port map (
            O => \N__33580\,
            I => \N__33574\
        );

    \I__7855\ : CascadeMux
    port map (
            O => \N__33577\,
            I => \N__33571\
        );

    \I__7854\ : CascadeBuf
    port map (
            O => \N__33574\,
            I => \N__33568\
        );

    \I__7853\ : CascadeBuf
    port map (
            O => \N__33571\,
            I => \N__33565\
        );

    \I__7852\ : CascadeMux
    port map (
            O => \N__33568\,
            I => \N__33562\
        );

    \I__7851\ : CascadeMux
    port map (
            O => \N__33565\,
            I => \N__33559\
        );

    \I__7850\ : CascadeBuf
    port map (
            O => \N__33562\,
            I => \N__33556\
        );

    \I__7849\ : CascadeBuf
    port map (
            O => \N__33559\,
            I => \N__33553\
        );

    \I__7848\ : CascadeMux
    port map (
            O => \N__33556\,
            I => \N__33550\
        );

    \I__7847\ : CascadeMux
    port map (
            O => \N__33553\,
            I => \N__33547\
        );

    \I__7846\ : CascadeBuf
    port map (
            O => \N__33550\,
            I => \N__33544\
        );

    \I__7845\ : CascadeBuf
    port map (
            O => \N__33547\,
            I => \N__33541\
        );

    \I__7844\ : CascadeMux
    port map (
            O => \N__33544\,
            I => \N__33538\
        );

    \I__7843\ : CascadeMux
    port map (
            O => \N__33541\,
            I => \N__33535\
        );

    \I__7842\ : CascadeBuf
    port map (
            O => \N__33538\,
            I => \N__33532\
        );

    \I__7841\ : CascadeBuf
    port map (
            O => \N__33535\,
            I => \N__33529\
        );

    \I__7840\ : CascadeMux
    port map (
            O => \N__33532\,
            I => \N__33526\
        );

    \I__7839\ : CascadeMux
    port map (
            O => \N__33529\,
            I => \N__33523\
        );

    \I__7838\ : InMux
    port map (
            O => \N__33526\,
            I => \N__33520\
        );

    \I__7837\ : InMux
    port map (
            O => \N__33523\,
            I => \N__33517\
        );

    \I__7836\ : LocalMux
    port map (
            O => \N__33520\,
            I => \indice_RNI3F233_0\
        );

    \I__7835\ : LocalMux
    port map (
            O => \N__33517\,
            I => \indice_RNI3F233_0\
        );

    \I__7834\ : InMux
    port map (
            O => \N__33512\,
            I => \N__33509\
        );

    \I__7833\ : LocalMux
    port map (
            O => \N__33509\,
            I => \N__33506\
        );

    \I__7832\ : Span4Mux_v
    port map (
            O => \N__33506\,
            I => \N__33503\
        );

    \I__7831\ : Span4Mux_h
    port map (
            O => \N__33503\,
            I => \N__33500\
        );

    \I__7830\ : Span4Mux_h
    port map (
            O => \N__33500\,
            I => \N__33497\
        );

    \I__7829\ : Odrv4
    port map (
            O => \N__33497\,
            I => \b2v_inst.addr_ram_iv_i_0_10\
        );

    \I__7828\ : CascadeMux
    port map (
            O => \N__33494\,
            I => \N__33491\
        );

    \I__7827\ : InMux
    port map (
            O => \N__33491\,
            I => \N__33488\
        );

    \I__7826\ : LocalMux
    port map (
            O => \N__33488\,
            I => \N__33485\
        );

    \I__7825\ : Span4Mux_h
    port map (
            O => \N__33485\,
            I => \N__33482\
        );

    \I__7824\ : Span4Mux_h
    port map (
            O => \N__33482\,
            I => \N__33479\
        );

    \I__7823\ : Odrv4
    port map (
            O => \N__33479\,
            I => \b2v_inst.addr_ram_iv_i_1_10\
        );

    \I__7822\ : CascadeMux
    port map (
            O => \N__33476\,
            I => \N__33472\
        );

    \I__7821\ : CascadeMux
    port map (
            O => \N__33475\,
            I => \N__33469\
        );

    \I__7820\ : CascadeBuf
    port map (
            O => \N__33472\,
            I => \N__33466\
        );

    \I__7819\ : CascadeBuf
    port map (
            O => \N__33469\,
            I => \N__33463\
        );

    \I__7818\ : CascadeMux
    port map (
            O => \N__33466\,
            I => \N__33460\
        );

    \I__7817\ : CascadeMux
    port map (
            O => \N__33463\,
            I => \N__33457\
        );

    \I__7816\ : CascadeBuf
    port map (
            O => \N__33460\,
            I => \N__33454\
        );

    \I__7815\ : CascadeBuf
    port map (
            O => \N__33457\,
            I => \N__33451\
        );

    \I__7814\ : CascadeMux
    port map (
            O => \N__33454\,
            I => \N__33448\
        );

    \I__7813\ : CascadeMux
    port map (
            O => \N__33451\,
            I => \N__33445\
        );

    \I__7812\ : CascadeBuf
    port map (
            O => \N__33448\,
            I => \N__33442\
        );

    \I__7811\ : CascadeBuf
    port map (
            O => \N__33445\,
            I => \N__33439\
        );

    \I__7810\ : CascadeMux
    port map (
            O => \N__33442\,
            I => \N__33436\
        );

    \I__7809\ : CascadeMux
    port map (
            O => \N__33439\,
            I => \N__33433\
        );

    \I__7808\ : CascadeBuf
    port map (
            O => \N__33436\,
            I => \N__33430\
        );

    \I__7807\ : CascadeBuf
    port map (
            O => \N__33433\,
            I => \N__33427\
        );

    \I__7806\ : CascadeMux
    port map (
            O => \N__33430\,
            I => \N__33424\
        );

    \I__7805\ : CascadeMux
    port map (
            O => \N__33427\,
            I => \N__33421\
        );

    \I__7804\ : CascadeBuf
    port map (
            O => \N__33424\,
            I => \N__33418\
        );

    \I__7803\ : CascadeBuf
    port map (
            O => \N__33421\,
            I => \N__33415\
        );

    \I__7802\ : CascadeMux
    port map (
            O => \N__33418\,
            I => \N__33412\
        );

    \I__7801\ : CascadeMux
    port map (
            O => \N__33415\,
            I => \N__33409\
        );

    \I__7800\ : InMux
    port map (
            O => \N__33412\,
            I => \N__33406\
        );

    \I__7799\ : InMux
    port map (
            O => \N__33409\,
            I => \N__33403\
        );

    \I__7798\ : LocalMux
    port map (
            O => \N__33406\,
            I => \N_37\
        );

    \I__7797\ : LocalMux
    port map (
            O => \N__33403\,
            I => \N_37\
        );

    \I__7796\ : CascadeMux
    port map (
            O => \N__33398\,
            I => \N__33394\
        );

    \I__7795\ : CascadeMux
    port map (
            O => \N__33397\,
            I => \N__33391\
        );

    \I__7794\ : InMux
    port map (
            O => \N__33394\,
            I => \N__33388\
        );

    \I__7793\ : InMux
    port map (
            O => \N__33391\,
            I => \N__33385\
        );

    \I__7792\ : LocalMux
    port map (
            O => \N__33388\,
            I => \N__33382\
        );

    \I__7791\ : LocalMux
    port map (
            O => \N__33385\,
            I => \N__33375\
        );

    \I__7790\ : Sp12to4
    port map (
            O => \N__33382\,
            I => \N__33375\
        );

    \I__7789\ : InMux
    port map (
            O => \N__33381\,
            I => \N__33372\
        );

    \I__7788\ : InMux
    port map (
            O => \N__33380\,
            I => \N__33369\
        );

    \I__7787\ : Span12Mux_h
    port map (
            O => \N__33375\,
            I => \N__33366\
        );

    \I__7786\ : LocalMux
    port map (
            O => \N__33372\,
            I => \N__33361\
        );

    \I__7785\ : LocalMux
    port map (
            O => \N__33369\,
            I => \N__33361\
        );

    \I__7784\ : Odrv12
    port map (
            O => \N__33366\,
            I => b2v_inst_data_a_escribir_8
        );

    \I__7783\ : Odrv12
    port map (
            O => \N__33361\,
            I => b2v_inst_data_a_escribir_8
        );

    \I__7782\ : InMux
    port map (
            O => \N__33356\,
            I => \N__33353\
        );

    \I__7781\ : LocalMux
    port map (
            O => \N__33353\,
            I => \N__33350\
        );

    \I__7780\ : Odrv4
    port map (
            O => \N__33350\,
            I => \N_112_i\
        );

    \I__7779\ : InMux
    port map (
            O => \N__33347\,
            I => \N__33344\
        );

    \I__7778\ : LocalMux
    port map (
            O => \N__33344\,
            I => \b2v_inst.un16_data_ram_cantidad_o_cry_3_c_RNIBDEOZ0\
        );

    \I__7777\ : CascadeMux
    port map (
            O => \N__33341\,
            I => \N__33338\
        );

    \I__7776\ : InMux
    port map (
            O => \N__33338\,
            I => \N__33333\
        );

    \I__7775\ : InMux
    port map (
            O => \N__33337\,
            I => \N__33330\
        );

    \I__7774\ : CascadeMux
    port map (
            O => \N__33336\,
            I => \N__33326\
        );

    \I__7773\ : LocalMux
    port map (
            O => \N__33333\,
            I => \N__33322\
        );

    \I__7772\ : LocalMux
    port map (
            O => \N__33330\,
            I => \N__33319\
        );

    \I__7771\ : CascadeMux
    port map (
            O => \N__33329\,
            I => \N__33316\
        );

    \I__7770\ : InMux
    port map (
            O => \N__33326\,
            I => \N__33313\
        );

    \I__7769\ : InMux
    port map (
            O => \N__33325\,
            I => \N__33310\
        );

    \I__7768\ : Span4Mux_v
    port map (
            O => \N__33322\,
            I => \N__33305\
        );

    \I__7767\ : Span4Mux_v
    port map (
            O => \N__33319\,
            I => \N__33305\
        );

    \I__7766\ : InMux
    port map (
            O => \N__33316\,
            I => \N__33302\
        );

    \I__7765\ : LocalMux
    port map (
            O => \N__33313\,
            I => \N__33297\
        );

    \I__7764\ : LocalMux
    port map (
            O => \N__33310\,
            I => \N__33297\
        );

    \I__7763\ : Sp12to4
    port map (
            O => \N__33305\,
            I => \N__33294\
        );

    \I__7762\ : LocalMux
    port map (
            O => \N__33302\,
            I => \N__33291\
        );

    \I__7761\ : Span4Mux_v
    port map (
            O => \N__33297\,
            I => \N__33288\
        );

    \I__7760\ : Span12Mux_h
    port map (
            O => \N__33294\,
            I => \N__33285\
        );

    \I__7759\ : Span4Mux_h
    port map (
            O => \N__33291\,
            I => \N__33280\
        );

    \I__7758\ : Span4Mux_h
    port map (
            O => \N__33288\,
            I => \N__33280\
        );

    \I__7757\ : Odrv12
    port map (
            O => \N__33285\,
            I => b2v_inst_data_a_escribir_4
        );

    \I__7756\ : Odrv4
    port map (
            O => \N__33280\,
            I => b2v_inst_data_a_escribir_4
        );

    \I__7755\ : InMux
    port map (
            O => \N__33275\,
            I => \N__33272\
        );

    \I__7754\ : LocalMux
    port map (
            O => \N__33272\,
            I => \N__33269\
        );

    \I__7753\ : Span4Mux_h
    port map (
            O => \N__33269\,
            I => \N__33266\
        );

    \I__7752\ : Odrv4
    port map (
            O => \N__33266\,
            I => \N_549_i\
        );

    \I__7751\ : InMux
    port map (
            O => \N__33263\,
            I => \N__33260\
        );

    \I__7750\ : LocalMux
    port map (
            O => \N__33260\,
            I => \b2v_inst.un16_data_ram_cantidad_o_cry_2_c_RNI9ADOZ0\
        );

    \I__7749\ : CascadeMux
    port map (
            O => \N__33257\,
            I => \N__33251\
        );

    \I__7748\ : InMux
    port map (
            O => \N__33256\,
            I => \N__33248\
        );

    \I__7747\ : CascadeMux
    port map (
            O => \N__33255\,
            I => \N__33245\
        );

    \I__7746\ : InMux
    port map (
            O => \N__33254\,
            I => \N__33241\
        );

    \I__7745\ : InMux
    port map (
            O => \N__33251\,
            I => \N__33238\
        );

    \I__7744\ : LocalMux
    port map (
            O => \N__33248\,
            I => \N__33235\
        );

    \I__7743\ : InMux
    port map (
            O => \N__33245\,
            I => \N__33232\
        );

    \I__7742\ : InMux
    port map (
            O => \N__33244\,
            I => \N__33229\
        );

    \I__7741\ : LocalMux
    port map (
            O => \N__33241\,
            I => \N__33226\
        );

    \I__7740\ : LocalMux
    port map (
            O => \N__33238\,
            I => \N__33223\
        );

    \I__7739\ : Span4Mux_h
    port map (
            O => \N__33235\,
            I => \N__33218\
        );

    \I__7738\ : LocalMux
    port map (
            O => \N__33232\,
            I => \N__33218\
        );

    \I__7737\ : LocalMux
    port map (
            O => \N__33229\,
            I => \N__33215\
        );

    \I__7736\ : Span4Mux_v
    port map (
            O => \N__33226\,
            I => \N__33212\
        );

    \I__7735\ : Span4Mux_v
    port map (
            O => \N__33223\,
            I => \N__33207\
        );

    \I__7734\ : Span4Mux_h
    port map (
            O => \N__33218\,
            I => \N__33207\
        );

    \I__7733\ : Span4Mux_h
    port map (
            O => \N__33215\,
            I => \N__33200\
        );

    \I__7732\ : Span4Mux_h
    port map (
            O => \N__33212\,
            I => \N__33200\
        );

    \I__7731\ : Span4Mux_h
    port map (
            O => \N__33207\,
            I => \N__33200\
        );

    \I__7730\ : Odrv4
    port map (
            O => \N__33200\,
            I => b2v_inst_data_a_escribir_3
        );

    \I__7729\ : InMux
    port map (
            O => \N__33197\,
            I => \N__33194\
        );

    \I__7728\ : LocalMux
    port map (
            O => \N__33194\,
            I => \N__33191\
        );

    \I__7727\ : Odrv4
    port map (
            O => \N__33191\,
            I => \N_551_i\
        );

    \I__7726\ : InMux
    port map (
            O => \N__33188\,
            I => \N__33184\
        );

    \I__7725\ : InMux
    port map (
            O => \N__33187\,
            I => \N__33181\
        );

    \I__7724\ : LocalMux
    port map (
            O => \N__33184\,
            I => \N__33177\
        );

    \I__7723\ : LocalMux
    port map (
            O => \N__33181\,
            I => \N__33174\
        );

    \I__7722\ : InMux
    port map (
            O => \N__33180\,
            I => \N__33171\
        );

    \I__7721\ : Span4Mux_v
    port map (
            O => \N__33177\,
            I => \N__33168\
        );

    \I__7720\ : Span4Mux_h
    port map (
            O => \N__33174\,
            I => \N__33164\
        );

    \I__7719\ : LocalMux
    port map (
            O => \N__33171\,
            I => \N__33159\
        );

    \I__7718\ : Sp12to4
    port map (
            O => \N__33168\,
            I => \N__33159\
        );

    \I__7717\ : InMux
    port map (
            O => \N__33167\,
            I => \N__33156\
        );

    \I__7716\ : Span4Mux_h
    port map (
            O => \N__33164\,
            I => \N__33153\
        );

    \I__7715\ : Odrv12
    port map (
            O => \N__33159\,
            I => \b2v_inst.N_481\
        );

    \I__7714\ : LocalMux
    port map (
            O => \N__33156\,
            I => \b2v_inst.N_481\
        );

    \I__7713\ : Odrv4
    port map (
            O => \N__33153\,
            I => \b2v_inst.N_481\
        );

    \I__7712\ : InMux
    port map (
            O => \N__33146\,
            I => \N__33143\
        );

    \I__7711\ : LocalMux
    port map (
            O => \N__33143\,
            I => \N_121_i\
        );

    \I__7710\ : CascadeMux
    port map (
            O => \N__33140\,
            I => \N__33136\
        );

    \I__7709\ : InMux
    port map (
            O => \N__33139\,
            I => \N__33132\
        );

    \I__7708\ : InMux
    port map (
            O => \N__33136\,
            I => \N__33128\
        );

    \I__7707\ : InMux
    port map (
            O => \N__33135\,
            I => \N__33125\
        );

    \I__7706\ : LocalMux
    port map (
            O => \N__33132\,
            I => \N__33121\
        );

    \I__7705\ : CascadeMux
    port map (
            O => \N__33131\,
            I => \N__33118\
        );

    \I__7704\ : LocalMux
    port map (
            O => \N__33128\,
            I => \N__33115\
        );

    \I__7703\ : LocalMux
    port map (
            O => \N__33125\,
            I => \N__33112\
        );

    \I__7702\ : InMux
    port map (
            O => \N__33124\,
            I => \N__33109\
        );

    \I__7701\ : Span4Mux_v
    port map (
            O => \N__33121\,
            I => \N__33106\
        );

    \I__7700\ : InMux
    port map (
            O => \N__33118\,
            I => \N__33103\
        );

    \I__7699\ : Span4Mux_h
    port map (
            O => \N__33115\,
            I => \N__33100\
        );

    \I__7698\ : Span4Mux_v
    port map (
            O => \N__33112\,
            I => \N__33097\
        );

    \I__7697\ : LocalMux
    port map (
            O => \N__33109\,
            I => \N__33094\
        );

    \I__7696\ : Span4Mux_h
    port map (
            O => \N__33106\,
            I => \N__33089\
        );

    \I__7695\ : LocalMux
    port map (
            O => \N__33103\,
            I => \N__33089\
        );

    \I__7694\ : Span4Mux_v
    port map (
            O => \N__33100\,
            I => \N__33084\
        );

    \I__7693\ : Span4Mux_h
    port map (
            O => \N__33097\,
            I => \N__33084\
        );

    \I__7692\ : Span12Mux_v
    port map (
            O => \N__33094\,
            I => \N__33081\
        );

    \I__7691\ : Span4Mux_h
    port map (
            O => \N__33089\,
            I => \N__33078\
        );

    \I__7690\ : Odrv4
    port map (
            O => \N__33084\,
            I => b2v_inst_data_a_escribir_2
        );

    \I__7689\ : Odrv12
    port map (
            O => \N__33081\,
            I => b2v_inst_data_a_escribir_2
        );

    \I__7688\ : Odrv4
    port map (
            O => \N__33078\,
            I => b2v_inst_data_a_escribir_2
        );

    \I__7687\ : InMux
    port map (
            O => \N__33071\,
            I => \N__33068\
        );

    \I__7686\ : LocalMux
    port map (
            O => \N__33068\,
            I => \N__33065\
        );

    \I__7685\ : Odrv4
    port map (
            O => \N__33065\,
            I => \N_118_i\
        );

    \I__7684\ : InMux
    port map (
            O => \N__33062\,
            I => \N__33058\
        );

    \I__7683\ : InMux
    port map (
            O => \N__33061\,
            I => \N__33055\
        );

    \I__7682\ : LocalMux
    port map (
            O => \N__33058\,
            I => \N__33051\
        );

    \I__7681\ : LocalMux
    port map (
            O => \N__33055\,
            I => \N__33047\
        );

    \I__7680\ : InMux
    port map (
            O => \N__33054\,
            I => \N__33044\
        );

    \I__7679\ : Span4Mux_h
    port map (
            O => \N__33051\,
            I => \N__33041\
        );

    \I__7678\ : InMux
    port map (
            O => \N__33050\,
            I => \N__33038\
        );

    \I__7677\ : Span4Mux_h
    port map (
            O => \N__33047\,
            I => \N__33035\
        );

    \I__7676\ : LocalMux
    port map (
            O => \N__33044\,
            I => \N__33030\
        );

    \I__7675\ : Span4Mux_h
    port map (
            O => \N__33041\,
            I => \N__33030\
        );

    \I__7674\ : LocalMux
    port map (
            O => \N__33038\,
            I => \N__33027\
        );

    \I__7673\ : Odrv4
    port map (
            O => \N__33035\,
            I => \SYNTHESIZED_WIRE_3_4\
        );

    \I__7672\ : Odrv4
    port map (
            O => \N__33030\,
            I => \SYNTHESIZED_WIRE_3_4\
        );

    \I__7671\ : Odrv4
    port map (
            O => \N__33027\,
            I => \SYNTHESIZED_WIRE_3_4\
        );

    \I__7670\ : InMux
    port map (
            O => \N__33020\,
            I => \N__33016\
        );

    \I__7669\ : InMux
    port map (
            O => \N__33019\,
            I => \N__33011\
        );

    \I__7668\ : LocalMux
    port map (
            O => \N__33016\,
            I => \N__33007\
        );

    \I__7667\ : InMux
    port map (
            O => \N__33015\,
            I => \N__33004\
        );

    \I__7666\ : InMux
    port map (
            O => \N__33014\,
            I => \N__33001\
        );

    \I__7665\ : LocalMux
    port map (
            O => \N__33011\,
            I => \N__32998\
        );

    \I__7664\ : CascadeMux
    port map (
            O => \N__33010\,
            I => \N__32995\
        );

    \I__7663\ : Span4Mux_v
    port map (
            O => \N__33007\,
            I => \N__32992\
        );

    \I__7662\ : LocalMux
    port map (
            O => \N__33004\,
            I => \N__32989\
        );

    \I__7661\ : LocalMux
    port map (
            O => \N__33001\,
            I => \N__32986\
        );

    \I__7660\ : Span4Mux_h
    port map (
            O => \N__32998\,
            I => \N__32983\
        );

    \I__7659\ : InMux
    port map (
            O => \N__32995\,
            I => \N__32980\
        );

    \I__7658\ : Span4Mux_h
    port map (
            O => \N__32992\,
            I => \N__32975\
        );

    \I__7657\ : Span4Mux_h
    port map (
            O => \N__32989\,
            I => \N__32975\
        );

    \I__7656\ : Odrv12
    port map (
            O => \N__32986\,
            I => \b2v_inst.reg_ancho_2Z0Z_4\
        );

    \I__7655\ : Odrv4
    port map (
            O => \N__32983\,
            I => \b2v_inst.reg_ancho_2Z0Z_4\
        );

    \I__7654\ : LocalMux
    port map (
            O => \N__32980\,
            I => \b2v_inst.reg_ancho_2Z0Z_4\
        );

    \I__7653\ : Odrv4
    port map (
            O => \N__32975\,
            I => \b2v_inst.reg_ancho_2Z0Z_4\
        );

    \I__7652\ : CEMux
    port map (
            O => \N__32966\,
            I => \N__32960\
        );

    \I__7651\ : CEMux
    port map (
            O => \N__32965\,
            I => \N__32955\
        );

    \I__7650\ : CEMux
    port map (
            O => \N__32964\,
            I => \N__32952\
        );

    \I__7649\ : CEMux
    port map (
            O => \N__32963\,
            I => \N__32949\
        );

    \I__7648\ : LocalMux
    port map (
            O => \N__32960\,
            I => \N__32946\
        );

    \I__7647\ : CEMux
    port map (
            O => \N__32959\,
            I => \N__32943\
        );

    \I__7646\ : CEMux
    port map (
            O => \N__32958\,
            I => \N__32940\
        );

    \I__7645\ : LocalMux
    port map (
            O => \N__32955\,
            I => \N__32937\
        );

    \I__7644\ : LocalMux
    port map (
            O => \N__32952\,
            I => \N__32934\
        );

    \I__7643\ : LocalMux
    port map (
            O => \N__32949\,
            I => \N__32931\
        );

    \I__7642\ : Span4Mux_v
    port map (
            O => \N__32946\,
            I => \N__32925\
        );

    \I__7641\ : LocalMux
    port map (
            O => \N__32943\,
            I => \N__32925\
        );

    \I__7640\ : LocalMux
    port map (
            O => \N__32940\,
            I => \N__32922\
        );

    \I__7639\ : Span4Mux_v
    port map (
            O => \N__32937\,
            I => \N__32919\
        );

    \I__7638\ : Span4Mux_v
    port map (
            O => \N__32934\,
            I => \N__32914\
        );

    \I__7637\ : Span4Mux_h
    port map (
            O => \N__32931\,
            I => \N__32914\
        );

    \I__7636\ : CEMux
    port map (
            O => \N__32930\,
            I => \N__32911\
        );

    \I__7635\ : Span4Mux_h
    port map (
            O => \N__32925\,
            I => \N__32900\
        );

    \I__7634\ : Span4Mux_v
    port map (
            O => \N__32922\,
            I => \N__32900\
        );

    \I__7633\ : Span4Mux_h
    port map (
            O => \N__32919\,
            I => \N__32900\
        );

    \I__7632\ : Span4Mux_v
    port map (
            O => \N__32914\,
            I => \N__32900\
        );

    \I__7631\ : LocalMux
    port map (
            O => \N__32911\,
            I => \N__32900\
        );

    \I__7630\ : Span4Mux_h
    port map (
            O => \N__32900\,
            I => \N__32893\
        );

    \I__7629\ : InMux
    port map (
            O => \N__32899\,
            I => \N__32890\
        );

    \I__7628\ : InMux
    port map (
            O => \N__32898\,
            I => \N__32885\
        );

    \I__7627\ : InMux
    port map (
            O => \N__32897\,
            I => \N__32885\
        );

    \I__7626\ : InMux
    port map (
            O => \N__32896\,
            I => \N__32882\
        );

    \I__7625\ : Odrv4
    port map (
            O => \N__32893\,
            I => \b2v_inst.stateZ0Z_23\
        );

    \I__7624\ : LocalMux
    port map (
            O => \N__32890\,
            I => \b2v_inst.stateZ0Z_23\
        );

    \I__7623\ : LocalMux
    port map (
            O => \N__32885\,
            I => \b2v_inst.stateZ0Z_23\
        );

    \I__7622\ : LocalMux
    port map (
            O => \N__32882\,
            I => \b2v_inst.stateZ0Z_23\
        );

    \I__7621\ : CascadeMux
    port map (
            O => \N__32873\,
            I => \N__32869\
        );

    \I__7620\ : CascadeMux
    port map (
            O => \N__32872\,
            I => \N__32866\
        );

    \I__7619\ : InMux
    port map (
            O => \N__32869\,
            I => \N__32863\
        );

    \I__7618\ : InMux
    port map (
            O => \N__32866\,
            I => \N__32860\
        );

    \I__7617\ : LocalMux
    port map (
            O => \N__32863\,
            I => \N__32854\
        );

    \I__7616\ : LocalMux
    port map (
            O => \N__32860\,
            I => \N__32854\
        );

    \I__7615\ : InMux
    port map (
            O => \N__32859\,
            I => \N__32850\
        );

    \I__7614\ : Span4Mux_h
    port map (
            O => \N__32854\,
            I => \N__32847\
        );

    \I__7613\ : InMux
    port map (
            O => \N__32853\,
            I => \N__32844\
        );

    \I__7612\ : LocalMux
    port map (
            O => \N__32850\,
            I => \N__32841\
        );

    \I__7611\ : Span4Mux_h
    port map (
            O => \N__32847\,
            I => \N__32836\
        );

    \I__7610\ : LocalMux
    port map (
            O => \N__32844\,
            I => \N__32836\
        );

    \I__7609\ : Span4Mux_h
    port map (
            O => \N__32841\,
            I => \N__32833\
        );

    \I__7608\ : Span4Mux_v
    port map (
            O => \N__32836\,
            I => \N__32830\
        );

    \I__7607\ : Odrv4
    port map (
            O => \N__32833\,
            I => b2v_inst_data_a_escribir_9
        );

    \I__7606\ : Odrv4
    port map (
            O => \N__32830\,
            I => b2v_inst_data_a_escribir_9
        );

    \I__7605\ : InMux
    port map (
            O => \N__32825\,
            I => \N__32822\
        );

    \I__7604\ : LocalMux
    port map (
            O => \N__32822\,
            I => \N_111_i\
        );

    \I__7603\ : InMux
    port map (
            O => \N__32819\,
            I => \N__32816\
        );

    \I__7602\ : LocalMux
    port map (
            O => \N__32816\,
            I => \N__32813\
        );

    \I__7601\ : Span4Mux_h
    port map (
            O => \N__32813\,
            I => \N__32810\
        );

    \I__7600\ : Span4Mux_h
    port map (
            O => \N__32810\,
            I => \N__32807\
        );

    \I__7599\ : Span4Mux_h
    port map (
            O => \N__32807\,
            I => \N__32804\
        );

    \I__7598\ : Odrv4
    port map (
            O => \N__32804\,
            I => \b2v_inst.addr_ram_iv_i_1_6\
        );

    \I__7597\ : CascadeMux
    port map (
            O => \N__32801\,
            I => \N__32798\
        );

    \I__7596\ : InMux
    port map (
            O => \N__32798\,
            I => \N__32795\
        );

    \I__7595\ : LocalMux
    port map (
            O => \N__32795\,
            I => \N__32792\
        );

    \I__7594\ : Span12Mux_h
    port map (
            O => \N__32792\,
            I => \N__32789\
        );

    \I__7593\ : Odrv12
    port map (
            O => \N__32789\,
            I => \b2v_inst.addr_ram_iv_i_0_6\
        );

    \I__7592\ : CascadeMux
    port map (
            O => \N__32786\,
            I => \N__32782\
        );

    \I__7591\ : CascadeMux
    port map (
            O => \N__32785\,
            I => \N__32779\
        );

    \I__7590\ : CascadeBuf
    port map (
            O => \N__32782\,
            I => \N__32776\
        );

    \I__7589\ : CascadeBuf
    port map (
            O => \N__32779\,
            I => \N__32773\
        );

    \I__7588\ : CascadeMux
    port map (
            O => \N__32776\,
            I => \N__32770\
        );

    \I__7587\ : CascadeMux
    port map (
            O => \N__32773\,
            I => \N__32767\
        );

    \I__7586\ : CascadeBuf
    port map (
            O => \N__32770\,
            I => \N__32764\
        );

    \I__7585\ : CascadeBuf
    port map (
            O => \N__32767\,
            I => \N__32761\
        );

    \I__7584\ : CascadeMux
    port map (
            O => \N__32764\,
            I => \N__32758\
        );

    \I__7583\ : CascadeMux
    port map (
            O => \N__32761\,
            I => \N__32755\
        );

    \I__7582\ : CascadeBuf
    port map (
            O => \N__32758\,
            I => \N__32752\
        );

    \I__7581\ : CascadeBuf
    port map (
            O => \N__32755\,
            I => \N__32749\
        );

    \I__7580\ : CascadeMux
    port map (
            O => \N__32752\,
            I => \N__32746\
        );

    \I__7579\ : CascadeMux
    port map (
            O => \N__32749\,
            I => \N__32743\
        );

    \I__7578\ : CascadeBuf
    port map (
            O => \N__32746\,
            I => \N__32740\
        );

    \I__7577\ : CascadeBuf
    port map (
            O => \N__32743\,
            I => \N__32737\
        );

    \I__7576\ : CascadeMux
    port map (
            O => \N__32740\,
            I => \N__32734\
        );

    \I__7575\ : CascadeMux
    port map (
            O => \N__32737\,
            I => \N__32731\
        );

    \I__7574\ : CascadeBuf
    port map (
            O => \N__32734\,
            I => \N__32728\
        );

    \I__7573\ : CascadeBuf
    port map (
            O => \N__32731\,
            I => \N__32725\
        );

    \I__7572\ : CascadeMux
    port map (
            O => \N__32728\,
            I => \N__32722\
        );

    \I__7571\ : CascadeMux
    port map (
            O => \N__32725\,
            I => \N__32719\
        );

    \I__7570\ : InMux
    port map (
            O => \N__32722\,
            I => \N__32716\
        );

    \I__7569\ : InMux
    port map (
            O => \N__32719\,
            I => \N__32713\
        );

    \I__7568\ : LocalMux
    port map (
            O => \N__32716\,
            I => \N__32710\
        );

    \I__7567\ : LocalMux
    port map (
            O => \N__32713\,
            I => \N_298\
        );

    \I__7566\ : Odrv4
    port map (
            O => \N__32710\,
            I => \N_298\
        );

    \I__7565\ : CascadeMux
    port map (
            O => \N__32705\,
            I => \N__32702\
        );

    \I__7564\ : InMux
    port map (
            O => \N__32702\,
            I => \N__32699\
        );

    \I__7563\ : LocalMux
    port map (
            O => \N__32699\,
            I => \N__32696\
        );

    \I__7562\ : Span4Mux_h
    port map (
            O => \N__32696\,
            I => \N__32693\
        );

    \I__7561\ : Odrv4
    port map (
            O => \N__32693\,
            I => \SYNTHESIZED_WIRE_1_0\
        );

    \I__7560\ : CascadeMux
    port map (
            O => \N__32690\,
            I => \N__32687\
        );

    \I__7559\ : InMux
    port map (
            O => \N__32687\,
            I => \N__32684\
        );

    \I__7558\ : LocalMux
    port map (
            O => \N__32684\,
            I => \N__32681\
        );

    \I__7557\ : Odrv12
    port map (
            O => \N__32681\,
            I => \SYNTHESIZED_WIRE_1_1\
        );

    \I__7556\ : CascadeMux
    port map (
            O => \N__32678\,
            I => \N__32675\
        );

    \I__7555\ : InMux
    port map (
            O => \N__32675\,
            I => \N__32672\
        );

    \I__7554\ : LocalMux
    port map (
            O => \N__32672\,
            I => \N__32669\
        );

    \I__7553\ : Span4Mux_h
    port map (
            O => \N__32669\,
            I => \N__32666\
        );

    \I__7552\ : Span4Mux_v
    port map (
            O => \N__32666\,
            I => \N__32663\
        );

    \I__7551\ : Odrv4
    port map (
            O => \N__32663\,
            I => \SYNTHESIZED_WIRE_1_4\
        );

    \I__7550\ : InMux
    port map (
            O => \N__32660\,
            I => \N__32657\
        );

    \I__7549\ : LocalMux
    port map (
            O => \N__32657\,
            I => \N__32653\
        );

    \I__7548\ : InMux
    port map (
            O => \N__32656\,
            I => \N__32649\
        );

    \I__7547\ : Span4Mux_h
    port map (
            O => \N__32653\,
            I => \N__32646\
        );

    \I__7546\ : InMux
    port map (
            O => \N__32652\,
            I => \N__32643\
        );

    \I__7545\ : LocalMux
    port map (
            O => \N__32649\,
            I => b2v_inst_cantidad_temp_2
        );

    \I__7544\ : Odrv4
    port map (
            O => \N__32646\,
            I => b2v_inst_cantidad_temp_2
        );

    \I__7543\ : LocalMux
    port map (
            O => \N__32643\,
            I => b2v_inst_cantidad_temp_2
        );

    \I__7542\ : InMux
    port map (
            O => \N__32636\,
            I => \b2v_inst.un16_data_ram_cantidad_o_cry_1\
        );

    \I__7541\ : InMux
    port map (
            O => \N__32633\,
            I => \b2v_inst.un16_data_ram_cantidad_o_cry_2\
        );

    \I__7540\ : InMux
    port map (
            O => \N__32630\,
            I => \N__32627\
        );

    \I__7539\ : LocalMux
    port map (
            O => \N__32627\,
            I => \N__32624\
        );

    \I__7538\ : Span4Mux_h
    port map (
            O => \N__32624\,
            I => \N__32620\
        );

    \I__7537\ : InMux
    port map (
            O => \N__32623\,
            I => \N__32616\
        );

    \I__7536\ : Span4Mux_h
    port map (
            O => \N__32620\,
            I => \N__32613\
        );

    \I__7535\ : InMux
    port map (
            O => \N__32619\,
            I => \N__32610\
        );

    \I__7534\ : LocalMux
    port map (
            O => \N__32616\,
            I => b2v_inst_cantidad_temp_4
        );

    \I__7533\ : Odrv4
    port map (
            O => \N__32613\,
            I => b2v_inst_cantidad_temp_4
        );

    \I__7532\ : LocalMux
    port map (
            O => \N__32610\,
            I => b2v_inst_cantidad_temp_4
        );

    \I__7531\ : InMux
    port map (
            O => \N__32603\,
            I => \b2v_inst.un16_data_ram_cantidad_o_cry_3\
        );

    \I__7530\ : CascadeMux
    port map (
            O => \N__32600\,
            I => \N__32596\
        );

    \I__7529\ : InMux
    port map (
            O => \N__32599\,
            I => \N__32593\
        );

    \I__7528\ : InMux
    port map (
            O => \N__32596\,
            I => \N__32590\
        );

    \I__7527\ : LocalMux
    port map (
            O => \N__32593\,
            I => \N__32587\
        );

    \I__7526\ : LocalMux
    port map (
            O => \N__32590\,
            I => \N__32583\
        );

    \I__7525\ : Span4Mux_v
    port map (
            O => \N__32587\,
            I => \N__32580\
        );

    \I__7524\ : InMux
    port map (
            O => \N__32586\,
            I => \N__32577\
        );

    \I__7523\ : Sp12to4
    port map (
            O => \N__32583\,
            I => \N__32572\
        );

    \I__7522\ : Sp12to4
    port map (
            O => \N__32580\,
            I => \N__32572\
        );

    \I__7521\ : LocalMux
    port map (
            O => \N__32577\,
            I => b2v_inst_cantidad_temp_5
        );

    \I__7520\ : Odrv12
    port map (
            O => \N__32572\,
            I => b2v_inst_cantidad_temp_5
        );

    \I__7519\ : InMux
    port map (
            O => \N__32567\,
            I => \b2v_inst.un16_data_ram_cantidad_o_cry_4\
        );

    \I__7518\ : InMux
    port map (
            O => \N__32564\,
            I => \N__32561\
        );

    \I__7517\ : LocalMux
    port map (
            O => \N__32561\,
            I => \b2v_inst.un16_data_ram_cantidad_o_cry_1_c_RNI77COZ0\
        );

    \I__7516\ : InMux
    port map (
            O => \N__32558\,
            I => \N__32555\
        );

    \I__7515\ : LocalMux
    port map (
            O => \N__32555\,
            I => \N__32552\
        );

    \I__7514\ : Span4Mux_h
    port map (
            O => \N__32552\,
            I => \N__32549\
        );

    \I__7513\ : Odrv4
    port map (
            O => \N__32549\,
            I => \N_553_i\
        );

    \I__7512\ : InMux
    port map (
            O => \N__32546\,
            I => \N__32530\
        );

    \I__7511\ : InMux
    port map (
            O => \N__32545\,
            I => \N__32530\
        );

    \I__7510\ : InMux
    port map (
            O => \N__32544\,
            I => \N__32525\
        );

    \I__7509\ : InMux
    port map (
            O => \N__32543\,
            I => \N__32525\
        );

    \I__7508\ : CascadeMux
    port map (
            O => \N__32542\,
            I => \N__32522\
        );

    \I__7507\ : InMux
    port map (
            O => \N__32541\,
            I => \N__32517\
        );

    \I__7506\ : InMux
    port map (
            O => \N__32540\,
            I => \N__32517\
        );

    \I__7505\ : InMux
    port map (
            O => \N__32539\,
            I => \N__32514\
        );

    \I__7504\ : InMux
    port map (
            O => \N__32538\,
            I => \N__32511\
        );

    \I__7503\ : InMux
    port map (
            O => \N__32537\,
            I => \N__32506\
        );

    \I__7502\ : InMux
    port map (
            O => \N__32536\,
            I => \N__32506\
        );

    \I__7501\ : InMux
    port map (
            O => \N__32535\,
            I => \N__32503\
        );

    \I__7500\ : LocalMux
    port map (
            O => \N__32530\,
            I => \N__32500\
        );

    \I__7499\ : LocalMux
    port map (
            O => \N__32525\,
            I => \N__32497\
        );

    \I__7498\ : InMux
    port map (
            O => \N__32522\,
            I => \N__32494\
        );

    \I__7497\ : LocalMux
    port map (
            O => \N__32517\,
            I => \N__32485\
        );

    \I__7496\ : LocalMux
    port map (
            O => \N__32514\,
            I => \N__32485\
        );

    \I__7495\ : LocalMux
    port map (
            O => \N__32511\,
            I => \N__32485\
        );

    \I__7494\ : LocalMux
    port map (
            O => \N__32506\,
            I => \N__32485\
        );

    \I__7493\ : LocalMux
    port map (
            O => \N__32503\,
            I => \N__32482\
        );

    \I__7492\ : Span4Mux_v
    port map (
            O => \N__32500\,
            I => \N__32477\
        );

    \I__7491\ : Span4Mux_v
    port map (
            O => \N__32497\,
            I => \N__32477\
        );

    \I__7490\ : LocalMux
    port map (
            O => \N__32494\,
            I => \N__32474\
        );

    \I__7489\ : Odrv12
    port map (
            O => \N__32485\,
            I => \b2v_inst.un2_valor_max1_THRU_CO\
        );

    \I__7488\ : Odrv12
    port map (
            O => \N__32482\,
            I => \b2v_inst.un2_valor_max1_THRU_CO\
        );

    \I__7487\ : Odrv4
    port map (
            O => \N__32477\,
            I => \b2v_inst.un2_valor_max1_THRU_CO\
        );

    \I__7486\ : Odrv4
    port map (
            O => \N__32474\,
            I => \b2v_inst.un2_valor_max1_THRU_CO\
        );

    \I__7485\ : InMux
    port map (
            O => \N__32465\,
            I => \N__32462\
        );

    \I__7484\ : LocalMux
    port map (
            O => \N__32462\,
            I => \b2v_inst.data_a_escribir_RNO_2Z0Z_3\
        );

    \I__7483\ : CascadeMux
    port map (
            O => \N__32459\,
            I => \N__32455\
        );

    \I__7482\ : CascadeMux
    port map (
            O => \N__32458\,
            I => \N__32452\
        );

    \I__7481\ : InMux
    port map (
            O => \N__32455\,
            I => \N__32449\
        );

    \I__7480\ : InMux
    port map (
            O => \N__32452\,
            I => \N__32445\
        );

    \I__7479\ : LocalMux
    port map (
            O => \N__32449\,
            I => \N__32442\
        );

    \I__7478\ : InMux
    port map (
            O => \N__32448\,
            I => \N__32439\
        );

    \I__7477\ : LocalMux
    port map (
            O => \N__32445\,
            I => \N__32435\
        );

    \I__7476\ : Span4Mux_h
    port map (
            O => \N__32442\,
            I => \N__32429\
        );

    \I__7475\ : LocalMux
    port map (
            O => \N__32439\,
            I => \N__32429\
        );

    \I__7474\ : InMux
    port map (
            O => \N__32438\,
            I => \N__32426\
        );

    \I__7473\ : Span4Mux_v
    port map (
            O => \N__32435\,
            I => \N__32423\
        );

    \I__7472\ : InMux
    port map (
            O => \N__32434\,
            I => \N__32420\
        );

    \I__7471\ : Span4Mux_v
    port map (
            O => \N__32429\,
            I => \N__32417\
        );

    \I__7470\ : LocalMux
    port map (
            O => \N__32426\,
            I => \b2v_inst.reg_ancho_2Z0Z_3\
        );

    \I__7469\ : Odrv4
    port map (
            O => \N__32423\,
            I => \b2v_inst.reg_ancho_2Z0Z_3\
        );

    \I__7468\ : LocalMux
    port map (
            O => \N__32420\,
            I => \b2v_inst.reg_ancho_2Z0Z_3\
        );

    \I__7467\ : Odrv4
    port map (
            O => \N__32417\,
            I => \b2v_inst.reg_ancho_2Z0Z_3\
        );

    \I__7466\ : InMux
    port map (
            O => \N__32408\,
            I => \N__32402\
        );

    \I__7465\ : InMux
    port map (
            O => \N__32407\,
            I => \N__32399\
        );

    \I__7464\ : InMux
    port map (
            O => \N__32406\,
            I => \N__32386\
        );

    \I__7463\ : InMux
    port map (
            O => \N__32405\,
            I => \N__32386\
        );

    \I__7462\ : LocalMux
    port map (
            O => \N__32402\,
            I => \N__32383\
        );

    \I__7461\ : LocalMux
    port map (
            O => \N__32399\,
            I => \N__32380\
        );

    \I__7460\ : InMux
    port map (
            O => \N__32398\,
            I => \N__32377\
        );

    \I__7459\ : InMux
    port map (
            O => \N__32397\,
            I => \N__32374\
        );

    \I__7458\ : InMux
    port map (
            O => \N__32396\,
            I => \N__32369\
        );

    \I__7457\ : InMux
    port map (
            O => \N__32395\,
            I => \N__32369\
        );

    \I__7456\ : InMux
    port map (
            O => \N__32394\,
            I => \N__32366\
        );

    \I__7455\ : InMux
    port map (
            O => \N__32393\,
            I => \N__32359\
        );

    \I__7454\ : InMux
    port map (
            O => \N__32392\,
            I => \N__32359\
        );

    \I__7453\ : InMux
    port map (
            O => \N__32391\,
            I => \N__32359\
        );

    \I__7452\ : LocalMux
    port map (
            O => \N__32386\,
            I => \N__32350\
        );

    \I__7451\ : Span4Mux_v
    port map (
            O => \N__32383\,
            I => \N__32350\
        );

    \I__7450\ : Span4Mux_h
    port map (
            O => \N__32380\,
            I => \N__32350\
        );

    \I__7449\ : LocalMux
    port map (
            O => \N__32377\,
            I => \N__32350\
        );

    \I__7448\ : LocalMux
    port map (
            O => \N__32374\,
            I => \N__32344\
        );

    \I__7447\ : LocalMux
    port map (
            O => \N__32369\,
            I => \N__32344\
        );

    \I__7446\ : LocalMux
    port map (
            O => \N__32366\,
            I => \N__32341\
        );

    \I__7445\ : LocalMux
    port map (
            O => \N__32359\,
            I => \N__32336\
        );

    \I__7444\ : Span4Mux_v
    port map (
            O => \N__32350\,
            I => \N__32336\
        );

    \I__7443\ : InMux
    port map (
            O => \N__32349\,
            I => \N__32333\
        );

    \I__7442\ : Odrv12
    port map (
            O => \N__32344\,
            I => \b2v_inst.un2_valor_max2_THRU_CO\
        );

    \I__7441\ : Odrv4
    port map (
            O => \N__32341\,
            I => \b2v_inst.un2_valor_max2_THRU_CO\
        );

    \I__7440\ : Odrv4
    port map (
            O => \N__32336\,
            I => \b2v_inst.un2_valor_max2_THRU_CO\
        );

    \I__7439\ : LocalMux
    port map (
            O => \N__32333\,
            I => \b2v_inst.un2_valor_max2_THRU_CO\
        );

    \I__7438\ : CascadeMux
    port map (
            O => \N__32324\,
            I => \N__32321\
        );

    \I__7437\ : InMux
    port map (
            O => \N__32321\,
            I => \N__32318\
        );

    \I__7436\ : LocalMux
    port map (
            O => \N__32318\,
            I => \N__32315\
        );

    \I__7435\ : Span4Mux_h
    port map (
            O => \N__32315\,
            I => \N__32312\
        );

    \I__7434\ : Odrv4
    port map (
            O => \N__32312\,
            I => \b2v_inst.N_264\
        );

    \I__7433\ : InMux
    port map (
            O => \N__32309\,
            I => \N__32306\
        );

    \I__7432\ : LocalMux
    port map (
            O => \N__32306\,
            I => \N__32302\
        );

    \I__7431\ : InMux
    port map (
            O => \N__32305\,
            I => \N__32298\
        );

    \I__7430\ : Span4Mux_h
    port map (
            O => \N__32302\,
            I => \N__32295\
        );

    \I__7429\ : InMux
    port map (
            O => \N__32301\,
            I => \N__32292\
        );

    \I__7428\ : LocalMux
    port map (
            O => \N__32298\,
            I => \b2v_inst.reg_ancho_3Z0Z_10\
        );

    \I__7427\ : Odrv4
    port map (
            O => \N__32295\,
            I => \b2v_inst.reg_ancho_3Z0Z_10\
        );

    \I__7426\ : LocalMux
    port map (
            O => \N__32292\,
            I => \b2v_inst.reg_ancho_3Z0Z_10\
        );

    \I__7425\ : InMux
    port map (
            O => \N__32285\,
            I => \N__32279\
        );

    \I__7424\ : InMux
    port map (
            O => \N__32284\,
            I => \N__32276\
        );

    \I__7423\ : InMux
    port map (
            O => \N__32283\,
            I => \N__32273\
        );

    \I__7422\ : InMux
    port map (
            O => \N__32282\,
            I => \N__32270\
        );

    \I__7421\ : LocalMux
    port map (
            O => \N__32279\,
            I => \N__32267\
        );

    \I__7420\ : LocalMux
    port map (
            O => \N__32276\,
            I => \N__32264\
        );

    \I__7419\ : LocalMux
    port map (
            O => \N__32273\,
            I => \N__32261\
        );

    \I__7418\ : LocalMux
    port map (
            O => \N__32270\,
            I => \N__32258\
        );

    \I__7417\ : Span4Mux_h
    port map (
            O => \N__32267\,
            I => \N__32255\
        );

    \I__7416\ : Span4Mux_h
    port map (
            O => \N__32264\,
            I => \N__32252\
        );

    \I__7415\ : Span4Mux_h
    port map (
            O => \N__32261\,
            I => \N__32249\
        );

    \I__7414\ : Span4Mux_h
    port map (
            O => \N__32258\,
            I => \N__32246\
        );

    \I__7413\ : Span4Mux_h
    port map (
            O => \N__32255\,
            I => \N__32241\
        );

    \I__7412\ : Span4Mux_v
    port map (
            O => \N__32252\,
            I => \N__32241\
        );

    \I__7411\ : Span4Mux_v
    port map (
            O => \N__32249\,
            I => \N__32236\
        );

    \I__7410\ : Span4Mux_h
    port map (
            O => \N__32246\,
            I => \N__32236\
        );

    \I__7409\ : Odrv4
    port map (
            O => \N__32241\,
            I => \SYNTHESIZED_WIRE_3_3\
        );

    \I__7408\ : Odrv4
    port map (
            O => \N__32236\,
            I => \SYNTHESIZED_WIRE_3_3\
        );

    \I__7407\ : InMux
    port map (
            O => \N__32231\,
            I => \N__32226\
        );

    \I__7406\ : InMux
    port map (
            O => \N__32230\,
            I => \N__32223\
        );

    \I__7405\ : InMux
    port map (
            O => \N__32229\,
            I => \N__32220\
        );

    \I__7404\ : LocalMux
    port map (
            O => \N__32226\,
            I => \N__32215\
        );

    \I__7403\ : LocalMux
    port map (
            O => \N__32223\,
            I => \N__32215\
        );

    \I__7402\ : LocalMux
    port map (
            O => \N__32220\,
            I => \b2v_inst.reg_ancho_3Z0Z_3\
        );

    \I__7401\ : Odrv4
    port map (
            O => \N__32215\,
            I => \b2v_inst.reg_ancho_3Z0Z_3\
        );

    \I__7400\ : InMux
    port map (
            O => \N__32210\,
            I => \N__32206\
        );

    \I__7399\ : InMux
    port map (
            O => \N__32209\,
            I => \N__32201\
        );

    \I__7398\ : LocalMux
    port map (
            O => \N__32206\,
            I => \N__32198\
        );

    \I__7397\ : InMux
    port map (
            O => \N__32205\,
            I => \N__32195\
        );

    \I__7396\ : InMux
    port map (
            O => \N__32204\,
            I => \N__32192\
        );

    \I__7395\ : LocalMux
    port map (
            O => \N__32201\,
            I => \N__32189\
        );

    \I__7394\ : Span4Mux_h
    port map (
            O => \N__32198\,
            I => \N__32186\
        );

    \I__7393\ : LocalMux
    port map (
            O => \N__32195\,
            I => \N__32183\
        );

    \I__7392\ : LocalMux
    port map (
            O => \N__32192\,
            I => \N__32180\
        );

    \I__7391\ : Span4Mux_v
    port map (
            O => \N__32189\,
            I => \N__32177\
        );

    \I__7390\ : Span4Mux_h
    port map (
            O => \N__32186\,
            I => \N__32172\
        );

    \I__7389\ : Span4Mux_h
    port map (
            O => \N__32183\,
            I => \N__32172\
        );

    \I__7388\ : Span4Mux_v
    port map (
            O => \N__32180\,
            I => \N__32169\
        );

    \I__7387\ : Span4Mux_v
    port map (
            O => \N__32177\,
            I => \N__32166\
        );

    \I__7386\ : Span4Mux_v
    port map (
            O => \N__32172\,
            I => \N__32163\
        );

    \I__7385\ : Span4Mux_h
    port map (
            O => \N__32169\,
            I => \N__32160\
        );

    \I__7384\ : Odrv4
    port map (
            O => \N__32166\,
            I => \SYNTHESIZED_WIRE_3_2\
        );

    \I__7383\ : Odrv4
    port map (
            O => \N__32163\,
            I => \SYNTHESIZED_WIRE_3_2\
        );

    \I__7382\ : Odrv4
    port map (
            O => \N__32160\,
            I => \SYNTHESIZED_WIRE_3_2\
        );

    \I__7381\ : InMux
    port map (
            O => \N__32153\,
            I => \N__32148\
        );

    \I__7380\ : InMux
    port map (
            O => \N__32152\,
            I => \N__32145\
        );

    \I__7379\ : InMux
    port map (
            O => \N__32151\,
            I => \N__32142\
        );

    \I__7378\ : LocalMux
    port map (
            O => \N__32148\,
            I => \N__32139\
        );

    \I__7377\ : LocalMux
    port map (
            O => \N__32145\,
            I => \b2v_inst.reg_ancho_3Z0Z_2\
        );

    \I__7376\ : LocalMux
    port map (
            O => \N__32142\,
            I => \b2v_inst.reg_ancho_3Z0Z_2\
        );

    \I__7375\ : Odrv4
    port map (
            O => \N__32139\,
            I => \b2v_inst.reg_ancho_3Z0Z_2\
        );

    \I__7374\ : InMux
    port map (
            O => \N__32132\,
            I => \N__32128\
        );

    \I__7373\ : InMux
    port map (
            O => \N__32131\,
            I => \N__32125\
        );

    \I__7372\ : LocalMux
    port map (
            O => \N__32128\,
            I => \N__32121\
        );

    \I__7371\ : LocalMux
    port map (
            O => \N__32125\,
            I => \N__32118\
        );

    \I__7370\ : InMux
    port map (
            O => \N__32124\,
            I => \N__32114\
        );

    \I__7369\ : Span4Mux_h
    port map (
            O => \N__32121\,
            I => \N__32111\
        );

    \I__7368\ : Span4Mux_v
    port map (
            O => \N__32118\,
            I => \N__32108\
        );

    \I__7367\ : InMux
    port map (
            O => \N__32117\,
            I => \N__32105\
        );

    \I__7366\ : LocalMux
    port map (
            O => \N__32114\,
            I => \N__32102\
        );

    \I__7365\ : Span4Mux_h
    port map (
            O => \N__32111\,
            I => \N__32099\
        );

    \I__7364\ : Span4Mux_v
    port map (
            O => \N__32108\,
            I => \N__32096\
        );

    \I__7363\ : LocalMux
    port map (
            O => \N__32105\,
            I => \N__32093\
        );

    \I__7362\ : Odrv12
    port map (
            O => \N__32102\,
            I => \SYNTHESIZED_WIRE_3_5\
        );

    \I__7361\ : Odrv4
    port map (
            O => \N__32099\,
            I => \SYNTHESIZED_WIRE_3_5\
        );

    \I__7360\ : Odrv4
    port map (
            O => \N__32096\,
            I => \SYNTHESIZED_WIRE_3_5\
        );

    \I__7359\ : Odrv4
    port map (
            O => \N__32093\,
            I => \SYNTHESIZED_WIRE_3_5\
        );

    \I__7358\ : CascadeMux
    port map (
            O => \N__32084\,
            I => \N__32079\
        );

    \I__7357\ : InMux
    port map (
            O => \N__32083\,
            I => \N__32076\
        );

    \I__7356\ : InMux
    port map (
            O => \N__32082\,
            I => \N__32073\
        );

    \I__7355\ : InMux
    port map (
            O => \N__32079\,
            I => \N__32070\
        );

    \I__7354\ : LocalMux
    port map (
            O => \N__32076\,
            I => \N__32065\
        );

    \I__7353\ : LocalMux
    port map (
            O => \N__32073\,
            I => \N__32065\
        );

    \I__7352\ : LocalMux
    port map (
            O => \N__32070\,
            I => \b2v_inst.reg_ancho_3Z0Z_5\
        );

    \I__7351\ : Odrv4
    port map (
            O => \N__32065\,
            I => \b2v_inst.reg_ancho_3Z0Z_5\
        );

    \I__7350\ : CEMux
    port map (
            O => \N__32060\,
            I => \N__32056\
        );

    \I__7349\ : CEMux
    port map (
            O => \N__32059\,
            I => \N__32053\
        );

    \I__7348\ : LocalMux
    port map (
            O => \N__32056\,
            I => \N__32048\
        );

    \I__7347\ : LocalMux
    port map (
            O => \N__32053\,
            I => \N__32045\
        );

    \I__7346\ : CEMux
    port map (
            O => \N__32052\,
            I => \N__32042\
        );

    \I__7345\ : InMux
    port map (
            O => \N__32051\,
            I => \N__32039\
        );

    \I__7344\ : Span4Mux_v
    port map (
            O => \N__32048\,
            I => \N__32036\
        );

    \I__7343\ : Span4Mux_v
    port map (
            O => \N__32045\,
            I => \N__32033\
        );

    \I__7342\ : LocalMux
    port map (
            O => \N__32042\,
            I => \N__32030\
        );

    \I__7341\ : LocalMux
    port map (
            O => \N__32039\,
            I => \N__32027\
        );

    \I__7340\ : Span4Mux_h
    port map (
            O => \N__32036\,
            I => \N__32021\
        );

    \I__7339\ : Span4Mux_h
    port map (
            O => \N__32033\,
            I => \N__32016\
        );

    \I__7338\ : Span4Mux_h
    port map (
            O => \N__32030\,
            I => \N__32016\
        );

    \I__7337\ : Span4Mux_h
    port map (
            O => \N__32027\,
            I => \N__32013\
        );

    \I__7336\ : InMux
    port map (
            O => \N__32026\,
            I => \N__32008\
        );

    \I__7335\ : InMux
    port map (
            O => \N__32025\,
            I => \N__32008\
        );

    \I__7334\ : InMux
    port map (
            O => \N__32024\,
            I => \N__32005\
        );

    \I__7333\ : Odrv4
    port map (
            O => \N__32021\,
            I => \b2v_inst.stateZ0Z_21\
        );

    \I__7332\ : Odrv4
    port map (
            O => \N__32016\,
            I => \b2v_inst.stateZ0Z_21\
        );

    \I__7331\ : Odrv4
    port map (
            O => \N__32013\,
            I => \b2v_inst.stateZ0Z_21\
        );

    \I__7330\ : LocalMux
    port map (
            O => \N__32008\,
            I => \b2v_inst.stateZ0Z_21\
        );

    \I__7329\ : LocalMux
    port map (
            O => \N__32005\,
            I => \b2v_inst.stateZ0Z_21\
        );

    \I__7328\ : InMux
    port map (
            O => \N__31994\,
            I => \N__31990\
        );

    \I__7327\ : InMux
    port map (
            O => \N__31993\,
            I => \N__31986\
        );

    \I__7326\ : LocalMux
    port map (
            O => \N__31990\,
            I => \N__31982\
        );

    \I__7325\ : InMux
    port map (
            O => \N__31989\,
            I => \N__31979\
        );

    \I__7324\ : LocalMux
    port map (
            O => \N__31986\,
            I => \N__31976\
        );

    \I__7323\ : InMux
    port map (
            O => \N__31985\,
            I => \N__31973\
        );

    \I__7322\ : Span4Mux_h
    port map (
            O => \N__31982\,
            I => \N__31966\
        );

    \I__7321\ : LocalMux
    port map (
            O => \N__31979\,
            I => \N__31966\
        );

    \I__7320\ : Span4Mux_v
    port map (
            O => \N__31976\,
            I => \N__31966\
        );

    \I__7319\ : LocalMux
    port map (
            O => \N__31973\,
            I => \N__31963\
        );

    \I__7318\ : Span4Mux_h
    port map (
            O => \N__31966\,
            I => \N__31958\
        );

    \I__7317\ : Span4Mux_h
    port map (
            O => \N__31963\,
            I => \N__31958\
        );

    \I__7316\ : Odrv4
    port map (
            O => \N__31958\,
            I => \SYNTHESIZED_WIRE_3_9\
        );

    \I__7315\ : InMux
    port map (
            O => \N__31955\,
            I => \N__31951\
        );

    \I__7314\ : InMux
    port map (
            O => \N__31954\,
            I => \N__31947\
        );

    \I__7313\ : LocalMux
    port map (
            O => \N__31951\,
            I => \N__31943\
        );

    \I__7312\ : InMux
    port map (
            O => \N__31950\,
            I => \N__31940\
        );

    \I__7311\ : LocalMux
    port map (
            O => \N__31947\,
            I => \N__31937\
        );

    \I__7310\ : InMux
    port map (
            O => \N__31946\,
            I => \N__31934\
        );

    \I__7309\ : Span4Mux_h
    port map (
            O => \N__31943\,
            I => \N__31931\
        );

    \I__7308\ : LocalMux
    port map (
            O => \N__31940\,
            I => \N__31928\
        );

    \I__7307\ : Odrv12
    port map (
            O => \N__31937\,
            I => \b2v_inst.reg_anteriorZ0Z_9\
        );

    \I__7306\ : LocalMux
    port map (
            O => \N__31934\,
            I => \b2v_inst.reg_anteriorZ0Z_9\
        );

    \I__7305\ : Odrv4
    port map (
            O => \N__31931\,
            I => \b2v_inst.reg_anteriorZ0Z_9\
        );

    \I__7304\ : Odrv4
    port map (
            O => \N__31928\,
            I => \b2v_inst.reg_anteriorZ0Z_9\
        );

    \I__7303\ : InMux
    port map (
            O => \N__31919\,
            I => \N__31914\
        );

    \I__7302\ : InMux
    port map (
            O => \N__31918\,
            I => \N__31909\
        );

    \I__7301\ : InMux
    port map (
            O => \N__31917\,
            I => \N__31909\
        );

    \I__7300\ : LocalMux
    port map (
            O => \N__31914\,
            I => \N__31889\
        );

    \I__7299\ : LocalMux
    port map (
            O => \N__31909\,
            I => \N__31889\
        );

    \I__7298\ : InMux
    port map (
            O => \N__31908\,
            I => \N__31876\
        );

    \I__7297\ : InMux
    port map (
            O => \N__31907\,
            I => \N__31876\
        );

    \I__7296\ : InMux
    port map (
            O => \N__31906\,
            I => \N__31876\
        );

    \I__7295\ : InMux
    port map (
            O => \N__31905\,
            I => \N__31876\
        );

    \I__7294\ : InMux
    port map (
            O => \N__31904\,
            I => \N__31876\
        );

    \I__7293\ : InMux
    port map (
            O => \N__31903\,
            I => \N__31876\
        );

    \I__7292\ : InMux
    port map (
            O => \N__31902\,
            I => \N__31873\
        );

    \I__7291\ : InMux
    port map (
            O => \N__31901\,
            I => \N__31864\
        );

    \I__7290\ : InMux
    port map (
            O => \N__31900\,
            I => \N__31864\
        );

    \I__7289\ : InMux
    port map (
            O => \N__31899\,
            I => \N__31864\
        );

    \I__7288\ : InMux
    port map (
            O => \N__31898\,
            I => \N__31864\
        );

    \I__7287\ : InMux
    port map (
            O => \N__31897\,
            I => \N__31859\
        );

    \I__7286\ : InMux
    port map (
            O => \N__31896\,
            I => \N__31859\
        );

    \I__7285\ : InMux
    port map (
            O => \N__31895\,
            I => \N__31853\
        );

    \I__7284\ : InMux
    port map (
            O => \N__31894\,
            I => \N__31853\
        );

    \I__7283\ : Span4Mux_v
    port map (
            O => \N__31889\,
            I => \N__31848\
        );

    \I__7282\ : LocalMux
    port map (
            O => \N__31876\,
            I => \N__31848\
        );

    \I__7281\ : LocalMux
    port map (
            O => \N__31873\,
            I => \N__31843\
        );

    \I__7280\ : LocalMux
    port map (
            O => \N__31864\,
            I => \N__31843\
        );

    \I__7279\ : LocalMux
    port map (
            O => \N__31859\,
            I => \N__31840\
        );

    \I__7278\ : InMux
    port map (
            O => \N__31858\,
            I => \N__31837\
        );

    \I__7277\ : LocalMux
    port map (
            O => \N__31853\,
            I => \N__31834\
        );

    \I__7276\ : Span4Mux_h
    port map (
            O => \N__31848\,
            I => \N__31828\
        );

    \I__7275\ : Span4Mux_v
    port map (
            O => \N__31843\,
            I => \N__31825\
        );

    \I__7274\ : Span4Mux_h
    port map (
            O => \N__31840\,
            I => \N__31820\
        );

    \I__7273\ : LocalMux
    port map (
            O => \N__31837\,
            I => \N__31820\
        );

    \I__7272\ : Span4Mux_v
    port map (
            O => \N__31834\,
            I => \N__31817\
        );

    \I__7271\ : InMux
    port map (
            O => \N__31833\,
            I => \N__31814\
        );

    \I__7270\ : InMux
    port map (
            O => \N__31832\,
            I => \N__31809\
        );

    \I__7269\ : InMux
    port map (
            O => \N__31831\,
            I => \N__31809\
        );

    \I__7268\ : Span4Mux_v
    port map (
            O => \N__31828\,
            I => \N__31802\
        );

    \I__7267\ : Span4Mux_h
    port map (
            O => \N__31825\,
            I => \N__31802\
        );

    \I__7266\ : Span4Mux_h
    port map (
            O => \N__31820\,
            I => \N__31802\
        );

    \I__7265\ : Sp12to4
    port map (
            O => \N__31817\,
            I => \N__31795\
        );

    \I__7264\ : LocalMux
    port map (
            O => \N__31814\,
            I => \N__31795\
        );

    \I__7263\ : LocalMux
    port map (
            O => \N__31809\,
            I => \N__31795\
        );

    \I__7262\ : Span4Mux_h
    port map (
            O => \N__31802\,
            I => \N__31792\
        );

    \I__7261\ : Span12Mux_h
    port map (
            O => \N__31795\,
            I => \N__31789\
        );

    \I__7260\ : Span4Mux_h
    port map (
            O => \N__31792\,
            I => \N__31786\
        );

    \I__7259\ : Odrv12
    port map (
            O => \N__31789\,
            I => \b2v_inst.ignorar_anteriorZ0\
        );

    \I__7258\ : Odrv4
    port map (
            O => \N__31786\,
            I => \b2v_inst.ignorar_anteriorZ0\
        );

    \I__7257\ : InMux
    port map (
            O => \N__31781\,
            I => \N__31777\
        );

    \I__7256\ : InMux
    port map (
            O => \N__31780\,
            I => \N__31773\
        );

    \I__7255\ : LocalMux
    port map (
            O => \N__31777\,
            I => \N__31769\
        );

    \I__7254\ : InMux
    port map (
            O => \N__31776\,
            I => \N__31766\
        );

    \I__7253\ : LocalMux
    port map (
            O => \N__31773\,
            I => \N__31763\
        );

    \I__7252\ : InMux
    port map (
            O => \N__31772\,
            I => \N__31760\
        );

    \I__7251\ : Span4Mux_v
    port map (
            O => \N__31769\,
            I => \N__31757\
        );

    \I__7250\ : LocalMux
    port map (
            O => \N__31766\,
            I => \N__31754\
        );

    \I__7249\ : Span4Mux_h
    port map (
            O => \N__31763\,
            I => \N__31751\
        );

    \I__7248\ : LocalMux
    port map (
            O => \N__31760\,
            I => \N__31748\
        );

    \I__7247\ : Span4Mux_h
    port map (
            O => \N__31757\,
            I => \N__31745\
        );

    \I__7246\ : Span4Mux_h
    port map (
            O => \N__31754\,
            I => \N__31742\
        );

    \I__7245\ : Span4Mux_v
    port map (
            O => \N__31751\,
            I => \N__31737\
        );

    \I__7244\ : Span4Mux_h
    port map (
            O => \N__31748\,
            I => \N__31737\
        );

    \I__7243\ : Odrv4
    port map (
            O => \N__31745\,
            I => \SYNTHESIZED_WIRE_3_10\
        );

    \I__7242\ : Odrv4
    port map (
            O => \N__31742\,
            I => \SYNTHESIZED_WIRE_3_10\
        );

    \I__7241\ : Odrv4
    port map (
            O => \N__31737\,
            I => \SYNTHESIZED_WIRE_3_10\
        );

    \I__7240\ : CascadeMux
    port map (
            O => \N__31730\,
            I => \N__31727\
        );

    \I__7239\ : InMux
    port map (
            O => \N__31727\,
            I => \N__31723\
        );

    \I__7238\ : InMux
    port map (
            O => \N__31726\,
            I => \N__31720\
        );

    \I__7237\ : LocalMux
    port map (
            O => \N__31723\,
            I => \N__31715\
        );

    \I__7236\ : LocalMux
    port map (
            O => \N__31720\,
            I => \N__31712\
        );

    \I__7235\ : InMux
    port map (
            O => \N__31719\,
            I => \N__31709\
        );

    \I__7234\ : InMux
    port map (
            O => \N__31718\,
            I => \N__31706\
        );

    \I__7233\ : Span4Mux_v
    port map (
            O => \N__31715\,
            I => \N__31703\
        );

    \I__7232\ : Span4Mux_h
    port map (
            O => \N__31712\,
            I => \N__31700\
        );

    \I__7231\ : LocalMux
    port map (
            O => \N__31709\,
            I => \N__31697\
        );

    \I__7230\ : LocalMux
    port map (
            O => \N__31706\,
            I => \b2v_inst.reg_anteriorZ0Z_10\
        );

    \I__7229\ : Odrv4
    port map (
            O => \N__31703\,
            I => \b2v_inst.reg_anteriorZ0Z_10\
        );

    \I__7228\ : Odrv4
    port map (
            O => \N__31700\,
            I => \b2v_inst.reg_anteriorZ0Z_10\
        );

    \I__7227\ : Odrv4
    port map (
            O => \N__31697\,
            I => \b2v_inst.reg_anteriorZ0Z_10\
        );

    \I__7226\ : CEMux
    port map (
            O => \N__31688\,
            I => \N__31683\
        );

    \I__7225\ : CEMux
    port map (
            O => \N__31687\,
            I => \N__31680\
        );

    \I__7224\ : CEMux
    port map (
            O => \N__31686\,
            I => \N__31677\
        );

    \I__7223\ : LocalMux
    port map (
            O => \N__31683\,
            I => \N__31674\
        );

    \I__7222\ : LocalMux
    port map (
            O => \N__31680\,
            I => \N__31668\
        );

    \I__7221\ : LocalMux
    port map (
            O => \N__31677\,
            I => \N__31663\
        );

    \I__7220\ : Span4Mux_v
    port map (
            O => \N__31674\,
            I => \N__31660\
        );

    \I__7219\ : CEMux
    port map (
            O => \N__31673\,
            I => \N__31657\
        );

    \I__7218\ : CEMux
    port map (
            O => \N__31672\,
            I => \N__31654\
        );

    \I__7217\ : CEMux
    port map (
            O => \N__31671\,
            I => \N__31651\
        );

    \I__7216\ : Span4Mux_h
    port map (
            O => \N__31668\,
            I => \N__31648\
        );

    \I__7215\ : CascadeMux
    port map (
            O => \N__31667\,
            I => \N__31645\
        );

    \I__7214\ : InMux
    port map (
            O => \N__31666\,
            I => \N__31642\
        );

    \I__7213\ : Span4Mux_v
    port map (
            O => \N__31663\,
            I => \N__31639\
        );

    \I__7212\ : Span4Mux_v
    port map (
            O => \N__31660\,
            I => \N__31634\
        );

    \I__7211\ : LocalMux
    port map (
            O => \N__31657\,
            I => \N__31634\
        );

    \I__7210\ : LocalMux
    port map (
            O => \N__31654\,
            I => \N__31631\
        );

    \I__7209\ : LocalMux
    port map (
            O => \N__31651\,
            I => \N__31626\
        );

    \I__7208\ : Span4Mux_v
    port map (
            O => \N__31648\,
            I => \N__31626\
        );

    \I__7207\ : InMux
    port map (
            O => \N__31645\,
            I => \N__31623\
        );

    \I__7206\ : LocalMux
    port map (
            O => \N__31642\,
            I => \N__31619\
        );

    \I__7205\ : Sp12to4
    port map (
            O => \N__31639\,
            I => \N__31614\
        );

    \I__7204\ : Sp12to4
    port map (
            O => \N__31634\,
            I => \N__31614\
        );

    \I__7203\ : Span4Mux_v
    port map (
            O => \N__31631\,
            I => \N__31610\
        );

    \I__7202\ : Span4Mux_h
    port map (
            O => \N__31626\,
            I => \N__31605\
        );

    \I__7201\ : LocalMux
    port map (
            O => \N__31623\,
            I => \N__31605\
        );

    \I__7200\ : InMux
    port map (
            O => \N__31622\,
            I => \N__31601\
        );

    \I__7199\ : Span4Mux_h
    port map (
            O => \N__31619\,
            I => \N__31598\
        );

    \I__7198\ : Span12Mux_h
    port map (
            O => \N__31614\,
            I => \N__31595\
        );

    \I__7197\ : InMux
    port map (
            O => \N__31613\,
            I => \N__31592\
        );

    \I__7196\ : Span4Mux_h
    port map (
            O => \N__31610\,
            I => \N__31587\
        );

    \I__7195\ : Span4Mux_v
    port map (
            O => \N__31605\,
            I => \N__31587\
        );

    \I__7194\ : InMux
    port map (
            O => \N__31604\,
            I => \N__31584\
        );

    \I__7193\ : LocalMux
    port map (
            O => \N__31601\,
            I => \b2v_inst.stateZ0Z_27\
        );

    \I__7192\ : Odrv4
    port map (
            O => \N__31598\,
            I => \b2v_inst.stateZ0Z_27\
        );

    \I__7191\ : Odrv12
    port map (
            O => \N__31595\,
            I => \b2v_inst.stateZ0Z_27\
        );

    \I__7190\ : LocalMux
    port map (
            O => \N__31592\,
            I => \b2v_inst.stateZ0Z_27\
        );

    \I__7189\ : Odrv4
    port map (
            O => \N__31587\,
            I => \b2v_inst.stateZ0Z_27\
        );

    \I__7188\ : LocalMux
    port map (
            O => \N__31584\,
            I => \b2v_inst.stateZ0Z_27\
        );

    \I__7187\ : InMux
    port map (
            O => \N__31571\,
            I => \N__31567\
        );

    \I__7186\ : InMux
    port map (
            O => \N__31570\,
            I => \N__31564\
        );

    \I__7185\ : LocalMux
    port map (
            O => \N__31567\,
            I => \N__31559\
        );

    \I__7184\ : LocalMux
    port map (
            O => \N__31564\,
            I => \N__31556\
        );

    \I__7183\ : InMux
    port map (
            O => \N__31563\,
            I => \N__31553\
        );

    \I__7182\ : InMux
    port map (
            O => \N__31562\,
            I => \N__31550\
        );

    \I__7181\ : Span4Mux_h
    port map (
            O => \N__31559\,
            I => \N__31543\
        );

    \I__7180\ : Span4Mux_v
    port map (
            O => \N__31556\,
            I => \N__31543\
        );

    \I__7179\ : LocalMux
    port map (
            O => \N__31553\,
            I => \N__31543\
        );

    \I__7178\ : LocalMux
    port map (
            O => \N__31550\,
            I => \N__31540\
        );

    \I__7177\ : Span4Mux_h
    port map (
            O => \N__31543\,
            I => \N__31537\
        );

    \I__7176\ : Span4Mux_h
    port map (
            O => \N__31540\,
            I => \N__31534\
        );

    \I__7175\ : Odrv4
    port map (
            O => \N__31537\,
            I => \SYNTHESIZED_WIRE_3_6\
        );

    \I__7174\ : Odrv4
    port map (
            O => \N__31534\,
            I => \SYNTHESIZED_WIRE_3_6\
        );

    \I__7173\ : CascadeMux
    port map (
            O => \N__31529\,
            I => \N__31526\
        );

    \I__7172\ : InMux
    port map (
            O => \N__31526\,
            I => \N__31522\
        );

    \I__7171\ : InMux
    port map (
            O => \N__31525\,
            I => \N__31519\
        );

    \I__7170\ : LocalMux
    port map (
            O => \N__31522\,
            I => \N__31515\
        );

    \I__7169\ : LocalMux
    port map (
            O => \N__31519\,
            I => \N__31511\
        );

    \I__7168\ : InMux
    port map (
            O => \N__31518\,
            I => \N__31508\
        );

    \I__7167\ : Span4Mux_h
    port map (
            O => \N__31515\,
            I => \N__31505\
        );

    \I__7166\ : InMux
    port map (
            O => \N__31514\,
            I => \N__31502\
        );

    \I__7165\ : Span4Mux_v
    port map (
            O => \N__31511\,
            I => \N__31499\
        );

    \I__7164\ : LocalMux
    port map (
            O => \N__31508\,
            I => \b2v_inst.reg_anteriorZ0Z_6\
        );

    \I__7163\ : Odrv4
    port map (
            O => \N__31505\,
            I => \b2v_inst.reg_anteriorZ0Z_6\
        );

    \I__7162\ : LocalMux
    port map (
            O => \N__31502\,
            I => \b2v_inst.reg_anteriorZ0Z_6\
        );

    \I__7161\ : Odrv4
    port map (
            O => \N__31499\,
            I => \b2v_inst.reg_anteriorZ0Z_6\
        );

    \I__7160\ : InMux
    port map (
            O => \N__31490\,
            I => \N__31484\
        );

    \I__7159\ : InMux
    port map (
            O => \N__31489\,
            I => \N__31480\
        );

    \I__7158\ : CascadeMux
    port map (
            O => \N__31488\,
            I => \N__31477\
        );

    \I__7157\ : InMux
    port map (
            O => \N__31487\,
            I => \N__31474\
        );

    \I__7156\ : LocalMux
    port map (
            O => \N__31484\,
            I => \N__31471\
        );

    \I__7155\ : InMux
    port map (
            O => \N__31483\,
            I => \N__31468\
        );

    \I__7154\ : LocalMux
    port map (
            O => \N__31480\,
            I => \N__31465\
        );

    \I__7153\ : InMux
    port map (
            O => \N__31477\,
            I => \N__31462\
        );

    \I__7152\ : LocalMux
    port map (
            O => \N__31474\,
            I => \N__31459\
        );

    \I__7151\ : Span4Mux_h
    port map (
            O => \N__31471\,
            I => \N__31450\
        );

    \I__7150\ : LocalMux
    port map (
            O => \N__31468\,
            I => \N__31450\
        );

    \I__7149\ : Span4Mux_v
    port map (
            O => \N__31465\,
            I => \N__31450\
        );

    \I__7148\ : LocalMux
    port map (
            O => \N__31462\,
            I => \N__31450\
        );

    \I__7147\ : Span4Mux_h
    port map (
            O => \N__31459\,
            I => \N__31445\
        );

    \I__7146\ : Span4Mux_v
    port map (
            O => \N__31450\,
            I => \N__31445\
        );

    \I__7145\ : Odrv4
    port map (
            O => \N__31445\,
            I => \b2v_inst.reg_ancho_2Z0Z_10\
        );

    \I__7144\ : InMux
    port map (
            O => \N__31442\,
            I => \N__31439\
        );

    \I__7143\ : LocalMux
    port map (
            O => \N__31439\,
            I => \N__31435\
        );

    \I__7142\ : InMux
    port map (
            O => \N__31438\,
            I => \N__31432\
        );

    \I__7141\ : Span4Mux_v
    port map (
            O => \N__31435\,
            I => \N__31427\
        );

    \I__7140\ : LocalMux
    port map (
            O => \N__31432\,
            I => \N__31427\
        );

    \I__7139\ : Span4Mux_h
    port map (
            O => \N__31427\,
            I => \N__31423\
        );

    \I__7138\ : InMux
    port map (
            O => \N__31426\,
            I => \N__31420\
        );

    \I__7137\ : Odrv4
    port map (
            O => \N__31423\,
            I => \b2v_inst.reg_ancho_3Z0Z_4\
        );

    \I__7136\ : LocalMux
    port map (
            O => \N__31420\,
            I => \b2v_inst.reg_ancho_3Z0Z_4\
        );

    \I__7135\ : InMux
    port map (
            O => \N__31415\,
            I => \N__31412\
        );

    \I__7134\ : LocalMux
    port map (
            O => \N__31412\,
            I => \N__31409\
        );

    \I__7133\ : Span4Mux_v
    port map (
            O => \N__31409\,
            I => \N__31406\
        );

    \I__7132\ : Span4Mux_h
    port map (
            O => \N__31406\,
            I => \N__31403\
        );

    \I__7131\ : Odrv4
    port map (
            O => \N__31403\,
            I => \b2v_inst.data_a_escribir11_3_and\
        );

    \I__7130\ : InMux
    port map (
            O => \N__31400\,
            I => \N__31397\
        );

    \I__7129\ : LocalMux
    port map (
            O => \N__31397\,
            I => \N__31391\
        );

    \I__7128\ : InMux
    port map (
            O => \N__31396\,
            I => \N__31388\
        );

    \I__7127\ : InMux
    port map (
            O => \N__31395\,
            I => \N__31385\
        );

    \I__7126\ : InMux
    port map (
            O => \N__31394\,
            I => \N__31382\
        );

    \I__7125\ : Span4Mux_v
    port map (
            O => \N__31391\,
            I => \N__31377\
        );

    \I__7124\ : LocalMux
    port map (
            O => \N__31388\,
            I => \N__31377\
        );

    \I__7123\ : LocalMux
    port map (
            O => \N__31385\,
            I => \N__31374\
        );

    \I__7122\ : LocalMux
    port map (
            O => \N__31382\,
            I => \N__31371\
        );

    \I__7121\ : Span4Mux_v
    port map (
            O => \N__31377\,
            I => \N__31368\
        );

    \I__7120\ : Span4Mux_v
    port map (
            O => \N__31374\,
            I => \N__31363\
        );

    \I__7119\ : Span4Mux_h
    port map (
            O => \N__31371\,
            I => \N__31363\
        );

    \I__7118\ : Span4Mux_h
    port map (
            O => \N__31368\,
            I => \N__31360\
        );

    \I__7117\ : Span4Mux_v
    port map (
            O => \N__31363\,
            I => \N__31357\
        );

    \I__7116\ : Odrv4
    port map (
            O => \N__31360\,
            I => \SYNTHESIZED_WIRE_3_1\
        );

    \I__7115\ : Odrv4
    port map (
            O => \N__31357\,
            I => \SYNTHESIZED_WIRE_3_1\
        );

    \I__7114\ : CascadeMux
    port map (
            O => \N__31352\,
            I => \N__31347\
        );

    \I__7113\ : InMux
    port map (
            O => \N__31351\,
            I => \N__31343\
        );

    \I__7112\ : InMux
    port map (
            O => \N__31350\,
            I => \N__31340\
        );

    \I__7111\ : InMux
    port map (
            O => \N__31347\,
            I => \N__31337\
        );

    \I__7110\ : InMux
    port map (
            O => \N__31346\,
            I => \N__31334\
        );

    \I__7109\ : LocalMux
    port map (
            O => \N__31343\,
            I => \N__31331\
        );

    \I__7108\ : LocalMux
    port map (
            O => \N__31340\,
            I => \N__31327\
        );

    \I__7107\ : LocalMux
    port map (
            O => \N__31337\,
            I => \N__31322\
        );

    \I__7106\ : LocalMux
    port map (
            O => \N__31334\,
            I => \N__31322\
        );

    \I__7105\ : Span4Mux_h
    port map (
            O => \N__31331\,
            I => \N__31319\
        );

    \I__7104\ : InMux
    port map (
            O => \N__31330\,
            I => \N__31316\
        );

    \I__7103\ : Span4Mux_v
    port map (
            O => \N__31327\,
            I => \N__31311\
        );

    \I__7102\ : Span4Mux_v
    port map (
            O => \N__31322\,
            I => \N__31311\
        );

    \I__7101\ : Odrv4
    port map (
            O => \N__31319\,
            I => \b2v_inst.reg_ancho_2Z0Z_1\
        );

    \I__7100\ : LocalMux
    port map (
            O => \N__31316\,
            I => \b2v_inst.reg_ancho_2Z0Z_1\
        );

    \I__7099\ : Odrv4
    port map (
            O => \N__31311\,
            I => \b2v_inst.reg_ancho_2Z0Z_1\
        );

    \I__7098\ : CascadeMux
    port map (
            O => \N__31304\,
            I => \N__31301\
        );

    \I__7097\ : InMux
    port map (
            O => \N__31301\,
            I => \N__31296\
        );

    \I__7096\ : InMux
    port map (
            O => \N__31300\,
            I => \N__31293\
        );

    \I__7095\ : InMux
    port map (
            O => \N__31299\,
            I => \N__31290\
        );

    \I__7094\ : LocalMux
    port map (
            O => \N__31296\,
            I => \N__31287\
        );

    \I__7093\ : LocalMux
    port map (
            O => \N__31293\,
            I => \N__31284\
        );

    \I__7092\ : LocalMux
    port map (
            O => \N__31290\,
            I => \N__31279\
        );

    \I__7091\ : Span4Mux_h
    port map (
            O => \N__31287\,
            I => \N__31276\
        );

    \I__7090\ : Span4Mux_h
    port map (
            O => \N__31284\,
            I => \N__31273\
        );

    \I__7089\ : InMux
    port map (
            O => \N__31283\,
            I => \N__31268\
        );

    \I__7088\ : InMux
    port map (
            O => \N__31282\,
            I => \N__31268\
        );

    \I__7087\ : Span4Mux_h
    port map (
            O => \N__31279\,
            I => \N__31265\
        );

    \I__7086\ : Odrv4
    port map (
            O => \N__31276\,
            I => \b2v_inst.reg_ancho_2Z0Z_2\
        );

    \I__7085\ : Odrv4
    port map (
            O => \N__31273\,
            I => \b2v_inst.reg_ancho_2Z0Z_2\
        );

    \I__7084\ : LocalMux
    port map (
            O => \N__31268\,
            I => \b2v_inst.reg_ancho_2Z0Z_2\
        );

    \I__7083\ : Odrv4
    port map (
            O => \N__31265\,
            I => \b2v_inst.reg_ancho_2Z0Z_2\
        );

    \I__7082\ : InMux
    port map (
            O => \N__31256\,
            I => \N__31252\
        );

    \I__7081\ : InMux
    port map (
            O => \N__31255\,
            I => \N__31249\
        );

    \I__7080\ : LocalMux
    port map (
            O => \N__31252\,
            I => \N__31246\
        );

    \I__7079\ : LocalMux
    port map (
            O => \N__31249\,
            I => \N__31242\
        );

    \I__7078\ : Span4Mux_v
    port map (
            O => \N__31246\,
            I => \N__31238\
        );

    \I__7077\ : InMux
    port map (
            O => \N__31245\,
            I => \N__31235\
        );

    \I__7076\ : Span4Mux_v
    port map (
            O => \N__31242\,
            I => \N__31232\
        );

    \I__7075\ : InMux
    port map (
            O => \N__31241\,
            I => \N__31229\
        );

    \I__7074\ : Span4Mux_h
    port map (
            O => \N__31238\,
            I => \N__31224\
        );

    \I__7073\ : LocalMux
    port map (
            O => \N__31235\,
            I => \N__31224\
        );

    \I__7072\ : Span4Mux_h
    port map (
            O => \N__31232\,
            I => \N__31220\
        );

    \I__7071\ : LocalMux
    port map (
            O => \N__31229\,
            I => \N__31217\
        );

    \I__7070\ : Span4Mux_h
    port map (
            O => \N__31224\,
            I => \N__31214\
        );

    \I__7069\ : InMux
    port map (
            O => \N__31223\,
            I => \N__31211\
        );

    \I__7068\ : Odrv4
    port map (
            O => \N__31220\,
            I => \b2v_inst.reg_ancho_1Z0Z_2\
        );

    \I__7067\ : Odrv12
    port map (
            O => \N__31217\,
            I => \b2v_inst.reg_ancho_1Z0Z_2\
        );

    \I__7066\ : Odrv4
    port map (
            O => \N__31214\,
            I => \b2v_inst.reg_ancho_1Z0Z_2\
        );

    \I__7065\ : LocalMux
    port map (
            O => \N__31211\,
            I => \b2v_inst.reg_ancho_1Z0Z_2\
        );

    \I__7064\ : InMux
    port map (
            O => \N__31202\,
            I => \N__31199\
        );

    \I__7063\ : LocalMux
    port map (
            O => \N__31199\,
            I => \N__31196\
        );

    \I__7062\ : Span4Mux_h
    port map (
            O => \N__31196\,
            I => \N__31192\
        );

    \I__7061\ : InMux
    port map (
            O => \N__31195\,
            I => \N__31189\
        );

    \I__7060\ : Odrv4
    port map (
            O => \N__31192\,
            I => \b2v_inst.eventosZ0Z_2\
        );

    \I__7059\ : LocalMux
    port map (
            O => \N__31189\,
            I => \b2v_inst.eventosZ0Z_2\
        );

    \I__7058\ : CascadeMux
    port map (
            O => \N__31184\,
            I => \b2v_inst.data_a_escribir_RNO_2Z0Z_2_cascade_\
        );

    \I__7057\ : InMux
    port map (
            O => \N__31181\,
            I => \N__31161\
        );

    \I__7056\ : InMux
    port map (
            O => \N__31180\,
            I => \N__31158\
        );

    \I__7055\ : InMux
    port map (
            O => \N__31179\,
            I => \N__31151\
        );

    \I__7054\ : InMux
    port map (
            O => \N__31178\,
            I => \N__31151\
        );

    \I__7053\ : InMux
    port map (
            O => \N__31177\,
            I => \N__31151\
        );

    \I__7052\ : InMux
    port map (
            O => \N__31176\,
            I => \N__31148\
        );

    \I__7051\ : InMux
    port map (
            O => \N__31175\,
            I => \N__31139\
        );

    \I__7050\ : InMux
    port map (
            O => \N__31174\,
            I => \N__31139\
        );

    \I__7049\ : InMux
    port map (
            O => \N__31173\,
            I => \N__31139\
        );

    \I__7048\ : InMux
    port map (
            O => \N__31172\,
            I => \N__31139\
        );

    \I__7047\ : InMux
    port map (
            O => \N__31171\,
            I => \N__31130\
        );

    \I__7046\ : InMux
    port map (
            O => \N__31170\,
            I => \N__31130\
        );

    \I__7045\ : InMux
    port map (
            O => \N__31169\,
            I => \N__31130\
        );

    \I__7044\ : InMux
    port map (
            O => \N__31168\,
            I => \N__31130\
        );

    \I__7043\ : InMux
    port map (
            O => \N__31167\,
            I => \N__31120\
        );

    \I__7042\ : InMux
    port map (
            O => \N__31166\,
            I => \N__31120\
        );

    \I__7041\ : InMux
    port map (
            O => \N__31165\,
            I => \N__31120\
        );

    \I__7040\ : InMux
    port map (
            O => \N__31164\,
            I => \N__31120\
        );

    \I__7039\ : LocalMux
    port map (
            O => \N__31161\,
            I => \N__31105\
        );

    \I__7038\ : LocalMux
    port map (
            O => \N__31158\,
            I => \N__31105\
        );

    \I__7037\ : LocalMux
    port map (
            O => \N__31151\,
            I => \N__31096\
        );

    \I__7036\ : LocalMux
    port map (
            O => \N__31148\,
            I => \N__31096\
        );

    \I__7035\ : LocalMux
    port map (
            O => \N__31139\,
            I => \N__31096\
        );

    \I__7034\ : LocalMux
    port map (
            O => \N__31130\,
            I => \N__31096\
        );

    \I__7033\ : InMux
    port map (
            O => \N__31129\,
            I => \N__31093\
        );

    \I__7032\ : LocalMux
    port map (
            O => \N__31120\,
            I => \N__31090\
        );

    \I__7031\ : InMux
    port map (
            O => \N__31119\,
            I => \N__31077\
        );

    \I__7030\ : InMux
    port map (
            O => \N__31118\,
            I => \N__31077\
        );

    \I__7029\ : InMux
    port map (
            O => \N__31117\,
            I => \N__31077\
        );

    \I__7028\ : InMux
    port map (
            O => \N__31116\,
            I => \N__31077\
        );

    \I__7027\ : InMux
    port map (
            O => \N__31115\,
            I => \N__31077\
        );

    \I__7026\ : InMux
    port map (
            O => \N__31114\,
            I => \N__31077\
        );

    \I__7025\ : InMux
    port map (
            O => \N__31113\,
            I => \N__31068\
        );

    \I__7024\ : InMux
    port map (
            O => \N__31112\,
            I => \N__31068\
        );

    \I__7023\ : InMux
    port map (
            O => \N__31111\,
            I => \N__31068\
        );

    \I__7022\ : InMux
    port map (
            O => \N__31110\,
            I => \N__31068\
        );

    \I__7021\ : Span4Mux_h
    port map (
            O => \N__31105\,
            I => \N__31061\
        );

    \I__7020\ : Span4Mux_v
    port map (
            O => \N__31096\,
            I => \N__31061\
        );

    \I__7019\ : LocalMux
    port map (
            O => \N__31093\,
            I => \N__31061\
        );

    \I__7018\ : Span4Mux_h
    port map (
            O => \N__31090\,
            I => \N__31056\
        );

    \I__7017\ : LocalMux
    port map (
            O => \N__31077\,
            I => \N__31056\
        );

    \I__7016\ : LocalMux
    port map (
            O => \N__31068\,
            I => \b2v_inst.data_a_escribir12_THRU_CO\
        );

    \I__7015\ : Odrv4
    port map (
            O => \N__31061\,
            I => \b2v_inst.data_a_escribir12_THRU_CO\
        );

    \I__7014\ : Odrv4
    port map (
            O => \N__31056\,
            I => \b2v_inst.data_a_escribir12_THRU_CO\
        );

    \I__7013\ : InMux
    port map (
            O => \N__31049\,
            I => \N__31046\
        );

    \I__7012\ : LocalMux
    port map (
            O => \N__31046\,
            I => \b2v_inst.un1_reg_anterior_0_i_1_2\
        );

    \I__7011\ : InMux
    port map (
            O => \N__31043\,
            I => \N__31038\
        );

    \I__7010\ : CascadeMux
    port map (
            O => \N__31042\,
            I => \N__31034\
        );

    \I__7009\ : InMux
    port map (
            O => \N__31041\,
            I => \N__31031\
        );

    \I__7008\ : LocalMux
    port map (
            O => \N__31038\,
            I => \N__31028\
        );

    \I__7007\ : InMux
    port map (
            O => \N__31037\,
            I => \N__31025\
        );

    \I__7006\ : InMux
    port map (
            O => \N__31034\,
            I => \N__31022\
        );

    \I__7005\ : LocalMux
    port map (
            O => \N__31031\,
            I => \N__31019\
        );

    \I__7004\ : Span4Mux_v
    port map (
            O => \N__31028\,
            I => \N__31014\
        );

    \I__7003\ : LocalMux
    port map (
            O => \N__31025\,
            I => \N__31014\
        );

    \I__7002\ : LocalMux
    port map (
            O => \N__31022\,
            I => \N__31011\
        );

    \I__7001\ : Span4Mux_v
    port map (
            O => \N__31019\,
            I => \N__31007\
        );

    \I__7000\ : Span4Mux_h
    port map (
            O => \N__31014\,
            I => \N__31002\
        );

    \I__6999\ : Span4Mux_v
    port map (
            O => \N__31011\,
            I => \N__31002\
        );

    \I__6998\ : InMux
    port map (
            O => \N__31010\,
            I => \N__30999\
        );

    \I__6997\ : Odrv4
    port map (
            O => \N__31007\,
            I => \b2v_inst.reg_ancho_1Z0Z_3\
        );

    \I__6996\ : Odrv4
    port map (
            O => \N__31002\,
            I => \b2v_inst.reg_ancho_1Z0Z_3\
        );

    \I__6995\ : LocalMux
    port map (
            O => \N__30999\,
            I => \b2v_inst.reg_ancho_1Z0Z_3\
        );

    \I__6994\ : CascadeMux
    port map (
            O => \N__30992\,
            I => \N__30984\
        );

    \I__6993\ : InMux
    port map (
            O => \N__30991\,
            I => \N__30972\
        );

    \I__6992\ : InMux
    port map (
            O => \N__30990\,
            I => \N__30972\
        );

    \I__6991\ : CascadeMux
    port map (
            O => \N__30989\,
            I => \N__30968\
        );

    \I__6990\ : CascadeMux
    port map (
            O => \N__30988\,
            I => \N__30965\
        );

    \I__6989\ : CascadeMux
    port map (
            O => \N__30987\,
            I => \N__30962\
        );

    \I__6988\ : InMux
    port map (
            O => \N__30984\,
            I => \N__30958\
        );

    \I__6987\ : CascadeMux
    port map (
            O => \N__30983\,
            I => \N__30953\
        );

    \I__6986\ : CascadeMux
    port map (
            O => \N__30982\,
            I => \N__30950\
        );

    \I__6985\ : CascadeMux
    port map (
            O => \N__30981\,
            I => \N__30947\
        );

    \I__6984\ : CascadeMux
    port map (
            O => \N__30980\,
            I => \N__30942\
        );

    \I__6983\ : CascadeMux
    port map (
            O => \N__30979\,
            I => \N__30938\
        );

    \I__6982\ : CascadeMux
    port map (
            O => \N__30978\,
            I => \N__30935\
        );

    \I__6981\ : InMux
    port map (
            O => \N__30977\,
            I => \N__30932\
        );

    \I__6980\ : LocalMux
    port map (
            O => \N__30972\,
            I => \N__30928\
        );

    \I__6979\ : InMux
    port map (
            O => \N__30971\,
            I => \N__30925\
        );

    \I__6978\ : InMux
    port map (
            O => \N__30968\,
            I => \N__30922\
        );

    \I__6977\ : InMux
    port map (
            O => \N__30965\,
            I => \N__30915\
        );

    \I__6976\ : InMux
    port map (
            O => \N__30962\,
            I => \N__30915\
        );

    \I__6975\ : InMux
    port map (
            O => \N__30961\,
            I => \N__30915\
        );

    \I__6974\ : LocalMux
    port map (
            O => \N__30958\,
            I => \N__30912\
        );

    \I__6973\ : InMux
    port map (
            O => \N__30957\,
            I => \N__30907\
        );

    \I__6972\ : InMux
    port map (
            O => \N__30956\,
            I => \N__30904\
        );

    \I__6971\ : InMux
    port map (
            O => \N__30953\,
            I => \N__30901\
        );

    \I__6970\ : InMux
    port map (
            O => \N__30950\,
            I => \N__30894\
        );

    \I__6969\ : InMux
    port map (
            O => \N__30947\,
            I => \N__30894\
        );

    \I__6968\ : InMux
    port map (
            O => \N__30946\,
            I => \N__30894\
        );

    \I__6967\ : InMux
    port map (
            O => \N__30945\,
            I => \N__30889\
        );

    \I__6966\ : InMux
    port map (
            O => \N__30942\,
            I => \N__30889\
        );

    \I__6965\ : InMux
    port map (
            O => \N__30941\,
            I => \N__30882\
        );

    \I__6964\ : InMux
    port map (
            O => \N__30938\,
            I => \N__30882\
        );

    \I__6963\ : InMux
    port map (
            O => \N__30935\,
            I => \N__30882\
        );

    \I__6962\ : LocalMux
    port map (
            O => \N__30932\,
            I => \N__30879\
        );

    \I__6961\ : CascadeMux
    port map (
            O => \N__30931\,
            I => \N__30876\
        );

    \I__6960\ : Span4Mux_v
    port map (
            O => \N__30928\,
            I => \N__30869\
        );

    \I__6959\ : LocalMux
    port map (
            O => \N__30925\,
            I => \N__30869\
        );

    \I__6958\ : LocalMux
    port map (
            O => \N__30922\,
            I => \N__30862\
        );

    \I__6957\ : LocalMux
    port map (
            O => \N__30915\,
            I => \N__30862\
        );

    \I__6956\ : Span4Mux_v
    port map (
            O => \N__30912\,
            I => \N__30862\
        );

    \I__6955\ : CascadeMux
    port map (
            O => \N__30911\,
            I => \N__30857\
        );

    \I__6954\ : CascadeMux
    port map (
            O => \N__30910\,
            I => \N__30854\
        );

    \I__6953\ : LocalMux
    port map (
            O => \N__30907\,
            I => \N__30849\
        );

    \I__6952\ : LocalMux
    port map (
            O => \N__30904\,
            I => \N__30849\
        );

    \I__6951\ : LocalMux
    port map (
            O => \N__30901\,
            I => \N__30846\
        );

    \I__6950\ : LocalMux
    port map (
            O => \N__30894\,
            I => \N__30843\
        );

    \I__6949\ : LocalMux
    port map (
            O => \N__30889\,
            I => \N__30840\
        );

    \I__6948\ : LocalMux
    port map (
            O => \N__30882\,
            I => \N__30837\
        );

    \I__6947\ : Span4Mux_v
    port map (
            O => \N__30879\,
            I => \N__30834\
        );

    \I__6946\ : InMux
    port map (
            O => \N__30876\,
            I => \N__30831\
        );

    \I__6945\ : InMux
    port map (
            O => \N__30875\,
            I => \N__30828\
        );

    \I__6944\ : InMux
    port map (
            O => \N__30874\,
            I => \N__30825\
        );

    \I__6943\ : Span4Mux_h
    port map (
            O => \N__30869\,
            I => \N__30820\
        );

    \I__6942\ : Span4Mux_h
    port map (
            O => \N__30862\,
            I => \N__30820\
        );

    \I__6941\ : InMux
    port map (
            O => \N__30861\,
            I => \N__30811\
        );

    \I__6940\ : InMux
    port map (
            O => \N__30860\,
            I => \N__30811\
        );

    \I__6939\ : InMux
    port map (
            O => \N__30857\,
            I => \N__30811\
        );

    \I__6938\ : InMux
    port map (
            O => \N__30854\,
            I => \N__30811\
        );

    \I__6937\ : Span4Mux_v
    port map (
            O => \N__30849\,
            I => \N__30806\
        );

    \I__6936\ : Span4Mux_v
    port map (
            O => \N__30846\,
            I => \N__30806\
        );

    \I__6935\ : Span4Mux_v
    port map (
            O => \N__30843\,
            I => \N__30799\
        );

    \I__6934\ : Span4Mux_v
    port map (
            O => \N__30840\,
            I => \N__30799\
        );

    \I__6933\ : Span4Mux_v
    port map (
            O => \N__30837\,
            I => \N__30799\
        );

    \I__6932\ : Span4Mux_h
    port map (
            O => \N__30834\,
            I => \N__30792\
        );

    \I__6931\ : LocalMux
    port map (
            O => \N__30831\,
            I => \N__30792\
        );

    \I__6930\ : LocalMux
    port map (
            O => \N__30828\,
            I => \N__30792\
        );

    \I__6929\ : LocalMux
    port map (
            O => \N__30825\,
            I => \N__30787\
        );

    \I__6928\ : Span4Mux_h
    port map (
            O => \N__30820\,
            I => \N__30787\
        );

    \I__6927\ : LocalMux
    port map (
            O => \N__30811\,
            I => \N__30780\
        );

    \I__6926\ : Sp12to4
    port map (
            O => \N__30806\,
            I => \N__30780\
        );

    \I__6925\ : Sp12to4
    port map (
            O => \N__30799\,
            I => \N__30780\
        );

    \I__6924\ : Span4Mux_h
    port map (
            O => \N__30792\,
            I => \N__30777\
        );

    \I__6923\ : Odrv4
    port map (
            O => \N__30787\,
            I => \b2v_inst.stateZ0Z_20\
        );

    \I__6922\ : Odrv12
    port map (
            O => \N__30780\,
            I => \b2v_inst.stateZ0Z_20\
        );

    \I__6921\ : Odrv4
    port map (
            O => \N__30777\,
            I => \b2v_inst.stateZ0Z_20\
        );

    \I__6920\ : InMux
    port map (
            O => \N__30770\,
            I => \N__30765\
        );

    \I__6919\ : InMux
    port map (
            O => \N__30769\,
            I => \N__30762\
        );

    \I__6918\ : InMux
    port map (
            O => \N__30768\,
            I => \N__30758\
        );

    \I__6917\ : LocalMux
    port map (
            O => \N__30765\,
            I => \N__30755\
        );

    \I__6916\ : LocalMux
    port map (
            O => \N__30762\,
            I => \N__30752\
        );

    \I__6915\ : InMux
    port map (
            O => \N__30761\,
            I => \N__30749\
        );

    \I__6914\ : LocalMux
    port map (
            O => \N__30758\,
            I => \N__30746\
        );

    \I__6913\ : Span4Mux_v
    port map (
            O => \N__30755\,
            I => \N__30743\
        );

    \I__6912\ : Span4Mux_h
    port map (
            O => \N__30752\,
            I => \N__30738\
        );

    \I__6911\ : LocalMux
    port map (
            O => \N__30749\,
            I => \N__30738\
        );

    \I__6910\ : Span4Mux_v
    port map (
            O => \N__30746\,
            I => \N__30733\
        );

    \I__6909\ : Span4Mux_h
    port map (
            O => \N__30743\,
            I => \N__30733\
        );

    \I__6908\ : Odrv4
    port map (
            O => \N__30738\,
            I => \b2v_inst.reg_anteriorZ0Z_8\
        );

    \I__6907\ : Odrv4
    port map (
            O => \N__30733\,
            I => \b2v_inst.reg_anteriorZ0Z_8\
        );

    \I__6906\ : InMux
    port map (
            O => \N__30728\,
            I => \N__30725\
        );

    \I__6905\ : LocalMux
    port map (
            O => \N__30725\,
            I => \N__30720\
        );

    \I__6904\ : InMux
    port map (
            O => \N__30724\,
            I => \N__30717\
        );

    \I__6903\ : InMux
    port map (
            O => \N__30723\,
            I => \N__30714\
        );

    \I__6902\ : Span4Mux_v
    port map (
            O => \N__30720\,
            I => \N__30709\
        );

    \I__6901\ : LocalMux
    port map (
            O => \N__30717\,
            I => \N__30709\
        );

    \I__6900\ : LocalMux
    port map (
            O => \N__30714\,
            I => \b2v_inst.reg_ancho_3Z0Z_8\
        );

    \I__6899\ : Odrv4
    port map (
            O => \N__30709\,
            I => \b2v_inst.reg_ancho_3Z0Z_8\
        );

    \I__6898\ : InMux
    port map (
            O => \N__30704\,
            I => \N__30701\
        );

    \I__6897\ : LocalMux
    port map (
            O => \N__30701\,
            I => \b2v_inst.N_544\
        );

    \I__6896\ : InMux
    port map (
            O => \N__30698\,
            I => \N__30695\
        );

    \I__6895\ : LocalMux
    port map (
            O => \N__30695\,
            I => \N__30692\
        );

    \I__6894\ : Span4Mux_v
    port map (
            O => \N__30692\,
            I => \N__30687\
        );

    \I__6893\ : InMux
    port map (
            O => \N__30691\,
            I => \N__30684\
        );

    \I__6892\ : InMux
    port map (
            O => \N__30690\,
            I => \N__30681\
        );

    \I__6891\ : Odrv4
    port map (
            O => \N__30687\,
            I => \b2v_inst.reg_ancho_3Z0Z_7\
        );

    \I__6890\ : LocalMux
    port map (
            O => \N__30684\,
            I => \b2v_inst.reg_ancho_3Z0Z_7\
        );

    \I__6889\ : LocalMux
    port map (
            O => \N__30681\,
            I => \b2v_inst.reg_ancho_3Z0Z_7\
        );

    \I__6888\ : CascadeMux
    port map (
            O => \N__30674\,
            I => \N__30671\
        );

    \I__6887\ : InMux
    port map (
            O => \N__30671\,
            I => \N__30664\
        );

    \I__6886\ : InMux
    port map (
            O => \N__30670\,
            I => \N__30664\
        );

    \I__6885\ : InMux
    port map (
            O => \N__30669\,
            I => \N__30661\
        );

    \I__6884\ : LocalMux
    port map (
            O => \N__30664\,
            I => \N__30658\
        );

    \I__6883\ : LocalMux
    port map (
            O => \N__30661\,
            I => \N__30654\
        );

    \I__6882\ : Span4Mux_h
    port map (
            O => \N__30658\,
            I => \N__30651\
        );

    \I__6881\ : InMux
    port map (
            O => \N__30657\,
            I => \N__30648\
        );

    \I__6880\ : Span4Mux_h
    port map (
            O => \N__30654\,
            I => \N__30645\
        );

    \I__6879\ : Odrv4
    port map (
            O => \N__30651\,
            I => \b2v_inst.reg_anteriorZ0Z_7\
        );

    \I__6878\ : LocalMux
    port map (
            O => \N__30648\,
            I => \b2v_inst.reg_anteriorZ0Z_7\
        );

    \I__6877\ : Odrv4
    port map (
            O => \N__30645\,
            I => \b2v_inst.reg_anteriorZ0Z_7\
        );

    \I__6876\ : InMux
    port map (
            O => \N__30638\,
            I => \N__30635\
        );

    \I__6875\ : LocalMux
    port map (
            O => \N__30635\,
            I => \b2v_inst.un1_reg_anterior_0_i_1_7\
        );

    \I__6874\ : CascadeMux
    port map (
            O => \N__30632\,
            I => \b2v_inst.data_a_escribir_RNO_0Z0Z_7_cascade_\
        );

    \I__6873\ : InMux
    port map (
            O => \N__30629\,
            I => \N__30615\
        );

    \I__6872\ : InMux
    port map (
            O => \N__30628\,
            I => \N__30615\
        );

    \I__6871\ : InMux
    port map (
            O => \N__30627\,
            I => \N__30615\
        );

    \I__6870\ : InMux
    port map (
            O => \N__30626\,
            I => \N__30601\
        );

    \I__6869\ : InMux
    port map (
            O => \N__30625\,
            I => \N__30601\
        );

    \I__6868\ : InMux
    port map (
            O => \N__30624\,
            I => \N__30594\
        );

    \I__6867\ : InMux
    port map (
            O => \N__30623\,
            I => \N__30594\
        );

    \I__6866\ : InMux
    port map (
            O => \N__30622\,
            I => \N__30594\
        );

    \I__6865\ : LocalMux
    port map (
            O => \N__30615\,
            I => \N__30591\
        );

    \I__6864\ : InMux
    port map (
            O => \N__30614\,
            I => \N__30584\
        );

    \I__6863\ : InMux
    port map (
            O => \N__30613\,
            I => \N__30584\
        );

    \I__6862\ : InMux
    port map (
            O => \N__30612\,
            I => \N__30584\
        );

    \I__6861\ : InMux
    port map (
            O => \N__30611\,
            I => \N__30577\
        );

    \I__6860\ : InMux
    port map (
            O => \N__30610\,
            I => \N__30577\
        );

    \I__6859\ : InMux
    port map (
            O => \N__30609\,
            I => \N__30577\
        );

    \I__6858\ : InMux
    port map (
            O => \N__30608\,
            I => \N__30570\
        );

    \I__6857\ : InMux
    port map (
            O => \N__30607\,
            I => \N__30570\
        );

    \I__6856\ : InMux
    port map (
            O => \N__30606\,
            I => \N__30570\
        );

    \I__6855\ : LocalMux
    port map (
            O => \N__30601\,
            I => \b2v_inst.N_711\
        );

    \I__6854\ : LocalMux
    port map (
            O => \N__30594\,
            I => \b2v_inst.N_711\
        );

    \I__6853\ : Odrv4
    port map (
            O => \N__30591\,
            I => \b2v_inst.N_711\
        );

    \I__6852\ : LocalMux
    port map (
            O => \N__30584\,
            I => \b2v_inst.N_711\
        );

    \I__6851\ : LocalMux
    port map (
            O => \N__30577\,
            I => \b2v_inst.N_711\
        );

    \I__6850\ : LocalMux
    port map (
            O => \N__30570\,
            I => \b2v_inst.N_711\
        );

    \I__6849\ : CEMux
    port map (
            O => \N__30557\,
            I => \N__30549\
        );

    \I__6848\ : CEMux
    port map (
            O => \N__30556\,
            I => \N__30546\
        );

    \I__6847\ : CEMux
    port map (
            O => \N__30555\,
            I => \N__30543\
        );

    \I__6846\ : CEMux
    port map (
            O => \N__30554\,
            I => \N__30540\
        );

    \I__6845\ : CEMux
    port map (
            O => \N__30553\,
            I => \N__30537\
        );

    \I__6844\ : CEMux
    port map (
            O => \N__30552\,
            I => \N__30534\
        );

    \I__6843\ : LocalMux
    port map (
            O => \N__30549\,
            I => \N__30531\
        );

    \I__6842\ : LocalMux
    port map (
            O => \N__30546\,
            I => \N__30528\
        );

    \I__6841\ : LocalMux
    port map (
            O => \N__30543\,
            I => \N__30525\
        );

    \I__6840\ : LocalMux
    port map (
            O => \N__30540\,
            I => \N__30522\
        );

    \I__6839\ : LocalMux
    port map (
            O => \N__30537\,
            I => \N__30517\
        );

    \I__6838\ : LocalMux
    port map (
            O => \N__30534\,
            I => \N__30517\
        );

    \I__6837\ : Span4Mux_h
    port map (
            O => \N__30531\,
            I => \N__30512\
        );

    \I__6836\ : Span4Mux_h
    port map (
            O => \N__30528\,
            I => \N__30512\
        );

    \I__6835\ : Odrv4
    port map (
            O => \N__30525\,
            I => \b2v_inst.un1_reset_inv_0\
        );

    \I__6834\ : Odrv4
    port map (
            O => \N__30522\,
            I => \b2v_inst.un1_reset_inv_0\
        );

    \I__6833\ : Odrv4
    port map (
            O => \N__30517\,
            I => \b2v_inst.un1_reset_inv_0\
        );

    \I__6832\ : Odrv4
    port map (
            O => \N__30512\,
            I => \b2v_inst.un1_reset_inv_0\
        );

    \I__6831\ : InMux
    port map (
            O => \N__30503\,
            I => \N__30500\
        );

    \I__6830\ : LocalMux
    port map (
            O => \N__30500\,
            I => \b2v_inst9.un1_cycle_counter_2_cry_1_THRU_CO\
        );

    \I__6829\ : CascadeMux
    port map (
            O => \N__30497\,
            I => \N__30494\
        );

    \I__6828\ : InMux
    port map (
            O => \N__30494\,
            I => \N__30488\
        );

    \I__6827\ : InMux
    port map (
            O => \N__30493\,
            I => \N__30485\
        );

    \I__6826\ : InMux
    port map (
            O => \N__30492\,
            I => \N__30480\
        );

    \I__6825\ : InMux
    port map (
            O => \N__30491\,
            I => \N__30480\
        );

    \I__6824\ : LocalMux
    port map (
            O => \N__30488\,
            I => \b2v_inst9.cycle_counterZ0Z_2\
        );

    \I__6823\ : LocalMux
    port map (
            O => \N__30485\,
            I => \b2v_inst9.cycle_counterZ0Z_2\
        );

    \I__6822\ : LocalMux
    port map (
            O => \N__30480\,
            I => \b2v_inst9.cycle_counterZ0Z_2\
        );

    \I__6821\ : InMux
    port map (
            O => \N__30473\,
            I => \N__30468\
        );

    \I__6820\ : InMux
    port map (
            O => \N__30472\,
            I => \N__30463\
        );

    \I__6819\ : InMux
    port map (
            O => \N__30471\,
            I => \N__30460\
        );

    \I__6818\ : LocalMux
    port map (
            O => \N__30468\,
            I => \N__30457\
        );

    \I__6817\ : InMux
    port map (
            O => \N__30467\,
            I => \N__30452\
        );

    \I__6816\ : InMux
    port map (
            O => \N__30466\,
            I => \N__30452\
        );

    \I__6815\ : LocalMux
    port map (
            O => \N__30463\,
            I => \N__30449\
        );

    \I__6814\ : LocalMux
    port map (
            O => \N__30460\,
            I => \N__30446\
        );

    \I__6813\ : Span4Mux_h
    port map (
            O => \N__30457\,
            I => \N__30443\
        );

    \I__6812\ : LocalMux
    port map (
            O => \N__30452\,
            I => \b2v_inst9.cycle_counter_RNIQAGDZ0Z_3\
        );

    \I__6811\ : Odrv4
    port map (
            O => \N__30449\,
            I => \b2v_inst9.cycle_counter_RNIQAGDZ0Z_3\
        );

    \I__6810\ : Odrv4
    port map (
            O => \N__30446\,
            I => \b2v_inst9.cycle_counter_RNIQAGDZ0Z_3\
        );

    \I__6809\ : Odrv4
    port map (
            O => \N__30443\,
            I => \b2v_inst9.cycle_counter_RNIQAGDZ0Z_3\
        );

    \I__6808\ : CascadeMux
    port map (
            O => \N__30434\,
            I => \N__30430\
        );

    \I__6807\ : InMux
    port map (
            O => \N__30433\,
            I => \N__30427\
        );

    \I__6806\ : InMux
    port map (
            O => \N__30430\,
            I => \N__30423\
        );

    \I__6805\ : LocalMux
    port map (
            O => \N__30427\,
            I => \N__30413\
        );

    \I__6804\ : InMux
    port map (
            O => \N__30426\,
            I => \N__30408\
        );

    \I__6803\ : LocalMux
    port map (
            O => \N__30423\,
            I => \N__30405\
        );

    \I__6802\ : InMux
    port map (
            O => \N__30422\,
            I => \N__30402\
        );

    \I__6801\ : InMux
    port map (
            O => \N__30421\,
            I => \N__30397\
        );

    \I__6800\ : InMux
    port map (
            O => \N__30420\,
            I => \N__30397\
        );

    \I__6799\ : InMux
    port map (
            O => \N__30419\,
            I => \N__30390\
        );

    \I__6798\ : InMux
    port map (
            O => \N__30418\,
            I => \N__30390\
        );

    \I__6797\ : InMux
    port map (
            O => \N__30417\,
            I => \N__30390\
        );

    \I__6796\ : InMux
    port map (
            O => \N__30416\,
            I => \N__30387\
        );

    \I__6795\ : Span4Mux_v
    port map (
            O => \N__30413\,
            I => \N__30384\
        );

    \I__6794\ : CascadeMux
    port map (
            O => \N__30412\,
            I => \N__30380\
        );

    \I__6793\ : CascadeMux
    port map (
            O => \N__30411\,
            I => \N__30372\
        );

    \I__6792\ : LocalMux
    port map (
            O => \N__30408\,
            I => \N__30368\
        );

    \I__6791\ : Span4Mux_v
    port map (
            O => \N__30405\,
            I => \N__30361\
        );

    \I__6790\ : LocalMux
    port map (
            O => \N__30402\,
            I => \N__30361\
        );

    \I__6789\ : LocalMux
    port map (
            O => \N__30397\,
            I => \N__30361\
        );

    \I__6788\ : LocalMux
    port map (
            O => \N__30390\,
            I => \N__30358\
        );

    \I__6787\ : LocalMux
    port map (
            O => \N__30387\,
            I => \N__30355\
        );

    \I__6786\ : Span4Mux_h
    port map (
            O => \N__30384\,
            I => \N__30352\
        );

    \I__6785\ : InMux
    port map (
            O => \N__30383\,
            I => \N__30343\
        );

    \I__6784\ : InMux
    port map (
            O => \N__30380\,
            I => \N__30343\
        );

    \I__6783\ : InMux
    port map (
            O => \N__30379\,
            I => \N__30343\
        );

    \I__6782\ : InMux
    port map (
            O => \N__30378\,
            I => \N__30343\
        );

    \I__6781\ : InMux
    port map (
            O => \N__30377\,
            I => \N__30338\
        );

    \I__6780\ : InMux
    port map (
            O => \N__30376\,
            I => \N__30338\
        );

    \I__6779\ : InMux
    port map (
            O => \N__30375\,
            I => \N__30335\
        );

    \I__6778\ : InMux
    port map (
            O => \N__30372\,
            I => \N__30330\
        );

    \I__6777\ : InMux
    port map (
            O => \N__30371\,
            I => \N__30330\
        );

    \I__6776\ : Span4Mux_v
    port map (
            O => \N__30368\,
            I => \N__30321\
        );

    \I__6775\ : Span4Mux_h
    port map (
            O => \N__30361\,
            I => \N__30321\
        );

    \I__6774\ : Span4Mux_v
    port map (
            O => \N__30358\,
            I => \N__30321\
        );

    \I__6773\ : Span4Mux_v
    port map (
            O => \N__30355\,
            I => \N__30321\
        );

    \I__6772\ : Odrv4
    port map (
            O => \N__30352\,
            I => \N_478\
        );

    \I__6771\ : LocalMux
    port map (
            O => \N__30343\,
            I => \N_478\
        );

    \I__6770\ : LocalMux
    port map (
            O => \N__30338\,
            I => \N_478\
        );

    \I__6769\ : LocalMux
    port map (
            O => \N__30335\,
            I => \N_478\
        );

    \I__6768\ : LocalMux
    port map (
            O => \N__30330\,
            I => \N_478\
        );

    \I__6767\ : Odrv4
    port map (
            O => \N__30321\,
            I => \N_478\
        );

    \I__6766\ : CascadeMux
    port map (
            O => \N__30308\,
            I => \N__30305\
        );

    \I__6765\ : InMux
    port map (
            O => \N__30305\,
            I => \N__30299\
        );

    \I__6764\ : InMux
    port map (
            O => \N__30304\,
            I => \N__30294\
        );

    \I__6763\ : InMux
    port map (
            O => \N__30303\,
            I => \N__30294\
        );

    \I__6762\ : InMux
    port map (
            O => \N__30302\,
            I => \N__30291\
        );

    \I__6761\ : LocalMux
    port map (
            O => \N__30299\,
            I => \N__30286\
        );

    \I__6760\ : LocalMux
    port map (
            O => \N__30294\,
            I => \N__30286\
        );

    \I__6759\ : LocalMux
    port map (
            O => \N__30291\,
            I => \b2v_inst9.cycle_counterZ0Z_0\
        );

    \I__6758\ : Odrv4
    port map (
            O => \N__30286\,
            I => \b2v_inst9.cycle_counterZ0Z_0\
        );

    \I__6757\ : InMux
    port map (
            O => \N__30281\,
            I => \N__30278\
        );

    \I__6756\ : LocalMux
    port map (
            O => \N__30278\,
            I => \N__30274\
        );

    \I__6755\ : CascadeMux
    port map (
            O => \N__30277\,
            I => \N__30271\
        );

    \I__6754\ : Span4Mux_h
    port map (
            O => \N__30274\,
            I => \N__30268\
        );

    \I__6753\ : InMux
    port map (
            O => \N__30271\,
            I => \N__30265\
        );

    \I__6752\ : Odrv4
    port map (
            O => \N__30268\,
            I => \SYNTHESIZED_WIRE_5_3\
        );

    \I__6751\ : LocalMux
    port map (
            O => \N__30265\,
            I => \SYNTHESIZED_WIRE_5_3\
        );

    \I__6750\ : InMux
    port map (
            O => \N__30260\,
            I => \N__30257\
        );

    \I__6749\ : LocalMux
    port map (
            O => \N__30257\,
            I => \N__30254\
        );

    \I__6748\ : Span4Mux_h
    port map (
            O => \N__30254\,
            I => \N__30251\
        );

    \I__6747\ : Odrv4
    port map (
            O => \N__30251\,
            I => \b2v_inst.pix_data_regZ0Z_3\
        );

    \I__6746\ : CEMux
    port map (
            O => \N__30248\,
            I => \N__30245\
        );

    \I__6745\ : LocalMux
    port map (
            O => \N__30245\,
            I => \N__30240\
        );

    \I__6744\ : CEMux
    port map (
            O => \N__30244\,
            I => \N__30237\
        );

    \I__6743\ : CEMux
    port map (
            O => \N__30243\,
            I => \N__30234\
        );

    \I__6742\ : Sp12to4
    port map (
            O => \N__30240\,
            I => \N__30227\
        );

    \I__6741\ : LocalMux
    port map (
            O => \N__30237\,
            I => \N__30227\
        );

    \I__6740\ : LocalMux
    port map (
            O => \N__30234\,
            I => \N__30224\
        );

    \I__6739\ : InMux
    port map (
            O => \N__30233\,
            I => \N__30221\
        );

    \I__6738\ : InMux
    port map (
            O => \N__30232\,
            I => \N__30218\
        );

    \I__6737\ : Span12Mux_h
    port map (
            O => \N__30227\,
            I => \N__30214\
        );

    \I__6736\ : Span4Mux_v
    port map (
            O => \N__30224\,
            I => \N__30211\
        );

    \I__6735\ : LocalMux
    port map (
            O => \N__30221\,
            I => \N__30208\
        );

    \I__6734\ : LocalMux
    port map (
            O => \N__30218\,
            I => \N__30205\
        );

    \I__6733\ : InMux
    port map (
            O => \N__30217\,
            I => \N__30202\
        );

    \I__6732\ : Odrv12
    port map (
            O => \N__30214\,
            I => \b2v_inst.stateZ0Z_24\
        );

    \I__6731\ : Odrv4
    port map (
            O => \N__30211\,
            I => \b2v_inst.stateZ0Z_24\
        );

    \I__6730\ : Odrv4
    port map (
            O => \N__30208\,
            I => \b2v_inst.stateZ0Z_24\
        );

    \I__6729\ : Odrv4
    port map (
            O => \N__30205\,
            I => \b2v_inst.stateZ0Z_24\
        );

    \I__6728\ : LocalMux
    port map (
            O => \N__30202\,
            I => \b2v_inst.stateZ0Z_24\
        );

    \I__6727\ : CascadeMux
    port map (
            O => \N__30191\,
            I => \N__30188\
        );

    \I__6726\ : InMux
    port map (
            O => \N__30188\,
            I => \N__30185\
        );

    \I__6725\ : LocalMux
    port map (
            O => \N__30185\,
            I => \N__30182\
        );

    \I__6724\ : Span4Mux_h
    port map (
            O => \N__30182\,
            I => \N__30179\
        );

    \I__6723\ : Odrv4
    port map (
            O => \N__30179\,
            I => \SYNTHESIZED_WIRE_1_2\
        );

    \I__6722\ : InMux
    port map (
            O => \N__30176\,
            I => \N__30172\
        );

    \I__6721\ : InMux
    port map (
            O => \N__30175\,
            I => \N__30168\
        );

    \I__6720\ : LocalMux
    port map (
            O => \N__30172\,
            I => \N__30165\
        );

    \I__6719\ : InMux
    port map (
            O => \N__30171\,
            I => \N__30162\
        );

    \I__6718\ : LocalMux
    port map (
            O => \N__30168\,
            I => \N__30159\
        );

    \I__6717\ : Span4Mux_v
    port map (
            O => \N__30165\,
            I => \N__30153\
        );

    \I__6716\ : LocalMux
    port map (
            O => \N__30162\,
            I => \N__30153\
        );

    \I__6715\ : Span12Mux_v
    port map (
            O => \N__30159\,
            I => \N__30150\
        );

    \I__6714\ : InMux
    port map (
            O => \N__30158\,
            I => \N__30147\
        );

    \I__6713\ : Span4Mux_v
    port map (
            O => \N__30153\,
            I => \N__30144\
        );

    \I__6712\ : Odrv12
    port map (
            O => \N__30150\,
            I => \b2v_inst.reg_anteriorZ0Z_4\
        );

    \I__6711\ : LocalMux
    port map (
            O => \N__30147\,
            I => \b2v_inst.reg_anteriorZ0Z_4\
        );

    \I__6710\ : Odrv4
    port map (
            O => \N__30144\,
            I => \b2v_inst.reg_anteriorZ0Z_4\
        );

    \I__6709\ : InMux
    port map (
            O => \N__30137\,
            I => \N__30133\
        );

    \I__6708\ : CascadeMux
    port map (
            O => \N__30136\,
            I => \N__30129\
        );

    \I__6707\ : LocalMux
    port map (
            O => \N__30133\,
            I => \N__30126\
        );

    \I__6706\ : InMux
    port map (
            O => \N__30132\,
            I => \N__30123\
        );

    \I__6705\ : InMux
    port map (
            O => \N__30129\,
            I => \N__30120\
        );

    \I__6704\ : Span4Mux_v
    port map (
            O => \N__30126\,
            I => \N__30115\
        );

    \I__6703\ : LocalMux
    port map (
            O => \N__30123\,
            I => \N__30115\
        );

    \I__6702\ : LocalMux
    port map (
            O => \N__30120\,
            I => \b2v_inst.reg_ancho_3Z0Z_9\
        );

    \I__6701\ : Odrv4
    port map (
            O => \N__30115\,
            I => \b2v_inst.reg_ancho_3Z0Z_9\
        );

    \I__6700\ : InMux
    port map (
            O => \N__30110\,
            I => \N__30106\
        );

    \I__6699\ : InMux
    port map (
            O => \N__30109\,
            I => \N__30103\
        );

    \I__6698\ : LocalMux
    port map (
            O => \N__30106\,
            I => \N__30100\
        );

    \I__6697\ : LocalMux
    port map (
            O => \N__30103\,
            I => \b2v_inst.eventosZ0Z_9\
        );

    \I__6696\ : Odrv4
    port map (
            O => \N__30100\,
            I => \b2v_inst.eventosZ0Z_9\
        );

    \I__6695\ : InMux
    port map (
            O => \N__30095\,
            I => \N__30092\
        );

    \I__6694\ : LocalMux
    port map (
            O => \N__30092\,
            I => \b2v_inst.N_545\
        );

    \I__6693\ : CascadeMux
    port map (
            O => \N__30089\,
            I => \b2v_inst.un1_reg_anterior_iv_0_0_0_9_cascade_\
        );

    \I__6692\ : InMux
    port map (
            O => \N__30086\,
            I => \N__30083\
        );

    \I__6691\ : LocalMux
    port map (
            O => \N__30083\,
            I => \N__30080\
        );

    \I__6690\ : Odrv4
    port map (
            O => \N__30080\,
            I => \b2v_inst.N_543\
        );

    \I__6689\ : CascadeMux
    port map (
            O => \N__30077\,
            I => \b2v_inst.un1_reg_anterior_iv_0_0_1_9_cascade_\
        );

    \I__6688\ : CascadeMux
    port map (
            O => \N__30074\,
            I => \N__30071\
        );

    \I__6687\ : InMux
    port map (
            O => \N__30071\,
            I => \N__30068\
        );

    \I__6686\ : LocalMux
    port map (
            O => \N__30068\,
            I => \N__30065\
        );

    \I__6685\ : Span4Mux_v
    port map (
            O => \N__30065\,
            I => \N__30062\
        );

    \I__6684\ : Odrv4
    port map (
            O => \N__30062\,
            I => \b2v_inst.valor_max2_6\
        );

    \I__6683\ : InMux
    port map (
            O => \N__30059\,
            I => \N__30056\
        );

    \I__6682\ : LocalMux
    port map (
            O => \N__30056\,
            I => \N__30053\
        );

    \I__6681\ : Odrv4
    port map (
            O => \N__30053\,
            I => \b2v_inst.un1_reg_anterior_iv_0_1_6\
        );

    \I__6680\ : InMux
    port map (
            O => \N__30050\,
            I => \N__30047\
        );

    \I__6679\ : LocalMux
    port map (
            O => \N__30047\,
            I => \N__30044\
        );

    \I__6678\ : Span4Mux_h
    port map (
            O => \N__30044\,
            I => \N__30041\
        );

    \I__6677\ : Odrv4
    port map (
            O => \N__30041\,
            I => \b2v_inst.data_a_escribir11_10_and\
        );

    \I__6676\ : InMux
    port map (
            O => \N__30038\,
            I => \N__30035\
        );

    \I__6675\ : LocalMux
    port map (
            O => \N__30035\,
            I => \N__30031\
        );

    \I__6674\ : InMux
    port map (
            O => \N__30034\,
            I => \N__30028\
        );

    \I__6673\ : Span4Mux_h
    port map (
            O => \N__30031\,
            I => \N__30025\
        );

    \I__6672\ : LocalMux
    port map (
            O => \N__30028\,
            I => \b2v_inst.eventosZ0Z_8\
        );

    \I__6671\ : Odrv4
    port map (
            O => \N__30025\,
            I => \b2v_inst.eventosZ0Z_8\
        );

    \I__6670\ : CascadeMux
    port map (
            O => \N__30020\,
            I => \b2v_inst.un1_reg_anterior_iv_0_0_0_8_cascade_\
        );

    \I__6669\ : InMux
    port map (
            O => \N__30017\,
            I => \N__30014\
        );

    \I__6668\ : LocalMux
    port map (
            O => \N__30014\,
            I => \N__30011\
        );

    \I__6667\ : Odrv12
    port map (
            O => \N__30011\,
            I => \b2v_inst.N_542\
        );

    \I__6666\ : CascadeMux
    port map (
            O => \N__30008\,
            I => \b2v_inst.un1_reg_anterior_iv_0_0_1_8_cascade_\
        );

    \I__6665\ : InMux
    port map (
            O => \N__30005\,
            I => \N__30000\
        );

    \I__6664\ : InMux
    port map (
            O => \N__30004\,
            I => \N__29997\
        );

    \I__6663\ : InMux
    port map (
            O => \N__30003\,
            I => \N__29994\
        );

    \I__6662\ : LocalMux
    port map (
            O => \N__30000\,
            I => \N__29989\
        );

    \I__6661\ : LocalMux
    port map (
            O => \N__29997\,
            I => \N__29989\
        );

    \I__6660\ : LocalMux
    port map (
            O => \N__29994\,
            I => \N__29984\
        );

    \I__6659\ : Span4Mux_h
    port map (
            O => \N__29989\,
            I => \N__29981\
        );

    \I__6658\ : InMux
    port map (
            O => \N__29988\,
            I => \N__29978\
        );

    \I__6657\ : InMux
    port map (
            O => \N__29987\,
            I => \N__29975\
        );

    \I__6656\ : Odrv4
    port map (
            O => \N__29984\,
            I => \b2v_inst.reg_ancho_1Z0Z_9\
        );

    \I__6655\ : Odrv4
    port map (
            O => \N__29981\,
            I => \b2v_inst.reg_ancho_1Z0Z_9\
        );

    \I__6654\ : LocalMux
    port map (
            O => \N__29978\,
            I => \b2v_inst.reg_ancho_1Z0Z_9\
        );

    \I__6653\ : LocalMux
    port map (
            O => \N__29975\,
            I => \b2v_inst.reg_ancho_1Z0Z_9\
        );

    \I__6652\ : InMux
    port map (
            O => \N__29966\,
            I => \N__29961\
        );

    \I__6651\ : InMux
    port map (
            O => \N__29965\,
            I => \N__29956\
        );

    \I__6650\ : InMux
    port map (
            O => \N__29964\,
            I => \N__29956\
        );

    \I__6649\ : LocalMux
    port map (
            O => \N__29961\,
            I => \N__29953\
        );

    \I__6648\ : LocalMux
    port map (
            O => \N__29956\,
            I => \N__29950\
        );

    \I__6647\ : Span4Mux_v
    port map (
            O => \N__29953\,
            I => \N__29945\
        );

    \I__6646\ : Span4Mux_h
    port map (
            O => \N__29950\,
            I => \N__29942\
        );

    \I__6645\ : InMux
    port map (
            O => \N__29949\,
            I => \N__29939\
        );

    \I__6644\ : InMux
    port map (
            O => \N__29948\,
            I => \N__29936\
        );

    \I__6643\ : Odrv4
    port map (
            O => \N__29945\,
            I => \b2v_inst.reg_ancho_1Z0Z_8\
        );

    \I__6642\ : Odrv4
    port map (
            O => \N__29942\,
            I => \b2v_inst.reg_ancho_1Z0Z_8\
        );

    \I__6641\ : LocalMux
    port map (
            O => \N__29939\,
            I => \b2v_inst.reg_ancho_1Z0Z_8\
        );

    \I__6640\ : LocalMux
    port map (
            O => \N__29936\,
            I => \b2v_inst.reg_ancho_1Z0Z_8\
        );

    \I__6639\ : InMux
    port map (
            O => \N__29927\,
            I => \N__29922\
        );

    \I__6638\ : CascadeMux
    port map (
            O => \N__29926\,
            I => \N__29919\
        );

    \I__6637\ : InMux
    port map (
            O => \N__29925\,
            I => \N__29916\
        );

    \I__6636\ : LocalMux
    port map (
            O => \N__29922\,
            I => \N__29913\
        );

    \I__6635\ : InMux
    port map (
            O => \N__29919\,
            I => \N__29910\
        );

    \I__6634\ : LocalMux
    port map (
            O => \N__29916\,
            I => \N__29906\
        );

    \I__6633\ : Span4Mux_v
    port map (
            O => \N__29913\,
            I => \N__29903\
        );

    \I__6632\ : LocalMux
    port map (
            O => \N__29910\,
            I => \N__29900\
        );

    \I__6631\ : CascadeMux
    port map (
            O => \N__29909\,
            I => \N__29896\
        );

    \I__6630\ : Span4Mux_v
    port map (
            O => \N__29906\,
            I => \N__29891\
        );

    \I__6629\ : Span4Mux_h
    port map (
            O => \N__29903\,
            I => \N__29891\
        );

    \I__6628\ : Span4Mux_h
    port map (
            O => \N__29900\,
            I => \N__29888\
        );

    \I__6627\ : InMux
    port map (
            O => \N__29899\,
            I => \N__29885\
        );

    \I__6626\ : InMux
    port map (
            O => \N__29896\,
            I => \N__29882\
        );

    \I__6625\ : Odrv4
    port map (
            O => \N__29891\,
            I => \b2v_inst.reg_ancho_2Z0Z_8\
        );

    \I__6624\ : Odrv4
    port map (
            O => \N__29888\,
            I => \b2v_inst.reg_ancho_2Z0Z_8\
        );

    \I__6623\ : LocalMux
    port map (
            O => \N__29885\,
            I => \b2v_inst.reg_ancho_2Z0Z_8\
        );

    \I__6622\ : LocalMux
    port map (
            O => \N__29882\,
            I => \b2v_inst.reg_ancho_2Z0Z_8\
        );

    \I__6621\ : CascadeMux
    port map (
            O => \N__29873\,
            I => \N__29870\
        );

    \I__6620\ : InMux
    port map (
            O => \N__29870\,
            I => \N__29867\
        );

    \I__6619\ : LocalMux
    port map (
            O => \N__29867\,
            I => \N__29864\
        );

    \I__6618\ : Span4Mux_h
    port map (
            O => \N__29864\,
            I => \N__29860\
        );

    \I__6617\ : InMux
    port map (
            O => \N__29863\,
            I => \N__29857\
        );

    \I__6616\ : Odrv4
    port map (
            O => \N__29860\,
            I => \b2v_inst.eventosZ0Z_3\
        );

    \I__6615\ : LocalMux
    port map (
            O => \N__29857\,
            I => \b2v_inst.eventosZ0Z_3\
        );

    \I__6614\ : InMux
    port map (
            O => \N__29852\,
            I => \N__29849\
        );

    \I__6613\ : LocalMux
    port map (
            O => \N__29849\,
            I => \N__29846\
        );

    \I__6612\ : Span4Mux_h
    port map (
            O => \N__29846\,
            I => \N__29843\
        );

    \I__6611\ : Odrv4
    port map (
            O => \N__29843\,
            I => \b2v_inst.un1_reg_anterior_0_i_1_3\
        );

    \I__6610\ : CascadeMux
    port map (
            O => \N__29840\,
            I => \N__29834\
        );

    \I__6609\ : InMux
    port map (
            O => \N__29839\,
            I => \N__29831\
        );

    \I__6608\ : InMux
    port map (
            O => \N__29838\,
            I => \N__29828\
        );

    \I__6607\ : InMux
    port map (
            O => \N__29837\,
            I => \N__29825\
        );

    \I__6606\ : InMux
    port map (
            O => \N__29834\,
            I => \N__29822\
        );

    \I__6605\ : LocalMux
    port map (
            O => \N__29831\,
            I => \N__29819\
        );

    \I__6604\ : LocalMux
    port map (
            O => \N__29828\,
            I => \N__29814\
        );

    \I__6603\ : LocalMux
    port map (
            O => \N__29825\,
            I => \N__29814\
        );

    \I__6602\ : LocalMux
    port map (
            O => \N__29822\,
            I => \N__29811\
        );

    \I__6601\ : Span4Mux_h
    port map (
            O => \N__29819\,
            I => \N__29806\
        );

    \I__6600\ : Span4Mux_v
    port map (
            O => \N__29814\,
            I => \N__29806\
        );

    \I__6599\ : Odrv4
    port map (
            O => \N__29811\,
            I => \b2v_inst.reg_anteriorZ0Z_2\
        );

    \I__6598\ : Odrv4
    port map (
            O => \N__29806\,
            I => \b2v_inst.reg_anteriorZ0Z_2\
        );

    \I__6597\ : InMux
    port map (
            O => \N__29801\,
            I => \N__29798\
        );

    \I__6596\ : LocalMux
    port map (
            O => \N__29798\,
            I => \N__29795\
        );

    \I__6595\ : Span4Mux_h
    port map (
            O => \N__29795\,
            I => \N__29792\
        );

    \I__6594\ : Odrv4
    port map (
            O => \N__29792\,
            I => \b2v_inst.data_a_escribir11_6_and\
        );

    \I__6593\ : InMux
    port map (
            O => \N__29789\,
            I => \N__29786\
        );

    \I__6592\ : LocalMux
    port map (
            O => \N__29786\,
            I => \N__29783\
        );

    \I__6591\ : Span4Mux_v
    port map (
            O => \N__29783\,
            I => \N__29780\
        );

    \I__6590\ : Sp12to4
    port map (
            O => \N__29780\,
            I => \N__29777\
        );

    \I__6589\ : Odrv12
    port map (
            O => \N__29777\,
            I => \b2v_inst.N_273\
        );

    \I__6588\ : CascadeMux
    port map (
            O => \N__29774\,
            I => \N__29771\
        );

    \I__6587\ : InMux
    port map (
            O => \N__29771\,
            I => \N__29768\
        );

    \I__6586\ : LocalMux
    port map (
            O => \N__29768\,
            I => \b2v_inst.un1_reg_anterior_iv_0_0_5\
        );

    \I__6585\ : InMux
    port map (
            O => \N__29765\,
            I => \N__29762\
        );

    \I__6584\ : LocalMux
    port map (
            O => \N__29762\,
            I => \N__29759\
        );

    \I__6583\ : Span4Mux_v
    port map (
            O => \N__29759\,
            I => \N__29756\
        );

    \I__6582\ : Odrv4
    port map (
            O => \N__29756\,
            I => \b2v_inst.N_267\
        );

    \I__6581\ : CascadeMux
    port map (
            O => \N__29753\,
            I => \b2v_inst.un1_reg_anterior_iv_0_1_5_cascade_\
        );

    \I__6580\ : CascadeMux
    port map (
            O => \N__29750\,
            I => \N__29747\
        );

    \I__6579\ : InMux
    port map (
            O => \N__29747\,
            I => \N__29744\
        );

    \I__6578\ : LocalMux
    port map (
            O => \N__29744\,
            I => \b2v_inst.data_a_escribir_RNO_0Z0Z_2\
        );

    \I__6577\ : CascadeMux
    port map (
            O => \N__29741\,
            I => \N__29738\
        );

    \I__6576\ : InMux
    port map (
            O => \N__29738\,
            I => \N__29733\
        );

    \I__6575\ : InMux
    port map (
            O => \N__29737\,
            I => \N__29730\
        );

    \I__6574\ : InMux
    port map (
            O => \N__29736\,
            I => \N__29727\
        );

    \I__6573\ : LocalMux
    port map (
            O => \N__29733\,
            I => \N__29718\
        );

    \I__6572\ : LocalMux
    port map (
            O => \N__29730\,
            I => \N__29718\
        );

    \I__6571\ : LocalMux
    port map (
            O => \N__29727\,
            I => \N__29718\
        );

    \I__6570\ : InMux
    port map (
            O => \N__29726\,
            I => \N__29715\
        );

    \I__6569\ : InMux
    port map (
            O => \N__29725\,
            I => \N__29712\
        );

    \I__6568\ : Span4Mux_v
    port map (
            O => \N__29718\,
            I => \N__29709\
        );

    \I__6567\ : LocalMux
    port map (
            O => \N__29715\,
            I => \b2v_inst.reg_ancho_2Z0Z_9\
        );

    \I__6566\ : LocalMux
    port map (
            O => \N__29712\,
            I => \b2v_inst.reg_ancho_2Z0Z_9\
        );

    \I__6565\ : Odrv4
    port map (
            O => \N__29709\,
            I => \b2v_inst.reg_ancho_2Z0Z_9\
        );

    \I__6564\ : InMux
    port map (
            O => \N__29702\,
            I => \N__29698\
        );

    \I__6563\ : InMux
    port map (
            O => \N__29701\,
            I => \N__29695\
        );

    \I__6562\ : LocalMux
    port map (
            O => \N__29698\,
            I => \N__29692\
        );

    \I__6561\ : LocalMux
    port map (
            O => \N__29695\,
            I => \N__29688\
        );

    \I__6560\ : Span4Mux_v
    port map (
            O => \N__29692\,
            I => \N__29685\
        );

    \I__6559\ : InMux
    port map (
            O => \N__29691\,
            I => \N__29682\
        );

    \I__6558\ : Odrv4
    port map (
            O => \N__29688\,
            I => \b2v_inst.reg_ancho_3Z0Z_1\
        );

    \I__6557\ : Odrv4
    port map (
            O => \N__29685\,
            I => \b2v_inst.reg_ancho_3Z0Z_1\
        );

    \I__6556\ : LocalMux
    port map (
            O => \N__29682\,
            I => \b2v_inst.reg_ancho_3Z0Z_1\
        );

    \I__6555\ : InMux
    port map (
            O => \N__29675\,
            I => \N__29671\
        );

    \I__6554\ : InMux
    port map (
            O => \N__29674\,
            I => \N__29668\
        );

    \I__6553\ : LocalMux
    port map (
            O => \N__29671\,
            I => \N__29665\
        );

    \I__6552\ : LocalMux
    port map (
            O => \N__29668\,
            I => \N__29661\
        );

    \I__6551\ : Span4Mux_v
    port map (
            O => \N__29665\,
            I => \N__29658\
        );

    \I__6550\ : InMux
    port map (
            O => \N__29664\,
            I => \N__29655\
        );

    \I__6549\ : Odrv4
    port map (
            O => \N__29661\,
            I => \b2v_inst.reg_ancho_3Z0Z_0\
        );

    \I__6548\ : Odrv4
    port map (
            O => \N__29658\,
            I => \b2v_inst.reg_ancho_3Z0Z_0\
        );

    \I__6547\ : LocalMux
    port map (
            O => \N__29655\,
            I => \b2v_inst.reg_ancho_3Z0Z_0\
        );

    \I__6546\ : InMux
    port map (
            O => \N__29648\,
            I => \N__29645\
        );

    \I__6545\ : LocalMux
    port map (
            O => \N__29645\,
            I => \N__29642\
        );

    \I__6544\ : Span4Mux_h
    port map (
            O => \N__29642\,
            I => \N__29639\
        );

    \I__6543\ : Odrv4
    port map (
            O => \N__29639\,
            I => \b2v_inst.data_a_escribir11_5_and\
        );

    \I__6542\ : InMux
    port map (
            O => \N__29636\,
            I => \N__29630\
        );

    \I__6541\ : InMux
    port map (
            O => \N__29635\,
            I => \N__29627\
        );

    \I__6540\ : InMux
    port map (
            O => \N__29634\,
            I => \N__29622\
        );

    \I__6539\ : InMux
    port map (
            O => \N__29633\,
            I => \N__29622\
        );

    \I__6538\ : LocalMux
    port map (
            O => \N__29630\,
            I => \N__29619\
        );

    \I__6537\ : LocalMux
    port map (
            O => \N__29627\,
            I => \N__29616\
        );

    \I__6536\ : LocalMux
    port map (
            O => \N__29622\,
            I => \N__29612\
        );

    \I__6535\ : Span4Mux_v
    port map (
            O => \N__29619\,
            I => \N__29609\
        );

    \I__6534\ : Span4Mux_v
    port map (
            O => \N__29616\,
            I => \N__29606\
        );

    \I__6533\ : InMux
    port map (
            O => \N__29615\,
            I => \N__29603\
        );

    \I__6532\ : Span4Mux_v
    port map (
            O => \N__29612\,
            I => \N__29600\
        );

    \I__6531\ : Odrv4
    port map (
            O => \N__29609\,
            I => \b2v_inst.reg_ancho_1Z0Z_4\
        );

    \I__6530\ : Odrv4
    port map (
            O => \N__29606\,
            I => \b2v_inst.reg_ancho_1Z0Z_4\
        );

    \I__6529\ : LocalMux
    port map (
            O => \N__29603\,
            I => \b2v_inst.reg_ancho_1Z0Z_4\
        );

    \I__6528\ : Odrv4
    port map (
            O => \N__29600\,
            I => \b2v_inst.reg_ancho_1Z0Z_4\
        );

    \I__6527\ : CascadeMux
    port map (
            O => \N__29591\,
            I => \N__29586\
        );

    \I__6526\ : CascadeMux
    port map (
            O => \N__29590\,
            I => \N__29583\
        );

    \I__6525\ : CascadeMux
    port map (
            O => \N__29589\,
            I => \N__29580\
        );

    \I__6524\ : InMux
    port map (
            O => \N__29586\,
            I => \N__29577\
        );

    \I__6523\ : InMux
    port map (
            O => \N__29583\,
            I => \N__29574\
        );

    \I__6522\ : InMux
    port map (
            O => \N__29580\,
            I => \N__29571\
        );

    \I__6521\ : LocalMux
    port map (
            O => \N__29577\,
            I => \N__29566\
        );

    \I__6520\ : LocalMux
    port map (
            O => \N__29574\,
            I => \N__29566\
        );

    \I__6519\ : LocalMux
    port map (
            O => \N__29571\,
            I => \b2v_inst.reg_ancho_3_i_4\
        );

    \I__6518\ : Odrv4
    port map (
            O => \N__29566\,
            I => \b2v_inst.reg_ancho_3_i_4\
        );

    \I__6517\ : CascadeMux
    port map (
            O => \N__29561\,
            I => \N__29556\
        );

    \I__6516\ : InMux
    port map (
            O => \N__29560\,
            I => \N__29553\
        );

    \I__6515\ : InMux
    port map (
            O => \N__29559\,
            I => \N__29548\
        );

    \I__6514\ : InMux
    port map (
            O => \N__29556\,
            I => \N__29545\
        );

    \I__6513\ : LocalMux
    port map (
            O => \N__29553\,
            I => \N__29542\
        );

    \I__6512\ : InMux
    port map (
            O => \N__29552\,
            I => \N__29539\
        );

    \I__6511\ : InMux
    port map (
            O => \N__29551\,
            I => \N__29536\
        );

    \I__6510\ : LocalMux
    port map (
            O => \N__29548\,
            I => \N__29533\
        );

    \I__6509\ : LocalMux
    port map (
            O => \N__29545\,
            I => \N__29530\
        );

    \I__6508\ : Span12Mux_h
    port map (
            O => \N__29542\,
            I => \N__29525\
        );

    \I__6507\ : LocalMux
    port map (
            O => \N__29539\,
            I => \N__29525\
        );

    \I__6506\ : LocalMux
    port map (
            O => \N__29536\,
            I => \N__29522\
        );

    \I__6505\ : Odrv4
    port map (
            O => \N__29533\,
            I => \b2v_inst.reg_ancho_1Z0Z_5\
        );

    \I__6504\ : Odrv4
    port map (
            O => \N__29530\,
            I => \b2v_inst.reg_ancho_1Z0Z_5\
        );

    \I__6503\ : Odrv12
    port map (
            O => \N__29525\,
            I => \b2v_inst.reg_ancho_1Z0Z_5\
        );

    \I__6502\ : Odrv4
    port map (
            O => \N__29522\,
            I => \b2v_inst.reg_ancho_1Z0Z_5\
        );

    \I__6501\ : CascadeMux
    port map (
            O => \N__29513\,
            I => \N__29509\
        );

    \I__6500\ : InMux
    port map (
            O => \N__29512\,
            I => \N__29506\
        );

    \I__6499\ : InMux
    port map (
            O => \N__29509\,
            I => \N__29502\
        );

    \I__6498\ : LocalMux
    port map (
            O => \N__29506\,
            I => \N__29499\
        );

    \I__6497\ : InMux
    port map (
            O => \N__29505\,
            I => \N__29496\
        );

    \I__6496\ : LocalMux
    port map (
            O => \N__29502\,
            I => \N__29493\
        );

    \I__6495\ : Odrv4
    port map (
            O => \N__29499\,
            I => \b2v_inst.reg_ancho_3_i_5\
        );

    \I__6494\ : LocalMux
    port map (
            O => \N__29496\,
            I => \b2v_inst.reg_ancho_3_i_5\
        );

    \I__6493\ : Odrv4
    port map (
            O => \N__29493\,
            I => \b2v_inst.reg_ancho_3_i_5\
        );

    \I__6492\ : InMux
    port map (
            O => \N__29486\,
            I => \N__29481\
        );

    \I__6491\ : InMux
    port map (
            O => \N__29485\,
            I => \N__29478\
        );

    \I__6490\ : InMux
    port map (
            O => \N__29484\,
            I => \N__29475\
        );

    \I__6489\ : LocalMux
    port map (
            O => \N__29481\,
            I => \N__29469\
        );

    \I__6488\ : LocalMux
    port map (
            O => \N__29478\,
            I => \N__29469\
        );

    \I__6487\ : LocalMux
    port map (
            O => \N__29475\,
            I => \N__29466\
        );

    \I__6486\ : InMux
    port map (
            O => \N__29474\,
            I => \N__29462\
        );

    \I__6485\ : Span4Mux_v
    port map (
            O => \N__29469\,
            I => \N__29457\
        );

    \I__6484\ : Span4Mux_h
    port map (
            O => \N__29466\,
            I => \N__29457\
        );

    \I__6483\ : InMux
    port map (
            O => \N__29465\,
            I => \N__29454\
        );

    \I__6482\ : LocalMux
    port map (
            O => \N__29462\,
            I => \N__29451\
        );

    \I__6481\ : Odrv4
    port map (
            O => \N__29457\,
            I => \b2v_inst.reg_ancho_1Z0Z_6\
        );

    \I__6480\ : LocalMux
    port map (
            O => \N__29454\,
            I => \b2v_inst.reg_ancho_1Z0Z_6\
        );

    \I__6479\ : Odrv12
    port map (
            O => \N__29451\,
            I => \b2v_inst.reg_ancho_1Z0Z_6\
        );

    \I__6478\ : InMux
    port map (
            O => \N__29444\,
            I => \N__29439\
        );

    \I__6477\ : InMux
    port map (
            O => \N__29443\,
            I => \N__29436\
        );

    \I__6476\ : InMux
    port map (
            O => \N__29442\,
            I => \N__29433\
        );

    \I__6475\ : LocalMux
    port map (
            O => \N__29439\,
            I => \b2v_inst.reg_ancho_3Z0Z_6\
        );

    \I__6474\ : LocalMux
    port map (
            O => \N__29436\,
            I => \b2v_inst.reg_ancho_3Z0Z_6\
        );

    \I__6473\ : LocalMux
    port map (
            O => \N__29433\,
            I => \b2v_inst.reg_ancho_3Z0Z_6\
        );

    \I__6472\ : InMux
    port map (
            O => \N__29426\,
            I => \N__29421\
        );

    \I__6471\ : CascadeMux
    port map (
            O => \N__29425\,
            I => \N__29418\
        );

    \I__6470\ : CascadeMux
    port map (
            O => \N__29424\,
            I => \N__29415\
        );

    \I__6469\ : LocalMux
    port map (
            O => \N__29421\,
            I => \N__29412\
        );

    \I__6468\ : InMux
    port map (
            O => \N__29418\,
            I => \N__29409\
        );

    \I__6467\ : InMux
    port map (
            O => \N__29415\,
            I => \N__29406\
        );

    \I__6466\ : Span4Mux_h
    port map (
            O => \N__29412\,
            I => \N__29401\
        );

    \I__6465\ : LocalMux
    port map (
            O => \N__29409\,
            I => \N__29401\
        );

    \I__6464\ : LocalMux
    port map (
            O => \N__29406\,
            I => \b2v_inst.reg_ancho_3_i_6\
        );

    \I__6463\ : Odrv4
    port map (
            O => \N__29401\,
            I => \b2v_inst.reg_ancho_3_i_6\
        );

    \I__6462\ : InMux
    port map (
            O => \N__29396\,
            I => \N__29392\
        );

    \I__6461\ : CascadeMux
    port map (
            O => \N__29395\,
            I => \N__29387\
        );

    \I__6460\ : LocalMux
    port map (
            O => \N__29392\,
            I => \N__29383\
        );

    \I__6459\ : InMux
    port map (
            O => \N__29391\,
            I => \N__29380\
        );

    \I__6458\ : InMux
    port map (
            O => \N__29390\,
            I => \N__29375\
        );

    \I__6457\ : InMux
    port map (
            O => \N__29387\,
            I => \N__29375\
        );

    \I__6456\ : InMux
    port map (
            O => \N__29386\,
            I => \N__29372\
        );

    \I__6455\ : Span4Mux_h
    port map (
            O => \N__29383\,
            I => \N__29369\
        );

    \I__6454\ : LocalMux
    port map (
            O => \N__29380\,
            I => \N__29366\
        );

    \I__6453\ : LocalMux
    port map (
            O => \N__29375\,
            I => \N__29363\
        );

    \I__6452\ : LocalMux
    port map (
            O => \N__29372\,
            I => \N__29360\
        );

    \I__6451\ : Odrv4
    port map (
            O => \N__29369\,
            I => \b2v_inst.reg_ancho_1Z0Z_7\
        );

    \I__6450\ : Odrv4
    port map (
            O => \N__29366\,
            I => \b2v_inst.reg_ancho_1Z0Z_7\
        );

    \I__6449\ : Odrv12
    port map (
            O => \N__29363\,
            I => \b2v_inst.reg_ancho_1Z0Z_7\
        );

    \I__6448\ : Odrv4
    port map (
            O => \N__29360\,
            I => \b2v_inst.reg_ancho_1Z0Z_7\
        );

    \I__6447\ : InMux
    port map (
            O => \N__29351\,
            I => \N__29346\
        );

    \I__6446\ : CascadeMux
    port map (
            O => \N__29350\,
            I => \N__29343\
        );

    \I__6445\ : CascadeMux
    port map (
            O => \N__29349\,
            I => \N__29340\
        );

    \I__6444\ : LocalMux
    port map (
            O => \N__29346\,
            I => \N__29337\
        );

    \I__6443\ : InMux
    port map (
            O => \N__29343\,
            I => \N__29334\
        );

    \I__6442\ : InMux
    port map (
            O => \N__29340\,
            I => \N__29331\
        );

    \I__6441\ : Span4Mux_h
    port map (
            O => \N__29337\,
            I => \N__29326\
        );

    \I__6440\ : LocalMux
    port map (
            O => \N__29334\,
            I => \N__29326\
        );

    \I__6439\ : LocalMux
    port map (
            O => \N__29331\,
            I => \b2v_inst.reg_ancho_3_i_7\
        );

    \I__6438\ : Odrv4
    port map (
            O => \N__29326\,
            I => \b2v_inst.reg_ancho_3_i_7\
        );

    \I__6437\ : CascadeMux
    port map (
            O => \N__29321\,
            I => \N__29316\
        );

    \I__6436\ : InMux
    port map (
            O => \N__29320\,
            I => \N__29313\
        );

    \I__6435\ : CascadeMux
    port map (
            O => \N__29319\,
            I => \N__29310\
        );

    \I__6434\ : InMux
    port map (
            O => \N__29316\,
            I => \N__29307\
        );

    \I__6433\ : LocalMux
    port map (
            O => \N__29313\,
            I => \N__29304\
        );

    \I__6432\ : InMux
    port map (
            O => \N__29310\,
            I => \N__29301\
        );

    \I__6431\ : LocalMux
    port map (
            O => \N__29307\,
            I => \N__29298\
        );

    \I__6430\ : Odrv4
    port map (
            O => \N__29304\,
            I => \b2v_inst.reg_ancho_3_i_8\
        );

    \I__6429\ : LocalMux
    port map (
            O => \N__29301\,
            I => \b2v_inst.reg_ancho_3_i_8\
        );

    \I__6428\ : Odrv4
    port map (
            O => \N__29298\,
            I => \b2v_inst.reg_ancho_3_i_8\
        );

    \I__6427\ : CascadeMux
    port map (
            O => \N__29291\,
            I => \N__29287\
        );

    \I__6426\ : CascadeMux
    port map (
            O => \N__29290\,
            I => \N__29283\
        );

    \I__6425\ : InMux
    port map (
            O => \N__29287\,
            I => \N__29280\
        );

    \I__6424\ : CascadeMux
    port map (
            O => \N__29286\,
            I => \N__29277\
        );

    \I__6423\ : InMux
    port map (
            O => \N__29283\,
            I => \N__29274\
        );

    \I__6422\ : LocalMux
    port map (
            O => \N__29280\,
            I => \N__29271\
        );

    \I__6421\ : InMux
    port map (
            O => \N__29277\,
            I => \N__29268\
        );

    \I__6420\ : LocalMux
    port map (
            O => \N__29274\,
            I => \N__29265\
        );

    \I__6419\ : Odrv4
    port map (
            O => \N__29271\,
            I => \b2v_inst.reg_ancho_3_i_9\
        );

    \I__6418\ : LocalMux
    port map (
            O => \N__29268\,
            I => \b2v_inst.reg_ancho_3_i_9\
        );

    \I__6417\ : Odrv4
    port map (
            O => \N__29265\,
            I => \b2v_inst.reg_ancho_3_i_9\
        );

    \I__6416\ : InMux
    port map (
            O => \N__29258\,
            I => \N__29253\
        );

    \I__6415\ : InMux
    port map (
            O => \N__29257\,
            I => \N__29250\
        );

    \I__6414\ : InMux
    port map (
            O => \N__29256\,
            I => \N__29247\
        );

    \I__6413\ : LocalMux
    port map (
            O => \N__29253\,
            I => \N__29240\
        );

    \I__6412\ : LocalMux
    port map (
            O => \N__29250\,
            I => \N__29240\
        );

    \I__6411\ : LocalMux
    port map (
            O => \N__29247\,
            I => \N__29237\
        );

    \I__6410\ : InMux
    port map (
            O => \N__29246\,
            I => \N__29234\
        );

    \I__6409\ : InMux
    port map (
            O => \N__29245\,
            I => \N__29231\
        );

    \I__6408\ : Span4Mux_v
    port map (
            O => \N__29240\,
            I => \N__29228\
        );

    \I__6407\ : Span4Mux_v
    port map (
            O => \N__29237\,
            I => \N__29225\
        );

    \I__6406\ : LocalMux
    port map (
            O => \N__29234\,
            I => \N__29220\
        );

    \I__6405\ : LocalMux
    port map (
            O => \N__29231\,
            I => \N__29220\
        );

    \I__6404\ : Odrv4
    port map (
            O => \N__29228\,
            I => \b2v_inst.reg_ancho_1Z0Z_10\
        );

    \I__6403\ : Odrv4
    port map (
            O => \N__29225\,
            I => \b2v_inst.reg_ancho_1Z0Z_10\
        );

    \I__6402\ : Odrv4
    port map (
            O => \N__29220\,
            I => \b2v_inst.reg_ancho_1Z0Z_10\
        );

    \I__6401\ : CascadeMux
    port map (
            O => \N__29213\,
            I => \N__29209\
        );

    \I__6400\ : CascadeMux
    port map (
            O => \N__29212\,
            I => \N__29205\
        );

    \I__6399\ : InMux
    port map (
            O => \N__29209\,
            I => \N__29202\
        );

    \I__6398\ : CascadeMux
    port map (
            O => \N__29208\,
            I => \N__29199\
        );

    \I__6397\ : InMux
    port map (
            O => \N__29205\,
            I => \N__29196\
        );

    \I__6396\ : LocalMux
    port map (
            O => \N__29202\,
            I => \N__29193\
        );

    \I__6395\ : InMux
    port map (
            O => \N__29199\,
            I => \N__29190\
        );

    \I__6394\ : LocalMux
    port map (
            O => \N__29196\,
            I => \N__29187\
        );

    \I__6393\ : Odrv4
    port map (
            O => \N__29193\,
            I => \b2v_inst.reg_ancho_3_i_10\
        );

    \I__6392\ : LocalMux
    port map (
            O => \N__29190\,
            I => \b2v_inst.reg_ancho_3_i_10\
        );

    \I__6391\ : Odrv4
    port map (
            O => \N__29187\,
            I => \b2v_inst.reg_ancho_3_i_10\
        );

    \I__6390\ : InMux
    port map (
            O => \N__29180\,
            I => \b2v_inst.valor_max_final40\
        );

    \I__6389\ : InMux
    port map (
            O => \N__29177\,
            I => \N__29174\
        );

    \I__6388\ : LocalMux
    port map (
            O => \N__29174\,
            I => \N__29171\
        );

    \I__6387\ : Span4Mux_v
    port map (
            O => \N__29171\,
            I => \N__29168\
        );

    \I__6386\ : Odrv4
    port map (
            O => \N__29168\,
            I => \b2v_inst.valor_max_final40_THRU_CO\
        );

    \I__6385\ : InMux
    port map (
            O => \N__29165\,
            I => \b2v_inst.un2_valor_max2\
        );

    \I__6384\ : InMux
    port map (
            O => \N__29162\,
            I => \N__29159\
        );

    \I__6383\ : LocalMux
    port map (
            O => \N__29159\,
            I => \N__29154\
        );

    \I__6382\ : InMux
    port map (
            O => \N__29158\,
            I => \N__29150\
        );

    \I__6381\ : InMux
    port map (
            O => \N__29157\,
            I => \N__29147\
        );

    \I__6380\ : Span4Mux_v
    port map (
            O => \N__29154\,
            I => \N__29144\
        );

    \I__6379\ : InMux
    port map (
            O => \N__29153\,
            I => \N__29141\
        );

    \I__6378\ : LocalMux
    port map (
            O => \N__29150\,
            I => \N__29138\
        );

    \I__6377\ : LocalMux
    port map (
            O => \N__29147\,
            I => \N__29135\
        );

    \I__6376\ : Span4Mux_h
    port map (
            O => \N__29144\,
            I => \N__29130\
        );

    \I__6375\ : LocalMux
    port map (
            O => \N__29141\,
            I => \N__29130\
        );

    \I__6374\ : Span4Mux_v
    port map (
            O => \N__29138\,
            I => \N__29127\
        );

    \I__6373\ : Odrv4
    port map (
            O => \N__29135\,
            I => \b2v_inst.reg_anteriorZ0Z_3\
        );

    \I__6372\ : Odrv4
    port map (
            O => \N__29130\,
            I => \b2v_inst.reg_anteriorZ0Z_3\
        );

    \I__6371\ : Odrv4
    port map (
            O => \N__29127\,
            I => \b2v_inst.reg_anteriorZ0Z_3\
        );

    \I__6370\ : CascadeMux
    port map (
            O => \N__29120\,
            I => \N__29117\
        );

    \I__6369\ : InMux
    port map (
            O => \N__29117\,
            I => \N__29114\
        );

    \I__6368\ : LocalMux
    port map (
            O => \N__29114\,
            I => \N__29111\
        );

    \I__6367\ : Span4Mux_v
    port map (
            O => \N__29111\,
            I => \N__29108\
        );

    \I__6366\ : Odrv4
    port map (
            O => \N__29108\,
            I => \b2v_inst.data_a_escribir_RNO_0Z0Z_3\
        );

    \I__6365\ : InMux
    port map (
            O => \N__29105\,
            I => \N__29102\
        );

    \I__6364\ : LocalMux
    port map (
            O => \N__29102\,
            I => \N__29098\
        );

    \I__6363\ : InMux
    port map (
            O => \N__29101\,
            I => \N__29094\
        );

    \I__6362\ : Span4Mux_h
    port map (
            O => \N__29098\,
            I => \N__29091\
        );

    \I__6361\ : InMux
    port map (
            O => \N__29097\,
            I => \N__29087\
        );

    \I__6360\ : LocalMux
    port map (
            O => \N__29094\,
            I => \N__29084\
        );

    \I__6359\ : Span4Mux_v
    port map (
            O => \N__29091\,
            I => \N__29081\
        );

    \I__6358\ : InMux
    port map (
            O => \N__29090\,
            I => \N__29078\
        );

    \I__6357\ : LocalMux
    port map (
            O => \N__29087\,
            I => \N__29073\
        );

    \I__6356\ : Span4Mux_v
    port map (
            O => \N__29084\,
            I => \N__29073\
        );

    \I__6355\ : Odrv4
    port map (
            O => \N__29081\,
            I => \b2v_inst.reg_anteriorZ0Z_5\
        );

    \I__6354\ : LocalMux
    port map (
            O => \N__29078\,
            I => \b2v_inst.reg_anteriorZ0Z_5\
        );

    \I__6353\ : Odrv4
    port map (
            O => \N__29073\,
            I => \b2v_inst.reg_anteriorZ0Z_5\
        );

    \I__6352\ : InMux
    port map (
            O => \N__29066\,
            I => \N__29062\
        );

    \I__6351\ : InMux
    port map (
            O => \N__29065\,
            I => \N__29057\
        );

    \I__6350\ : LocalMux
    port map (
            O => \N__29062\,
            I => \N__29054\
        );

    \I__6349\ : InMux
    port map (
            O => \N__29061\,
            I => \N__29049\
        );

    \I__6348\ : InMux
    port map (
            O => \N__29060\,
            I => \N__29049\
        );

    \I__6347\ : LocalMux
    port map (
            O => \N__29057\,
            I => \N__29046\
        );

    \I__6346\ : Span4Mux_v
    port map (
            O => \N__29054\,
            I => \N__29042\
        );

    \I__6345\ : LocalMux
    port map (
            O => \N__29049\,
            I => \N__29039\
        );

    \I__6344\ : Span4Mux_v
    port map (
            O => \N__29046\,
            I => \N__29036\
        );

    \I__6343\ : InMux
    port map (
            O => \N__29045\,
            I => \N__29033\
        );

    \I__6342\ : Odrv4
    port map (
            O => \N__29042\,
            I => \b2v_inst.reg_ancho_1Z0Z_0\
        );

    \I__6341\ : Odrv12
    port map (
            O => \N__29039\,
            I => \b2v_inst.reg_ancho_1Z0Z_0\
        );

    \I__6340\ : Odrv4
    port map (
            O => \N__29036\,
            I => \b2v_inst.reg_ancho_1Z0Z_0\
        );

    \I__6339\ : LocalMux
    port map (
            O => \N__29033\,
            I => \b2v_inst.reg_ancho_1Z0Z_0\
        );

    \I__6338\ : CascadeMux
    port map (
            O => \N__29024\,
            I => \N__29019\
        );

    \I__6337\ : InMux
    port map (
            O => \N__29023\,
            I => \N__29016\
        );

    \I__6336\ : CascadeMux
    port map (
            O => \N__29022\,
            I => \N__29013\
        );

    \I__6335\ : InMux
    port map (
            O => \N__29019\,
            I => \N__29010\
        );

    \I__6334\ : LocalMux
    port map (
            O => \N__29016\,
            I => \N__29007\
        );

    \I__6333\ : InMux
    port map (
            O => \N__29013\,
            I => \N__29004\
        );

    \I__6332\ : LocalMux
    port map (
            O => \N__29010\,
            I => \N__29001\
        );

    \I__6331\ : Odrv4
    port map (
            O => \N__29007\,
            I => \b2v_inst.reg_ancho_3_i_0\
        );

    \I__6330\ : LocalMux
    port map (
            O => \N__29004\,
            I => \b2v_inst.reg_ancho_3_i_0\
        );

    \I__6329\ : Odrv4
    port map (
            O => \N__29001\,
            I => \b2v_inst.reg_ancho_3_i_0\
        );

    \I__6328\ : InMux
    port map (
            O => \N__28994\,
            I => \N__28991\
        );

    \I__6327\ : LocalMux
    port map (
            O => \N__28991\,
            I => \N__28987\
        );

    \I__6326\ : InMux
    port map (
            O => \N__28990\,
            I => \N__28984\
        );

    \I__6325\ : Span4Mux_v
    port map (
            O => \N__28987\,
            I => \N__28977\
        );

    \I__6324\ : LocalMux
    port map (
            O => \N__28984\,
            I => \N__28977\
        );

    \I__6323\ : InMux
    port map (
            O => \N__28983\,
            I => \N__28972\
        );

    \I__6322\ : InMux
    port map (
            O => \N__28982\,
            I => \N__28972\
        );

    \I__6321\ : Span4Mux_v
    port map (
            O => \N__28977\,
            I => \N__28968\
        );

    \I__6320\ : LocalMux
    port map (
            O => \N__28972\,
            I => \N__28965\
        );

    \I__6319\ : InMux
    port map (
            O => \N__28971\,
            I => \N__28962\
        );

    \I__6318\ : Span4Mux_h
    port map (
            O => \N__28968\,
            I => \N__28959\
        );

    \I__6317\ : Odrv12
    port map (
            O => \N__28965\,
            I => \b2v_inst.reg_ancho_1Z0Z_1\
        );

    \I__6316\ : LocalMux
    port map (
            O => \N__28962\,
            I => \b2v_inst.reg_ancho_1Z0Z_1\
        );

    \I__6315\ : Odrv4
    port map (
            O => \N__28959\,
            I => \b2v_inst.reg_ancho_1Z0Z_1\
        );

    \I__6314\ : CascadeMux
    port map (
            O => \N__28952\,
            I => \N__28948\
        );

    \I__6313\ : CascadeMux
    port map (
            O => \N__28951\,
            I => \N__28945\
        );

    \I__6312\ : InMux
    port map (
            O => \N__28948\,
            I => \N__28941\
        );

    \I__6311\ : InMux
    port map (
            O => \N__28945\,
            I => \N__28938\
        );

    \I__6310\ : CascadeMux
    port map (
            O => \N__28944\,
            I => \N__28935\
        );

    \I__6309\ : LocalMux
    port map (
            O => \N__28941\,
            I => \N__28932\
        );

    \I__6308\ : LocalMux
    port map (
            O => \N__28938\,
            I => \N__28929\
        );

    \I__6307\ : InMux
    port map (
            O => \N__28935\,
            I => \N__28926\
        );

    \I__6306\ : Span4Mux_h
    port map (
            O => \N__28932\,
            I => \N__28923\
        );

    \I__6305\ : Odrv4
    port map (
            O => \N__28929\,
            I => \b2v_inst.reg_ancho_3_i_1\
        );

    \I__6304\ : LocalMux
    port map (
            O => \N__28926\,
            I => \b2v_inst.reg_ancho_3_i_1\
        );

    \I__6303\ : Odrv4
    port map (
            O => \N__28923\,
            I => \b2v_inst.reg_ancho_3_i_1\
        );

    \I__6302\ : CascadeMux
    port map (
            O => \N__28916\,
            I => \N__28912\
        );

    \I__6301\ : CascadeMux
    port map (
            O => \N__28915\,
            I => \N__28908\
        );

    \I__6300\ : InMux
    port map (
            O => \N__28912\,
            I => \N__28905\
        );

    \I__6299\ : CascadeMux
    port map (
            O => \N__28911\,
            I => \N__28902\
        );

    \I__6298\ : InMux
    port map (
            O => \N__28908\,
            I => \N__28899\
        );

    \I__6297\ : LocalMux
    port map (
            O => \N__28905\,
            I => \N__28896\
        );

    \I__6296\ : InMux
    port map (
            O => \N__28902\,
            I => \N__28893\
        );

    \I__6295\ : LocalMux
    port map (
            O => \N__28899\,
            I => \N__28890\
        );

    \I__6294\ : Odrv4
    port map (
            O => \N__28896\,
            I => \b2v_inst.reg_ancho_3_i_2\
        );

    \I__6293\ : LocalMux
    port map (
            O => \N__28893\,
            I => \b2v_inst.reg_ancho_3_i_2\
        );

    \I__6292\ : Odrv4
    port map (
            O => \N__28890\,
            I => \b2v_inst.reg_ancho_3_i_2\
        );

    \I__6291\ : CascadeMux
    port map (
            O => \N__28883\,
            I => \N__28878\
        );

    \I__6290\ : InMux
    port map (
            O => \N__28882\,
            I => \N__28875\
        );

    \I__6289\ : CascadeMux
    port map (
            O => \N__28881\,
            I => \N__28872\
        );

    \I__6288\ : InMux
    port map (
            O => \N__28878\,
            I => \N__28869\
        );

    \I__6287\ : LocalMux
    port map (
            O => \N__28875\,
            I => \N__28866\
        );

    \I__6286\ : InMux
    port map (
            O => \N__28872\,
            I => \N__28863\
        );

    \I__6285\ : LocalMux
    port map (
            O => \N__28869\,
            I => \N__28860\
        );

    \I__6284\ : Odrv4
    port map (
            O => \N__28866\,
            I => \b2v_inst.reg_ancho_3_i_3\
        );

    \I__6283\ : LocalMux
    port map (
            O => \N__28863\,
            I => \b2v_inst.reg_ancho_3_i_3\
        );

    \I__6282\ : Odrv4
    port map (
            O => \N__28860\,
            I => \b2v_inst.reg_ancho_3_i_3\
        );

    \I__6281\ : InMux
    port map (
            O => \N__28853\,
            I => \N__28849\
        );

    \I__6280\ : InMux
    port map (
            O => \N__28852\,
            I => \N__28846\
        );

    \I__6279\ : LocalMux
    port map (
            O => \N__28849\,
            I => \SYNTHESIZED_WIRE_5_7\
        );

    \I__6278\ : LocalMux
    port map (
            O => \N__28846\,
            I => \SYNTHESIZED_WIRE_5_7\
        );

    \I__6277\ : InMux
    port map (
            O => \N__28841\,
            I => \N__28836\
        );

    \I__6276\ : InMux
    port map (
            O => \N__28840\,
            I => \N__28833\
        );

    \I__6275\ : InMux
    port map (
            O => \N__28839\,
            I => \N__28830\
        );

    \I__6274\ : LocalMux
    port map (
            O => \N__28836\,
            I => \SYNTHESIZED_WIRE_5_6\
        );

    \I__6273\ : LocalMux
    port map (
            O => \N__28833\,
            I => \SYNTHESIZED_WIRE_5_6\
        );

    \I__6272\ : LocalMux
    port map (
            O => \N__28830\,
            I => \SYNTHESIZED_WIRE_5_6\
        );

    \I__6271\ : InMux
    port map (
            O => \N__28823\,
            I => \N__28820\
        );

    \I__6270\ : LocalMux
    port map (
            O => \N__28820\,
            I => \b2v_inst.un12_pix_count_intlto7_N_3LZ0Z3\
        );

    \I__6269\ : InMux
    port map (
            O => \N__28817\,
            I => \N__28814\
        );

    \I__6268\ : LocalMux
    port map (
            O => \N__28814\,
            I => \N__28810\
        );

    \I__6267\ : InMux
    port map (
            O => \N__28813\,
            I => \N__28807\
        );

    \I__6266\ : Odrv12
    port map (
            O => \N__28810\,
            I => \SYNTHESIZED_WIRE_10_5\
        );

    \I__6265\ : LocalMux
    port map (
            O => \N__28807\,
            I => \SYNTHESIZED_WIRE_10_5\
        );

    \I__6264\ : InMux
    port map (
            O => \N__28802\,
            I => \N__28799\
        );

    \I__6263\ : LocalMux
    port map (
            O => \N__28799\,
            I => \N__28796\
        );

    \I__6262\ : Span4Mux_h
    port map (
            O => \N__28796\,
            I => \N__28792\
        );

    \I__6261\ : InMux
    port map (
            O => \N__28795\,
            I => \N__28789\
        );

    \I__6260\ : Odrv4
    port map (
            O => \N__28792\,
            I => \SYNTHESIZED_WIRE_5_5\
        );

    \I__6259\ : LocalMux
    port map (
            O => \N__28789\,
            I => \SYNTHESIZED_WIRE_5_5\
        );

    \I__6258\ : CEMux
    port map (
            O => \N__28784\,
            I => \N__28780\
        );

    \I__6257\ : CEMux
    port map (
            O => \N__28783\,
            I => \N__28776\
        );

    \I__6256\ : LocalMux
    port map (
            O => \N__28780\,
            I => \N__28773\
        );

    \I__6255\ : CEMux
    port map (
            O => \N__28779\,
            I => \N__28770\
        );

    \I__6254\ : LocalMux
    port map (
            O => \N__28776\,
            I => \N__28767\
        );

    \I__6253\ : Span4Mux_v
    port map (
            O => \N__28773\,
            I => \N__28764\
        );

    \I__6252\ : LocalMux
    port map (
            O => \N__28770\,
            I => \N__28761\
        );

    \I__6251\ : Sp12to4
    port map (
            O => \N__28767\,
            I => \N__28757\
        );

    \I__6250\ : Span4Mux_h
    port map (
            O => \N__28764\,
            I => \N__28752\
        );

    \I__6249\ : Span4Mux_h
    port map (
            O => \N__28761\,
            I => \N__28752\
        );

    \I__6248\ : CascadeMux
    port map (
            O => \N__28760\,
            I => \N__28748\
        );

    \I__6247\ : Span12Mux_h
    port map (
            O => \N__28757\,
            I => \N__28745\
        );

    \I__6246\ : Span4Mux_h
    port map (
            O => \N__28752\,
            I => \N__28742\
        );

    \I__6245\ : InMux
    port map (
            O => \N__28751\,
            I => \N__28739\
        );

    \I__6244\ : InMux
    port map (
            O => \N__28748\,
            I => \N__28736\
        );

    \I__6243\ : Odrv12
    port map (
            O => \N__28745\,
            I => \b2v_inst4.pix_count_int_0_sqmuxa\
        );

    \I__6242\ : Odrv4
    port map (
            O => \N__28742\,
            I => \b2v_inst4.pix_count_int_0_sqmuxa\
        );

    \I__6241\ : LocalMux
    port map (
            O => \N__28739\,
            I => \b2v_inst4.pix_count_int_0_sqmuxa\
        );

    \I__6240\ : LocalMux
    port map (
            O => \N__28736\,
            I => \b2v_inst4.pix_count_int_0_sqmuxa\
        );

    \I__6239\ : CascadeMux
    port map (
            O => \N__28727\,
            I => \N__28723\
        );

    \I__6238\ : InMux
    port map (
            O => \N__28726\,
            I => \N__28720\
        );

    \I__6237\ : InMux
    port map (
            O => \N__28723\,
            I => \N__28717\
        );

    \I__6236\ : LocalMux
    port map (
            O => \N__28720\,
            I => \N__28712\
        );

    \I__6235\ : LocalMux
    port map (
            O => \N__28717\,
            I => \N__28712\
        );

    \I__6234\ : Odrv4
    port map (
            O => \N__28712\,
            I => \b2v_inst9.N_175_i\
        );

    \I__6233\ : InMux
    port map (
            O => \N__28709\,
            I => \N__28704\
        );

    \I__6232\ : InMux
    port map (
            O => \N__28708\,
            I => \N__28699\
        );

    \I__6231\ : InMux
    port map (
            O => \N__28707\,
            I => \N__28699\
        );

    \I__6230\ : LocalMux
    port map (
            O => \N__28704\,
            I => \b2v_inst9.bit_counterZ0Z_0\
        );

    \I__6229\ : LocalMux
    port map (
            O => \N__28699\,
            I => \b2v_inst9.bit_counterZ0Z_0\
        );

    \I__6228\ : InMux
    port map (
            O => \N__28694\,
            I => \N__28689\
        );

    \I__6227\ : InMux
    port map (
            O => \N__28693\,
            I => \N__28684\
        );

    \I__6226\ : InMux
    port map (
            O => \N__28692\,
            I => \N__28684\
        );

    \I__6225\ : LocalMux
    port map (
            O => \N__28689\,
            I => \b2v_inst9.bit_counterZ1Z_1\
        );

    \I__6224\ : LocalMux
    port map (
            O => \N__28684\,
            I => \b2v_inst9.bit_counterZ1Z_1\
        );

    \I__6223\ : InMux
    port map (
            O => \N__28679\,
            I => \b2v_inst9.un1_bit_counter_3_cry_0\
        );

    \I__6222\ : CascadeMux
    port map (
            O => \N__28676\,
            I => \N__28672\
        );

    \I__6221\ : InMux
    port map (
            O => \N__28675\,
            I => \N__28668\
        );

    \I__6220\ : InMux
    port map (
            O => \N__28672\,
            I => \N__28663\
        );

    \I__6219\ : InMux
    port map (
            O => \N__28671\,
            I => \N__28663\
        );

    \I__6218\ : LocalMux
    port map (
            O => \N__28668\,
            I => \b2v_inst9.bit_counterZ0Z_2\
        );

    \I__6217\ : LocalMux
    port map (
            O => \N__28663\,
            I => \b2v_inst9.bit_counterZ0Z_2\
        );

    \I__6216\ : InMux
    port map (
            O => \N__28658\,
            I => \b2v_inst9.un1_bit_counter_3_cry_1\
        );

    \I__6215\ : InMux
    port map (
            O => \N__28655\,
            I => \N__28647\
        );

    \I__6214\ : InMux
    port map (
            O => \N__28654\,
            I => \N__28647\
        );

    \I__6213\ : InMux
    port map (
            O => \N__28653\,
            I => \N__28642\
        );

    \I__6212\ : InMux
    port map (
            O => \N__28652\,
            I => \N__28642\
        );

    \I__6211\ : LocalMux
    port map (
            O => \N__28647\,
            I => \b2v_inst9.fsm_state_RNIND1P1Z0Z_0\
        );

    \I__6210\ : LocalMux
    port map (
            O => \N__28642\,
            I => \b2v_inst9.fsm_state_RNIND1P1Z0Z_0\
        );

    \I__6209\ : InMux
    port map (
            O => \N__28637\,
            I => \b2v_inst9.un1_bit_counter_3_cry_2\
        );

    \I__6208\ : InMux
    port map (
            O => \N__28634\,
            I => \N__28629\
        );

    \I__6207\ : InMux
    port map (
            O => \N__28633\,
            I => \N__28624\
        );

    \I__6206\ : InMux
    port map (
            O => \N__28632\,
            I => \N__28624\
        );

    \I__6205\ : LocalMux
    port map (
            O => \N__28629\,
            I => \b2v_inst9.bit_counterZ0Z_3\
        );

    \I__6204\ : LocalMux
    port map (
            O => \N__28624\,
            I => \b2v_inst9.bit_counterZ0Z_3\
        );

    \I__6203\ : InMux
    port map (
            O => \N__28619\,
            I => \N__28616\
        );

    \I__6202\ : LocalMux
    port map (
            O => \N__28616\,
            I => \N__28611\
        );

    \I__6201\ : InMux
    port map (
            O => \N__28615\,
            I => \N__28607\
        );

    \I__6200\ : InMux
    port map (
            O => \N__28614\,
            I => \N__28604\
        );

    \I__6199\ : Span4Mux_h
    port map (
            O => \N__28611\,
            I => \N__28601\
        );

    \I__6198\ : InMux
    port map (
            O => \N__28610\,
            I => \N__28598\
        );

    \I__6197\ : LocalMux
    port map (
            O => \N__28607\,
            I => \b2v_inst.reg_anteriorZ0Z_0\
        );

    \I__6196\ : LocalMux
    port map (
            O => \N__28604\,
            I => \b2v_inst.reg_anteriorZ0Z_0\
        );

    \I__6195\ : Odrv4
    port map (
            O => \N__28601\,
            I => \b2v_inst.reg_anteriorZ0Z_0\
        );

    \I__6194\ : LocalMux
    port map (
            O => \N__28598\,
            I => \b2v_inst.reg_anteriorZ0Z_0\
        );

    \I__6193\ : InMux
    port map (
            O => \N__28589\,
            I => \N__28585\
        );

    \I__6192\ : InMux
    port map (
            O => \N__28588\,
            I => \N__28581\
        );

    \I__6191\ : LocalMux
    port map (
            O => \N__28585\,
            I => \N__28578\
        );

    \I__6190\ : InMux
    port map (
            O => \N__28584\,
            I => \N__28575\
        );

    \I__6189\ : LocalMux
    port map (
            O => \N__28581\,
            I => \N__28571\
        );

    \I__6188\ : Span4Mux_h
    port map (
            O => \N__28578\,
            I => \N__28566\
        );

    \I__6187\ : LocalMux
    port map (
            O => \N__28575\,
            I => \N__28566\
        );

    \I__6186\ : InMux
    port map (
            O => \N__28574\,
            I => \N__28563\
        );

    \I__6185\ : Span4Mux_h
    port map (
            O => \N__28571\,
            I => \N__28558\
        );

    \I__6184\ : Span4Mux_v
    port map (
            O => \N__28566\,
            I => \N__28558\
        );

    \I__6183\ : LocalMux
    port map (
            O => \N__28563\,
            I => \b2v_inst.reg_anteriorZ0Z_1\
        );

    \I__6182\ : Odrv4
    port map (
            O => \N__28558\,
            I => \b2v_inst.reg_anteriorZ0Z_1\
        );

    \I__6181\ : InMux
    port map (
            O => \N__28553\,
            I => \N__28550\
        );

    \I__6180\ : LocalMux
    port map (
            O => \N__28550\,
            I => \N__28547\
        );

    \I__6179\ : Span4Mux_v
    port map (
            O => \N__28547\,
            I => \N__28543\
        );

    \I__6178\ : InMux
    port map (
            O => \N__28546\,
            I => \N__28540\
        );

    \I__6177\ : Span4Mux_h
    port map (
            O => \N__28543\,
            I => \N__28537\
        );

    \I__6176\ : LocalMux
    port map (
            O => \N__28540\,
            I => \N__28534\
        );

    \I__6175\ : Odrv4
    port map (
            O => \N__28537\,
            I => \b2v_inst.N_654_2\
        );

    \I__6174\ : Odrv4
    port map (
            O => \N__28534\,
            I => \b2v_inst.N_654_2\
        );

    \I__6173\ : CascadeMux
    port map (
            O => \N__28529\,
            I => \b2v_inst.un1_reset_inv_0_0_tz_cascade_\
        );

    \I__6172\ : InMux
    port map (
            O => \N__28526\,
            I => \N__28522\
        );

    \I__6171\ : InMux
    port map (
            O => \N__28525\,
            I => \N__28518\
        );

    \I__6170\ : LocalMux
    port map (
            O => \N__28522\,
            I => \N__28515\
        );

    \I__6169\ : InMux
    port map (
            O => \N__28521\,
            I => \N__28511\
        );

    \I__6168\ : LocalMux
    port map (
            O => \N__28518\,
            I => \N__28508\
        );

    \I__6167\ : Span4Mux_h
    port map (
            O => \N__28515\,
            I => \N__28505\
        );

    \I__6166\ : InMux
    port map (
            O => \N__28514\,
            I => \N__28502\
        );

    \I__6165\ : LocalMux
    port map (
            O => \N__28511\,
            I => \N__28497\
        );

    \I__6164\ : Span12Mux_h
    port map (
            O => \N__28508\,
            I => \N__28497\
        );

    \I__6163\ : Odrv4
    port map (
            O => \N__28505\,
            I => \b2v_inst.N_482\
        );

    \I__6162\ : LocalMux
    port map (
            O => \N__28502\,
            I => \b2v_inst.N_482\
        );

    \I__6161\ : Odrv12
    port map (
            O => \N__28497\,
            I => \b2v_inst.N_482\
        );

    \I__6160\ : CascadeMux
    port map (
            O => \N__28490\,
            I => \N__28487\
        );

    \I__6159\ : InMux
    port map (
            O => \N__28487\,
            I => \N__28484\
        );

    \I__6158\ : LocalMux
    port map (
            O => \N__28484\,
            I => \N__28481\
        );

    \I__6157\ : Span4Mux_h
    port map (
            O => \N__28481\,
            I => \N__28477\
        );

    \I__6156\ : InMux
    port map (
            O => \N__28480\,
            I => \N__28474\
        );

    \I__6155\ : Odrv4
    port map (
            O => \N__28477\,
            I => \b2v_inst.eventosZ0Z_7\
        );

    \I__6154\ : LocalMux
    port map (
            O => \N__28474\,
            I => \b2v_inst.eventosZ0Z_7\
        );

    \I__6153\ : InMux
    port map (
            O => \N__28469\,
            I => \N__28466\
        );

    \I__6152\ : LocalMux
    port map (
            O => \N__28466\,
            I => \b2v_inst.data_a_escribir_RNO_2Z0Z_7\
        );

    \I__6151\ : InMux
    port map (
            O => \N__28463\,
            I => \b2v_inst9.un1_cycle_counter_2_cry_0\
        );

    \I__6150\ : InMux
    port map (
            O => \N__28460\,
            I => \b2v_inst9.un1_cycle_counter_2_cry_1\
        );

    \I__6149\ : InMux
    port map (
            O => \N__28457\,
            I => \b2v_inst9.un1_cycle_counter_2_cry_2\
        );

    \I__6148\ : CascadeMux
    port map (
            O => \N__28454\,
            I => \N__28449\
        );

    \I__6147\ : InMux
    port map (
            O => \N__28453\,
            I => \N__28446\
        );

    \I__6146\ : InMux
    port map (
            O => \N__28452\,
            I => \N__28441\
        );

    \I__6145\ : InMux
    port map (
            O => \N__28449\,
            I => \N__28441\
        );

    \I__6144\ : LocalMux
    port map (
            O => \N__28446\,
            I => \b2v_inst9.cycle_counterZ0Z_3\
        );

    \I__6143\ : LocalMux
    port map (
            O => \N__28441\,
            I => \b2v_inst9.cycle_counterZ0Z_3\
        );

    \I__6142\ : CascadeMux
    port map (
            O => \N__28436\,
            I => \b2v_inst9.cycle_counter_RNIQAGDZ0Z_3_cascade_\
        );

    \I__6141\ : InMux
    port map (
            O => \N__28433\,
            I => \N__28430\
        );

    \I__6140\ : LocalMux
    port map (
            O => \N__28430\,
            I => \b2v_inst9.un1_cycle_counter_2_cry_0_THRU_CO\
        );

    \I__6139\ : CascadeMux
    port map (
            O => \N__28427\,
            I => \N__28422\
        );

    \I__6138\ : CascadeMux
    port map (
            O => \N__28426\,
            I => \N__28419\
        );

    \I__6137\ : InMux
    port map (
            O => \N__28425\,
            I => \N__28409\
        );

    \I__6136\ : InMux
    port map (
            O => \N__28422\,
            I => \N__28409\
        );

    \I__6135\ : InMux
    port map (
            O => \N__28419\,
            I => \N__28409\
        );

    \I__6134\ : InMux
    port map (
            O => \N__28418\,
            I => \N__28409\
        );

    \I__6133\ : LocalMux
    port map (
            O => \N__28409\,
            I => \b2v_inst9.cycle_counterZ0Z_1\
        );

    \I__6132\ : CascadeMux
    port map (
            O => \N__28406\,
            I => \N__28402\
        );

    \I__6131\ : CascadeMux
    port map (
            O => \N__28405\,
            I => \N__28399\
        );

    \I__6130\ : InMux
    port map (
            O => \N__28402\,
            I => \N__28396\
        );

    \I__6129\ : InMux
    port map (
            O => \N__28399\,
            I => \N__28393\
        );

    \I__6128\ : LocalMux
    port map (
            O => \N__28396\,
            I => \N__28390\
        );

    \I__6127\ : LocalMux
    port map (
            O => \N__28393\,
            I => \b2v_inst.reg_anterior_i_9\
        );

    \I__6126\ : Odrv4
    port map (
            O => \N__28390\,
            I => \b2v_inst.reg_anterior_i_9\
        );

    \I__6125\ : CascadeMux
    port map (
            O => \N__28385\,
            I => \N__28381\
        );

    \I__6124\ : CascadeMux
    port map (
            O => \N__28384\,
            I => \N__28378\
        );

    \I__6123\ : InMux
    port map (
            O => \N__28381\,
            I => \N__28375\
        );

    \I__6122\ : InMux
    port map (
            O => \N__28378\,
            I => \N__28372\
        );

    \I__6121\ : LocalMux
    port map (
            O => \N__28375\,
            I => \N__28369\
        );

    \I__6120\ : LocalMux
    port map (
            O => \N__28372\,
            I => \b2v_inst.reg_anterior_i_10\
        );

    \I__6119\ : Odrv4
    port map (
            O => \N__28369\,
            I => \b2v_inst.reg_anterior_i_10\
        );

    \I__6118\ : InMux
    port map (
            O => \N__28364\,
            I => \N__28361\
        );

    \I__6117\ : LocalMux
    port map (
            O => \N__28361\,
            I => \N__28358\
        );

    \I__6116\ : Odrv4
    port map (
            O => \N__28358\,
            I => \b2v_inst.valor_max_final43_THRU_CO\
        );

    \I__6115\ : CascadeMux
    port map (
            O => \N__28355\,
            I => \N__28352\
        );

    \I__6114\ : InMux
    port map (
            O => \N__28352\,
            I => \N__28349\
        );

    \I__6113\ : LocalMux
    port map (
            O => \N__28349\,
            I => \N__28346\
        );

    \I__6112\ : Odrv12
    port map (
            O => \N__28346\,
            I => \b2v_inst.m54_ns_1\
        );

    \I__6111\ : InMux
    port map (
            O => \N__28343\,
            I => \b2v_inst.valor_max_final41\
        );

    \I__6110\ : InMux
    port map (
            O => \N__28340\,
            I => \N__28334\
        );

    \I__6109\ : InMux
    port map (
            O => \N__28339\,
            I => \N__28328\
        );

    \I__6108\ : InMux
    port map (
            O => \N__28338\,
            I => \N__28325\
        );

    \I__6107\ : InMux
    port map (
            O => \N__28337\,
            I => \N__28322\
        );

    \I__6106\ : LocalMux
    port map (
            O => \N__28334\,
            I => \N__28319\
        );

    \I__6105\ : InMux
    port map (
            O => \N__28333\,
            I => \N__28314\
        );

    \I__6104\ : InMux
    port map (
            O => \N__28332\,
            I => \N__28314\
        );

    \I__6103\ : InMux
    port map (
            O => \N__28331\,
            I => \N__28310\
        );

    \I__6102\ : LocalMux
    port map (
            O => \N__28328\,
            I => \N__28307\
        );

    \I__6101\ : LocalMux
    port map (
            O => \N__28325\,
            I => \N__28304\
        );

    \I__6100\ : LocalMux
    port map (
            O => \N__28322\,
            I => \N__28301\
        );

    \I__6099\ : Span4Mux_h
    port map (
            O => \N__28319\,
            I => \N__28298\
        );

    \I__6098\ : LocalMux
    port map (
            O => \N__28314\,
            I => \N__28294\
        );

    \I__6097\ : InMux
    port map (
            O => \N__28313\,
            I => \N__28290\
        );

    \I__6096\ : LocalMux
    port map (
            O => \N__28310\,
            I => \N__28287\
        );

    \I__6095\ : Span4Mux_h
    port map (
            O => \N__28307\,
            I => \N__28282\
        );

    \I__6094\ : Span4Mux_h
    port map (
            O => \N__28304\,
            I => \N__28282\
        );

    \I__6093\ : Span4Mux_h
    port map (
            O => \N__28301\,
            I => \N__28277\
        );

    \I__6092\ : Span4Mux_h
    port map (
            O => \N__28298\,
            I => \N__28277\
        );

    \I__6091\ : InMux
    port map (
            O => \N__28297\,
            I => \N__28274\
        );

    \I__6090\ : Span4Mux_h
    port map (
            O => \N__28294\,
            I => \N__28271\
        );

    \I__6089\ : InMux
    port map (
            O => \N__28293\,
            I => \N__28268\
        );

    \I__6088\ : LocalMux
    port map (
            O => \N__28290\,
            I => \b2v_inst.stateZ0Z_6\
        );

    \I__6087\ : Odrv12
    port map (
            O => \N__28287\,
            I => \b2v_inst.stateZ0Z_6\
        );

    \I__6086\ : Odrv4
    port map (
            O => \N__28282\,
            I => \b2v_inst.stateZ0Z_6\
        );

    \I__6085\ : Odrv4
    port map (
            O => \N__28277\,
            I => \b2v_inst.stateZ0Z_6\
        );

    \I__6084\ : LocalMux
    port map (
            O => \N__28274\,
            I => \b2v_inst.stateZ0Z_6\
        );

    \I__6083\ : Odrv4
    port map (
            O => \N__28271\,
            I => \b2v_inst.stateZ0Z_6\
        );

    \I__6082\ : LocalMux
    port map (
            O => \N__28268\,
            I => \b2v_inst.stateZ0Z_6\
        );

    \I__6081\ : InMux
    port map (
            O => \N__28253\,
            I => \N__28249\
        );

    \I__6080\ : CascadeMux
    port map (
            O => \N__28252\,
            I => \N__28246\
        );

    \I__6079\ : LocalMux
    port map (
            O => \N__28249\,
            I => \N__28243\
        );

    \I__6078\ : InMux
    port map (
            O => \N__28246\,
            I => \N__28240\
        );

    \I__6077\ : Span4Mux_h
    port map (
            O => \N__28243\,
            I => \N__28235\
        );

    \I__6076\ : LocalMux
    port map (
            O => \N__28240\,
            I => \N__28230\
        );

    \I__6075\ : InMux
    port map (
            O => \N__28239\,
            I => \N__28225\
        );

    \I__6074\ : InMux
    port map (
            O => \N__28238\,
            I => \N__28225\
        );

    \I__6073\ : Span4Mux_h
    port map (
            O => \N__28235\,
            I => \N__28222\
        );

    \I__6072\ : InMux
    port map (
            O => \N__28234\,
            I => \N__28217\
        );

    \I__6071\ : InMux
    port map (
            O => \N__28233\,
            I => \N__28217\
        );

    \I__6070\ : Odrv4
    port map (
            O => \N__28230\,
            I => \b2v_inst.stateZ0Z_10\
        );

    \I__6069\ : LocalMux
    port map (
            O => \N__28225\,
            I => \b2v_inst.stateZ0Z_10\
        );

    \I__6068\ : Odrv4
    port map (
            O => \N__28222\,
            I => \b2v_inst.stateZ0Z_10\
        );

    \I__6067\ : LocalMux
    port map (
            O => \N__28217\,
            I => \b2v_inst.stateZ0Z_10\
        );

    \I__6066\ : InMux
    port map (
            O => \N__28208\,
            I => \N__28198\
        );

    \I__6065\ : InMux
    port map (
            O => \N__28207\,
            I => \N__28192\
        );

    \I__6064\ : InMux
    port map (
            O => \N__28206\,
            I => \N__28192\
        );

    \I__6063\ : InMux
    port map (
            O => \N__28205\,
            I => \N__28189\
        );

    \I__6062\ : InMux
    port map (
            O => \N__28204\,
            I => \N__28186\
        );

    \I__6061\ : InMux
    port map (
            O => \N__28203\,
            I => \N__28178\
        );

    \I__6060\ : InMux
    port map (
            O => \N__28202\,
            I => \N__28178\
        );

    \I__6059\ : CascadeMux
    port map (
            O => \N__28201\,
            I => \N__28175\
        );

    \I__6058\ : LocalMux
    port map (
            O => \N__28198\,
            I => \N__28170\
        );

    \I__6057\ : InMux
    port map (
            O => \N__28197\,
            I => \N__28167\
        );

    \I__6056\ : LocalMux
    port map (
            O => \N__28192\,
            I => \N__28164\
        );

    \I__6055\ : LocalMux
    port map (
            O => \N__28189\,
            I => \N__28161\
        );

    \I__6054\ : LocalMux
    port map (
            O => \N__28186\,
            I => \N__28158\
        );

    \I__6053\ : InMux
    port map (
            O => \N__28185\,
            I => \N__28151\
        );

    \I__6052\ : InMux
    port map (
            O => \N__28184\,
            I => \N__28151\
        );

    \I__6051\ : InMux
    port map (
            O => \N__28183\,
            I => \N__28151\
        );

    \I__6050\ : LocalMux
    port map (
            O => \N__28178\,
            I => \N__28148\
        );

    \I__6049\ : InMux
    port map (
            O => \N__28175\,
            I => \N__28145\
        );

    \I__6048\ : InMux
    port map (
            O => \N__28174\,
            I => \N__28142\
        );

    \I__6047\ : InMux
    port map (
            O => \N__28173\,
            I => \N__28139\
        );

    \I__6046\ : Span4Mux_v
    port map (
            O => \N__28170\,
            I => \N__28133\
        );

    \I__6045\ : LocalMux
    port map (
            O => \N__28167\,
            I => \N__28130\
        );

    \I__6044\ : Span4Mux_h
    port map (
            O => \N__28164\,
            I => \N__28127\
        );

    \I__6043\ : Span4Mux_v
    port map (
            O => \N__28161\,
            I => \N__28116\
        );

    \I__6042\ : Span4Mux_v
    port map (
            O => \N__28158\,
            I => \N__28116\
        );

    \I__6041\ : LocalMux
    port map (
            O => \N__28151\,
            I => \N__28116\
        );

    \I__6040\ : Span4Mux_h
    port map (
            O => \N__28148\,
            I => \N__28116\
        );

    \I__6039\ : LocalMux
    port map (
            O => \N__28145\,
            I => \N__28116\
        );

    \I__6038\ : LocalMux
    port map (
            O => \N__28142\,
            I => \N__28113\
        );

    \I__6037\ : LocalMux
    port map (
            O => \N__28139\,
            I => \N__28110\
        );

    \I__6036\ : InMux
    port map (
            O => \N__28138\,
            I => \N__28107\
        );

    \I__6035\ : InMux
    port map (
            O => \N__28137\,
            I => \N__28102\
        );

    \I__6034\ : InMux
    port map (
            O => \N__28136\,
            I => \N__28102\
        );

    \I__6033\ : Span4Mux_h
    port map (
            O => \N__28133\,
            I => \N__28099\
        );

    \I__6032\ : Span4Mux_h
    port map (
            O => \N__28130\,
            I => \N__28096\
        );

    \I__6031\ : Span4Mux_h
    port map (
            O => \N__28127\,
            I => \N__28091\
        );

    \I__6030\ : Span4Mux_h
    port map (
            O => \N__28116\,
            I => \N__28091\
        );

    \I__6029\ : Odrv12
    port map (
            O => \N__28113\,
            I => \b2v_inst.stateZ0Z_29\
        );

    \I__6028\ : Odrv4
    port map (
            O => \N__28110\,
            I => \b2v_inst.stateZ0Z_29\
        );

    \I__6027\ : LocalMux
    port map (
            O => \N__28107\,
            I => \b2v_inst.stateZ0Z_29\
        );

    \I__6026\ : LocalMux
    port map (
            O => \N__28102\,
            I => \b2v_inst.stateZ0Z_29\
        );

    \I__6025\ : Odrv4
    port map (
            O => \N__28099\,
            I => \b2v_inst.stateZ0Z_29\
        );

    \I__6024\ : Odrv4
    port map (
            O => \N__28096\,
            I => \b2v_inst.stateZ0Z_29\
        );

    \I__6023\ : Odrv4
    port map (
            O => \N__28091\,
            I => \b2v_inst.stateZ0Z_29\
        );

    \I__6022\ : InMux
    port map (
            O => \N__28076\,
            I => \N__28073\
        );

    \I__6021\ : LocalMux
    port map (
            O => \N__28073\,
            I => \N__28070\
        );

    \I__6020\ : Odrv4
    port map (
            O => \N__28070\,
            I => \b2v_inst.state_ns_a3_i_0_a2_1_4_1\
        );

    \I__6019\ : CascadeMux
    port map (
            O => \N__28067\,
            I => \N__28061\
        );

    \I__6018\ : InMux
    port map (
            O => \N__28066\,
            I => \N__28058\
        );

    \I__6017\ : InMux
    port map (
            O => \N__28065\,
            I => \N__28053\
        );

    \I__6016\ : InMux
    port map (
            O => \N__28064\,
            I => \N__28053\
        );

    \I__6015\ : InMux
    port map (
            O => \N__28061\,
            I => \N__28050\
        );

    \I__6014\ : LocalMux
    port map (
            O => \N__28058\,
            I => \N__28047\
        );

    \I__6013\ : LocalMux
    port map (
            O => \N__28053\,
            I => \N__28040\
        );

    \I__6012\ : LocalMux
    port map (
            O => \N__28050\,
            I => \N__28040\
        );

    \I__6011\ : Span4Mux_h
    port map (
            O => \N__28047\,
            I => \N__28037\
        );

    \I__6010\ : InMux
    port map (
            O => \N__28046\,
            I => \N__28032\
        );

    \I__6009\ : InMux
    port map (
            O => \N__28045\,
            I => \N__28032\
        );

    \I__6008\ : Odrv12
    port map (
            O => \N__28040\,
            I => b2v_inst_state_3
        );

    \I__6007\ : Odrv4
    port map (
            O => \N__28037\,
            I => b2v_inst_state_3
        );

    \I__6006\ : LocalMux
    port map (
            O => \N__28032\,
            I => b2v_inst_state_3
        );

    \I__6005\ : InMux
    port map (
            O => \N__28025\,
            I => \N__28022\
        );

    \I__6004\ : LocalMux
    port map (
            O => \N__28022\,
            I => \b2v_inst.N_694\
        );

    \I__6003\ : CascadeMux
    port map (
            O => \N__28019\,
            I => \b2v_inst.N_695_cascade_\
        );

    \I__6002\ : InMux
    port map (
            O => \N__28016\,
            I => \N__28013\
        );

    \I__6001\ : LocalMux
    port map (
            O => \N__28013\,
            I => \N__28010\
        );

    \I__6000\ : Span4Mux_h
    port map (
            O => \N__28010\,
            I => \N__28007\
        );

    \I__5999\ : Odrv4
    port map (
            O => \N__28007\,
            I => \b2v_inst.state_ns_a3_i_0_1_1\
        );

    \I__5998\ : InMux
    port map (
            O => \N__28004\,
            I => \N__27998\
        );

    \I__5997\ : InMux
    port map (
            O => \N__28003\,
            I => \N__27998\
        );

    \I__5996\ : LocalMux
    port map (
            O => \N__27998\,
            I => \N__27994\
        );

    \I__5995\ : InMux
    port map (
            O => \N__27997\,
            I => \N__27990\
        );

    \I__5994\ : Span4Mux_h
    port map (
            O => \N__27994\,
            I => \N__27987\
        );

    \I__5993\ : InMux
    port map (
            O => \N__27993\,
            I => \N__27984\
        );

    \I__5992\ : LocalMux
    port map (
            O => \N__27990\,
            I => \N__27980\
        );

    \I__5991\ : Span4Mux_h
    port map (
            O => \N__27987\,
            I => \N__27975\
        );

    \I__5990\ : LocalMux
    port map (
            O => \N__27984\,
            I => \N__27975\
        );

    \I__5989\ : InMux
    port map (
            O => \N__27983\,
            I => \N__27972\
        );

    \I__5988\ : Span4Mux_v
    port map (
            O => \N__27980\,
            I => \N__27967\
        );

    \I__5987\ : Span4Mux_h
    port map (
            O => \N__27975\,
            I => \N__27967\
        );

    \I__5986\ : LocalMux
    port map (
            O => \N__27972\,
            I => \b2v_inst.un2_cuentalto10_i_a2_8\
        );

    \I__5985\ : Odrv4
    port map (
            O => \N__27967\,
            I => \b2v_inst.un2_cuentalto10_i_a2_8\
        );

    \I__5984\ : InMux
    port map (
            O => \N__27962\,
            I => \N__27954\
        );

    \I__5983\ : InMux
    port map (
            O => \N__27961\,
            I => \N__27954\
        );

    \I__5982\ : InMux
    port map (
            O => \N__27960\,
            I => \N__27951\
        );

    \I__5981\ : InMux
    port map (
            O => \N__27959\,
            I => \N__27947\
        );

    \I__5980\ : LocalMux
    port map (
            O => \N__27954\,
            I => \N__27944\
        );

    \I__5979\ : LocalMux
    port map (
            O => \N__27951\,
            I => \N__27941\
        );

    \I__5978\ : InMux
    port map (
            O => \N__27950\,
            I => \N__27938\
        );

    \I__5977\ : LocalMux
    port map (
            O => \N__27947\,
            I => \N__27935\
        );

    \I__5976\ : Span4Mux_h
    port map (
            O => \N__27944\,
            I => \N__27932\
        );

    \I__5975\ : Span4Mux_v
    port map (
            O => \N__27941\,
            I => \N__27925\
        );

    \I__5974\ : LocalMux
    port map (
            O => \N__27938\,
            I => \N__27925\
        );

    \I__5973\ : Span4Mux_h
    port map (
            O => \N__27935\,
            I => \N__27925\
        );

    \I__5972\ : Odrv4
    port map (
            O => \N__27932\,
            I => \b2v_inst.un2_cuentalto10_i_a2_7\
        );

    \I__5971\ : Odrv4
    port map (
            O => \N__27925\,
            I => \b2v_inst.un2_cuentalto10_i_a2_7\
        );

    \I__5970\ : CascadeMux
    port map (
            O => \N__27920\,
            I => \N__27914\
        );

    \I__5969\ : InMux
    port map (
            O => \N__27919\,
            I => \N__27911\
        );

    \I__5968\ : InMux
    port map (
            O => \N__27918\,
            I => \N__27902\
        );

    \I__5967\ : InMux
    port map (
            O => \N__27917\,
            I => \N__27902\
        );

    \I__5966\ : InMux
    port map (
            O => \N__27914\,
            I => \N__27902\
        );

    \I__5965\ : LocalMux
    port map (
            O => \N__27911\,
            I => \N__27899\
        );

    \I__5964\ : InMux
    port map (
            O => \N__27910\,
            I => \N__27896\
        );

    \I__5963\ : CascadeMux
    port map (
            O => \N__27909\,
            I => \N__27893\
        );

    \I__5962\ : LocalMux
    port map (
            O => \N__27902\,
            I => \N__27890\
        );

    \I__5961\ : Span4Mux_h
    port map (
            O => \N__27899\,
            I => \N__27887\
        );

    \I__5960\ : LocalMux
    port map (
            O => \N__27896\,
            I => \N__27883\
        );

    \I__5959\ : InMux
    port map (
            O => \N__27893\,
            I => \N__27880\
        );

    \I__5958\ : Span4Mux_v
    port map (
            O => \N__27890\,
            I => \N__27877\
        );

    \I__5957\ : Span4Mux_v
    port map (
            O => \N__27887\,
            I => \N__27874\
        );

    \I__5956\ : InMux
    port map (
            O => \N__27886\,
            I => \N__27871\
        );

    \I__5955\ : Span4Mux_v
    port map (
            O => \N__27883\,
            I => \N__27866\
        );

    \I__5954\ : LocalMux
    port map (
            O => \N__27880\,
            I => \N__27866\
        );

    \I__5953\ : Sp12to4
    port map (
            O => \N__27877\,
            I => \N__27859\
        );

    \I__5952\ : Sp12to4
    port map (
            O => \N__27874\,
            I => \N__27859\
        );

    \I__5951\ : LocalMux
    port map (
            O => \N__27871\,
            I => \N__27859\
        );

    \I__5950\ : Span4Mux_h
    port map (
            O => \N__27866\,
            I => \N__27856\
        );

    \I__5949\ : Span12Mux_h
    port map (
            O => \N__27859\,
            I => \N__27853\
        );

    \I__5948\ : Span4Mux_h
    port map (
            O => \N__27856\,
            I => \N__27850\
        );

    \I__5947\ : Odrv12
    port map (
            O => \N__27853\,
            I => \b2v_inst.state_32_repZ0Z1\
        );

    \I__5946\ : Odrv4
    port map (
            O => \N__27850\,
            I => \b2v_inst.state_32_repZ0Z1\
        );

    \I__5945\ : CascadeMux
    port map (
            O => \N__27845\,
            I => \N__27841\
        );

    \I__5944\ : InMux
    port map (
            O => \N__27844\,
            I => \N__27834\
        );

    \I__5943\ : InMux
    port map (
            O => \N__27841\,
            I => \N__27830\
        );

    \I__5942\ : InMux
    port map (
            O => \N__27840\,
            I => \N__27827\
        );

    \I__5941\ : InMux
    port map (
            O => \N__27839\,
            I => \N__27822\
        );

    \I__5940\ : InMux
    port map (
            O => \N__27838\,
            I => \N__27822\
        );

    \I__5939\ : InMux
    port map (
            O => \N__27837\,
            I => \N__27819\
        );

    \I__5938\ : LocalMux
    port map (
            O => \N__27834\,
            I => \N__27816\
        );

    \I__5937\ : InMux
    port map (
            O => \N__27833\,
            I => \N__27813\
        );

    \I__5936\ : LocalMux
    port map (
            O => \N__27830\,
            I => \N__27808\
        );

    \I__5935\ : LocalMux
    port map (
            O => \N__27827\,
            I => \N__27808\
        );

    \I__5934\ : LocalMux
    port map (
            O => \N__27822\,
            I => \N__27805\
        );

    \I__5933\ : LocalMux
    port map (
            O => \N__27819\,
            I => \N__27802\
        );

    \I__5932\ : Span4Mux_v
    port map (
            O => \N__27816\,
            I => \N__27799\
        );

    \I__5931\ : LocalMux
    port map (
            O => \N__27813\,
            I => \N__27796\
        );

    \I__5930\ : Span4Mux_v
    port map (
            O => \N__27808\,
            I => \N__27793\
        );

    \I__5929\ : Span4Mux_h
    port map (
            O => \N__27805\,
            I => \N__27788\
        );

    \I__5928\ : Span4Mux_v
    port map (
            O => \N__27802\,
            I => \N__27788\
        );

    \I__5927\ : Span4Mux_v
    port map (
            O => \N__27799\,
            I => \N__27782\
        );

    \I__5926\ : Span4Mux_v
    port map (
            O => \N__27796\,
            I => \N__27782\
        );

    \I__5925\ : Span4Mux_v
    port map (
            O => \N__27793\,
            I => \N__27779\
        );

    \I__5924\ : Span4Mux_h
    port map (
            O => \N__27788\,
            I => \N__27776\
        );

    \I__5923\ : InMux
    port map (
            O => \N__27787\,
            I => \N__27773\
        );

    \I__5922\ : Sp12to4
    port map (
            O => \N__27782\,
            I => \N__27768\
        );

    \I__5921\ : Sp12to4
    port map (
            O => \N__27779\,
            I => \N__27768\
        );

    \I__5920\ : Span4Mux_h
    port map (
            O => \N__27776\,
            I => \N__27763\
        );

    \I__5919\ : LocalMux
    port map (
            O => \N__27773\,
            I => \N__27763\
        );

    \I__5918\ : Span12Mux_h
    port map (
            O => \N__27768\,
            I => \N__27760\
        );

    \I__5917\ : Sp12to4
    port map (
            O => \N__27763\,
            I => \N__27757\
        );

    \I__5916\ : Span12Mux_v
    port map (
            O => \N__27760\,
            I => \N__27754\
        );

    \I__5915\ : Span12Mux_v
    port map (
            O => \N__27757\,
            I => \N__27751\
        );

    \I__5914\ : Odrv12
    port map (
            O => \N__27754\,
            I => reset_c
        );

    \I__5913\ : Odrv12
    port map (
            O => \N__27751\,
            I => reset_c
        );

    \I__5912\ : CascadeMux
    port map (
            O => \N__27746\,
            I => \N__27742\
        );

    \I__5911\ : InMux
    port map (
            O => \N__27745\,
            I => \N__27739\
        );

    \I__5910\ : InMux
    port map (
            O => \N__27742\,
            I => \N__27736\
        );

    \I__5909\ : LocalMux
    port map (
            O => \N__27739\,
            I => \N__27733\
        );

    \I__5908\ : LocalMux
    port map (
            O => \N__27736\,
            I => \b2v_inst.reg_anterior_i_1\
        );

    \I__5907\ : Odrv4
    port map (
            O => \N__27733\,
            I => \b2v_inst.reg_anterior_i_1\
        );

    \I__5906\ : CascadeMux
    port map (
            O => \N__27728\,
            I => \N__27724\
        );

    \I__5905\ : InMux
    port map (
            O => \N__27727\,
            I => \N__27721\
        );

    \I__5904\ : InMux
    port map (
            O => \N__27724\,
            I => \N__27718\
        );

    \I__5903\ : LocalMux
    port map (
            O => \N__27721\,
            I => \N__27715\
        );

    \I__5902\ : LocalMux
    port map (
            O => \N__27718\,
            I => \b2v_inst.reg_anterior_i_2\
        );

    \I__5901\ : Odrv4
    port map (
            O => \N__27715\,
            I => \b2v_inst.reg_anterior_i_2\
        );

    \I__5900\ : CascadeMux
    port map (
            O => \N__27710\,
            I => \N__27706\
        );

    \I__5899\ : InMux
    port map (
            O => \N__27709\,
            I => \N__27703\
        );

    \I__5898\ : InMux
    port map (
            O => \N__27706\,
            I => \N__27700\
        );

    \I__5897\ : LocalMux
    port map (
            O => \N__27703\,
            I => \N__27697\
        );

    \I__5896\ : LocalMux
    port map (
            O => \N__27700\,
            I => \b2v_inst.reg_anterior_i_3\
        );

    \I__5895\ : Odrv4
    port map (
            O => \N__27697\,
            I => \b2v_inst.reg_anterior_i_3\
        );

    \I__5894\ : CascadeMux
    port map (
            O => \N__27692\,
            I => \N__27688\
        );

    \I__5893\ : CascadeMux
    port map (
            O => \N__27691\,
            I => \N__27685\
        );

    \I__5892\ : InMux
    port map (
            O => \N__27688\,
            I => \N__27682\
        );

    \I__5891\ : InMux
    port map (
            O => \N__27685\,
            I => \N__27679\
        );

    \I__5890\ : LocalMux
    port map (
            O => \N__27682\,
            I => \N__27676\
        );

    \I__5889\ : LocalMux
    port map (
            O => \N__27679\,
            I => \b2v_inst.reg_anterior_i_4\
        );

    \I__5888\ : Odrv4
    port map (
            O => \N__27676\,
            I => \b2v_inst.reg_anterior_i_4\
        );

    \I__5887\ : CascadeMux
    port map (
            O => \N__27671\,
            I => \N__27667\
        );

    \I__5886\ : CascadeMux
    port map (
            O => \N__27670\,
            I => \N__27664\
        );

    \I__5885\ : InMux
    port map (
            O => \N__27667\,
            I => \N__27661\
        );

    \I__5884\ : InMux
    port map (
            O => \N__27664\,
            I => \N__27658\
        );

    \I__5883\ : LocalMux
    port map (
            O => \N__27661\,
            I => \N__27655\
        );

    \I__5882\ : LocalMux
    port map (
            O => \N__27658\,
            I => \b2v_inst.reg_anterior_i_5\
        );

    \I__5881\ : Odrv4
    port map (
            O => \N__27655\,
            I => \b2v_inst.reg_anterior_i_5\
        );

    \I__5880\ : CascadeMux
    port map (
            O => \N__27650\,
            I => \N__27646\
        );

    \I__5879\ : InMux
    port map (
            O => \N__27649\,
            I => \N__27643\
        );

    \I__5878\ : InMux
    port map (
            O => \N__27646\,
            I => \N__27640\
        );

    \I__5877\ : LocalMux
    port map (
            O => \N__27643\,
            I => \N__27637\
        );

    \I__5876\ : LocalMux
    port map (
            O => \N__27640\,
            I => \b2v_inst.reg_anterior_i_6\
        );

    \I__5875\ : Odrv4
    port map (
            O => \N__27637\,
            I => \b2v_inst.reg_anterior_i_6\
        );

    \I__5874\ : CascadeMux
    port map (
            O => \N__27632\,
            I => \N__27628\
        );

    \I__5873\ : CascadeMux
    port map (
            O => \N__27631\,
            I => \N__27625\
        );

    \I__5872\ : InMux
    port map (
            O => \N__27628\,
            I => \N__27622\
        );

    \I__5871\ : InMux
    port map (
            O => \N__27625\,
            I => \N__27619\
        );

    \I__5870\ : LocalMux
    port map (
            O => \N__27622\,
            I => \N__27616\
        );

    \I__5869\ : LocalMux
    port map (
            O => \N__27619\,
            I => \b2v_inst.reg_anterior_i_7\
        );

    \I__5868\ : Odrv4
    port map (
            O => \N__27616\,
            I => \b2v_inst.reg_anterior_i_7\
        );

    \I__5867\ : CascadeMux
    port map (
            O => \N__27611\,
            I => \N__27607\
        );

    \I__5866\ : CascadeMux
    port map (
            O => \N__27610\,
            I => \N__27604\
        );

    \I__5865\ : InMux
    port map (
            O => \N__27607\,
            I => \N__27601\
        );

    \I__5864\ : InMux
    port map (
            O => \N__27604\,
            I => \N__27598\
        );

    \I__5863\ : LocalMux
    port map (
            O => \N__27601\,
            I => \N__27595\
        );

    \I__5862\ : LocalMux
    port map (
            O => \N__27598\,
            I => \b2v_inst.reg_anterior_i_8\
        );

    \I__5861\ : Odrv4
    port map (
            O => \N__27595\,
            I => \b2v_inst.reg_anterior_i_8\
        );

    \I__5860\ : CascadeMux
    port map (
            O => \N__27590\,
            I => \N__27587\
        );

    \I__5859\ : InMux
    port map (
            O => \N__27587\,
            I => \N__27582\
        );

    \I__5858\ : InMux
    port map (
            O => \N__27586\,
            I => \N__27579\
        );

    \I__5857\ : InMux
    port map (
            O => \N__27585\,
            I => \N__27576\
        );

    \I__5856\ : LocalMux
    port map (
            O => \N__27582\,
            I => \N__27572\
        );

    \I__5855\ : LocalMux
    port map (
            O => \N__27579\,
            I => \N__27569\
        );

    \I__5854\ : LocalMux
    port map (
            O => \N__27576\,
            I => \N__27566\
        );

    \I__5853\ : InMux
    port map (
            O => \N__27575\,
            I => \N__27563\
        );

    \I__5852\ : Span4Mux_h
    port map (
            O => \N__27572\,
            I => \N__27559\
        );

    \I__5851\ : Span4Mux_v
    port map (
            O => \N__27569\,
            I => \N__27552\
        );

    \I__5850\ : Span4Mux_h
    port map (
            O => \N__27566\,
            I => \N__27552\
        );

    \I__5849\ : LocalMux
    port map (
            O => \N__27563\,
            I => \N__27552\
        );

    \I__5848\ : InMux
    port map (
            O => \N__27562\,
            I => \N__27549\
        );

    \I__5847\ : Odrv4
    port map (
            O => \N__27559\,
            I => \b2v_inst.reg_ancho_2Z0Z_7\
        );

    \I__5846\ : Odrv4
    port map (
            O => \N__27552\,
            I => \b2v_inst.reg_ancho_2Z0Z_7\
        );

    \I__5845\ : LocalMux
    port map (
            O => \N__27549\,
            I => \b2v_inst.reg_ancho_2Z0Z_7\
        );

    \I__5844\ : InMux
    port map (
            O => \N__27542\,
            I => \b2v_inst.valor_max_final43\
        );

    \I__5843\ : InMux
    port map (
            O => \N__27539\,
            I => \N__27536\
        );

    \I__5842\ : LocalMux
    port map (
            O => \N__27536\,
            I => \b2v_inst.data_a_escribir_RNO_0Z0Z_0\
        );

    \I__5841\ : InMux
    port map (
            O => \N__27533\,
            I => \N__27530\
        );

    \I__5840\ : LocalMux
    port map (
            O => \N__27530\,
            I => \b2v_inst.data_a_escribir_RNO_0Z0Z_1\
        );

    \I__5839\ : InMux
    port map (
            O => \N__27527\,
            I => \N__27524\
        );

    \I__5838\ : LocalMux
    port map (
            O => \N__27524\,
            I => \N__27521\
        );

    \I__5837\ : Span4Mux_v
    port map (
            O => \N__27521\,
            I => \N__27517\
        );

    \I__5836\ : InMux
    port map (
            O => \N__27520\,
            I => \N__27514\
        );

    \I__5835\ : Sp12to4
    port map (
            O => \N__27517\,
            I => \N__27511\
        );

    \I__5834\ : LocalMux
    port map (
            O => \N__27514\,
            I => \b2v_inst.eventosZ0Z_5\
        );

    \I__5833\ : Odrv12
    port map (
            O => \N__27511\,
            I => \b2v_inst.eventosZ0Z_5\
        );

    \I__5832\ : CascadeMux
    port map (
            O => \N__27506\,
            I => \N__27502\
        );

    \I__5831\ : InMux
    port map (
            O => \N__27505\,
            I => \N__27499\
        );

    \I__5830\ : InMux
    port map (
            O => \N__27502\,
            I => \N__27496\
        );

    \I__5829\ : LocalMux
    port map (
            O => \N__27499\,
            I => \N__27493\
        );

    \I__5828\ : LocalMux
    port map (
            O => \N__27496\,
            I => \b2v_inst.reg_anterior_i_0\
        );

    \I__5827\ : Odrv4
    port map (
            O => \N__27493\,
            I => \b2v_inst.reg_anterior_i_0\
        );

    \I__5826\ : InMux
    port map (
            O => \N__27488\,
            I => \N__27483\
        );

    \I__5825\ : InMux
    port map (
            O => \N__27487\,
            I => \N__27480\
        );

    \I__5824\ : InMux
    port map (
            O => \N__27486\,
            I => \N__27476\
        );

    \I__5823\ : LocalMux
    port map (
            O => \N__27483\,
            I => \N__27471\
        );

    \I__5822\ : LocalMux
    port map (
            O => \N__27480\,
            I => \N__27471\
        );

    \I__5821\ : InMux
    port map (
            O => \N__27479\,
            I => \N__27468\
        );

    \I__5820\ : LocalMux
    port map (
            O => \N__27476\,
            I => \N__27465\
        );

    \I__5819\ : Span4Mux_v
    port map (
            O => \N__27471\,
            I => \N__27460\
        );

    \I__5818\ : LocalMux
    port map (
            O => \N__27468\,
            I => \N__27460\
        );

    \I__5817\ : Span4Mux_v
    port map (
            O => \N__27465\,
            I => \N__27455\
        );

    \I__5816\ : Span4Mux_h
    port map (
            O => \N__27460\,
            I => \N__27455\
        );

    \I__5815\ : Span4Mux_h
    port map (
            O => \N__27455\,
            I => \N__27452\
        );

    \I__5814\ : Odrv4
    port map (
            O => \N__27452\,
            I => \SYNTHESIZED_WIRE_3_0\
        );

    \I__5813\ : InMux
    port map (
            O => \N__27449\,
            I => \N__27445\
        );

    \I__5812\ : CascadeMux
    port map (
            O => \N__27448\,
            I => \N__27442\
        );

    \I__5811\ : LocalMux
    port map (
            O => \N__27445\,
            I => \N__27438\
        );

    \I__5810\ : InMux
    port map (
            O => \N__27442\,
            I => \N__27435\
        );

    \I__5809\ : CascadeMux
    port map (
            O => \N__27441\,
            I => \N__27431\
        );

    \I__5808\ : Span4Mux_v
    port map (
            O => \N__27438\,
            I => \N__27425\
        );

    \I__5807\ : LocalMux
    port map (
            O => \N__27435\,
            I => \N__27425\
        );

    \I__5806\ : CascadeMux
    port map (
            O => \N__27434\,
            I => \N__27422\
        );

    \I__5805\ : InMux
    port map (
            O => \N__27431\,
            I => \N__27419\
        );

    \I__5804\ : InMux
    port map (
            O => \N__27430\,
            I => \N__27416\
        );

    \I__5803\ : Span4Mux_v
    port map (
            O => \N__27425\,
            I => \N__27413\
        );

    \I__5802\ : InMux
    port map (
            O => \N__27422\,
            I => \N__27410\
        );

    \I__5801\ : LocalMux
    port map (
            O => \N__27419\,
            I => \N__27405\
        );

    \I__5800\ : LocalMux
    port map (
            O => \N__27416\,
            I => \N__27405\
        );

    \I__5799\ : Odrv4
    port map (
            O => \N__27413\,
            I => \b2v_inst.reg_ancho_2Z0Z_0\
        );

    \I__5798\ : LocalMux
    port map (
            O => \N__27410\,
            I => \b2v_inst.reg_ancho_2Z0Z_0\
        );

    \I__5797\ : Odrv4
    port map (
            O => \N__27405\,
            I => \b2v_inst.reg_ancho_2Z0Z_0\
        );

    \I__5796\ : InMux
    port map (
            O => \N__27398\,
            I => \N__27395\
        );

    \I__5795\ : LocalMux
    port map (
            O => \N__27395\,
            I => \N__27390\
        );

    \I__5794\ : CascadeMux
    port map (
            O => \N__27394\,
            I => \N__27387\
        );

    \I__5793\ : InMux
    port map (
            O => \N__27393\,
            I => \N__27384\
        );

    \I__5792\ : Span4Mux_v
    port map (
            O => \N__27390\,
            I => \N__27380\
        );

    \I__5791\ : InMux
    port map (
            O => \N__27387\,
            I => \N__27377\
        );

    \I__5790\ : LocalMux
    port map (
            O => \N__27384\,
            I => \N__27374\
        );

    \I__5789\ : InMux
    port map (
            O => \N__27383\,
            I => \N__27371\
        );

    \I__5788\ : Span4Mux_h
    port map (
            O => \N__27380\,
            I => \N__27365\
        );

    \I__5787\ : LocalMux
    port map (
            O => \N__27377\,
            I => \N__27365\
        );

    \I__5786\ : Span4Mux_h
    port map (
            O => \N__27374\,
            I => \N__27360\
        );

    \I__5785\ : LocalMux
    port map (
            O => \N__27371\,
            I => \N__27360\
        );

    \I__5784\ : InMux
    port map (
            O => \N__27370\,
            I => \N__27357\
        );

    \I__5783\ : Odrv4
    port map (
            O => \N__27365\,
            I => \b2v_inst.reg_ancho_2Z0Z_5\
        );

    \I__5782\ : Odrv4
    port map (
            O => \N__27360\,
            I => \b2v_inst.reg_ancho_2Z0Z_5\
        );

    \I__5781\ : LocalMux
    port map (
            O => \N__27357\,
            I => \b2v_inst.reg_ancho_2Z0Z_5\
        );

    \I__5780\ : InMux
    port map (
            O => \N__27350\,
            I => \N__27345\
        );

    \I__5779\ : CascadeMux
    port map (
            O => \N__27349\,
            I => \N__27342\
        );

    \I__5778\ : CascadeMux
    port map (
            O => \N__27348\,
            I => \N__27339\
        );

    \I__5777\ : LocalMux
    port map (
            O => \N__27345\,
            I => \N__27336\
        );

    \I__5776\ : InMux
    port map (
            O => \N__27342\,
            I => \N__27333\
        );

    \I__5775\ : InMux
    port map (
            O => \N__27339\,
            I => \N__27330\
        );

    \I__5774\ : Span4Mux_h
    port map (
            O => \N__27336\,
            I => \N__27327\
        );

    \I__5773\ : LocalMux
    port map (
            O => \N__27333\,
            I => \N__27324\
        );

    \I__5772\ : LocalMux
    port map (
            O => \N__27330\,
            I => \N__27321\
        );

    \I__5771\ : Span4Mux_v
    port map (
            O => \N__27327\,
            I => \N__27312\
        );

    \I__5770\ : Span4Mux_v
    port map (
            O => \N__27324\,
            I => \N__27312\
        );

    \I__5769\ : Span4Mux_v
    port map (
            O => \N__27321\,
            I => \N__27312\
        );

    \I__5768\ : InMux
    port map (
            O => \N__27320\,
            I => \N__27309\
        );

    \I__5767\ : InMux
    port map (
            O => \N__27319\,
            I => \N__27306\
        );

    \I__5766\ : Odrv4
    port map (
            O => \N__27312\,
            I => \b2v_inst.reg_ancho_2Z0Z_6\
        );

    \I__5765\ : LocalMux
    port map (
            O => \N__27309\,
            I => \b2v_inst.reg_ancho_2Z0Z_6\
        );

    \I__5764\ : LocalMux
    port map (
            O => \N__27306\,
            I => \b2v_inst.reg_ancho_2Z0Z_6\
        );

    \I__5763\ : InMux
    port map (
            O => \N__27299\,
            I => \b2v_inst.valor_max_final42\
        );

    \I__5762\ : InMux
    port map (
            O => \N__27296\,
            I => \N__27293\
        );

    \I__5761\ : LocalMux
    port map (
            O => \N__27293\,
            I => \N__27290\
        );

    \I__5760\ : Span4Mux_h
    port map (
            O => \N__27290\,
            I => \N__27287\
        );

    \I__5759\ : Odrv4
    port map (
            O => \N__27287\,
            I => \b2v_inst.data_a_escribir11_7_and\
        );

    \I__5758\ : InMux
    port map (
            O => \N__27284\,
            I => \N__27280\
        );

    \I__5757\ : InMux
    port map (
            O => \N__27283\,
            I => \N__27277\
        );

    \I__5756\ : LocalMux
    port map (
            O => \N__27280\,
            I => \N__27271\
        );

    \I__5755\ : LocalMux
    port map (
            O => \N__27277\,
            I => \N__27271\
        );

    \I__5754\ : InMux
    port map (
            O => \N__27276\,
            I => \N__27267\
        );

    \I__5753\ : Span4Mux_v
    port map (
            O => \N__27271\,
            I => \N__27264\
        );

    \I__5752\ : InMux
    port map (
            O => \N__27270\,
            I => \N__27261\
        );

    \I__5751\ : LocalMux
    port map (
            O => \N__27267\,
            I => \N__27254\
        );

    \I__5750\ : Sp12to4
    port map (
            O => \N__27264\,
            I => \N__27254\
        );

    \I__5749\ : LocalMux
    port map (
            O => \N__27261\,
            I => \N__27254\
        );

    \I__5748\ : Odrv12
    port map (
            O => \N__27254\,
            I => \SYNTHESIZED_WIRE_3_7\
        );

    \I__5747\ : InMux
    port map (
            O => \N__27251\,
            I => \N__27245\
        );

    \I__5746\ : InMux
    port map (
            O => \N__27250\,
            I => \N__27242\
        );

    \I__5745\ : InMux
    port map (
            O => \N__27249\,
            I => \N__27239\
        );

    \I__5744\ : InMux
    port map (
            O => \N__27248\,
            I => \N__27236\
        );

    \I__5743\ : LocalMux
    port map (
            O => \N__27245\,
            I => \N__27233\
        );

    \I__5742\ : LocalMux
    port map (
            O => \N__27242\,
            I => \N__27228\
        );

    \I__5741\ : LocalMux
    port map (
            O => \N__27239\,
            I => \N__27228\
        );

    \I__5740\ : LocalMux
    port map (
            O => \N__27236\,
            I => \N__27225\
        );

    \I__5739\ : Span4Mux_v
    port map (
            O => \N__27233\,
            I => \N__27222\
        );

    \I__5738\ : Span4Mux_v
    port map (
            O => \N__27228\,
            I => \N__27217\
        );

    \I__5737\ : Span4Mux_h
    port map (
            O => \N__27225\,
            I => \N__27217\
        );

    \I__5736\ : Span4Mux_h
    port map (
            O => \N__27222\,
            I => \N__27214\
        );

    \I__5735\ : Span4Mux_h
    port map (
            O => \N__27217\,
            I => \N__27211\
        );

    \I__5734\ : Odrv4
    port map (
            O => \N__27214\,
            I => \SYNTHESIZED_WIRE_3_8\
        );

    \I__5733\ : Odrv4
    port map (
            O => \N__27211\,
            I => \SYNTHESIZED_WIRE_3_8\
        );

    \I__5732\ : CascadeMux
    port map (
            O => \N__27206\,
            I => \N__27200\
        );

    \I__5731\ : CascadeMux
    port map (
            O => \N__27205\,
            I => \N__27197\
        );

    \I__5730\ : CascadeMux
    port map (
            O => \N__27204\,
            I => \N__27193\
        );

    \I__5729\ : InMux
    port map (
            O => \N__27203\,
            I => \N__27183\
        );

    \I__5728\ : InMux
    port map (
            O => \N__27200\,
            I => \N__27183\
        );

    \I__5727\ : InMux
    port map (
            O => \N__27197\,
            I => \N__27179\
        );

    \I__5726\ : InMux
    port map (
            O => \N__27196\,
            I => \N__27174\
        );

    \I__5725\ : InMux
    port map (
            O => \N__27193\,
            I => \N__27174\
        );

    \I__5724\ : InMux
    port map (
            O => \N__27192\,
            I => \N__27171\
        );

    \I__5723\ : InMux
    port map (
            O => \N__27191\,
            I => \N__27168\
        );

    \I__5722\ : InMux
    port map (
            O => \N__27190\,
            I => \N__27163\
        );

    \I__5721\ : InMux
    port map (
            O => \N__27189\,
            I => \N__27163\
        );

    \I__5720\ : CascadeMux
    port map (
            O => \N__27188\,
            I => \N__27159\
        );

    \I__5719\ : LocalMux
    port map (
            O => \N__27183\,
            I => \N__27156\
        );

    \I__5718\ : CascadeMux
    port map (
            O => \N__27182\,
            I => \N__27153\
        );

    \I__5717\ : LocalMux
    port map (
            O => \N__27179\,
            I => \N__27150\
        );

    \I__5716\ : LocalMux
    port map (
            O => \N__27174\,
            I => \N__27147\
        );

    \I__5715\ : LocalMux
    port map (
            O => \N__27171\,
            I => \N__27143\
        );

    \I__5714\ : LocalMux
    port map (
            O => \N__27168\,
            I => \N__27138\
        );

    \I__5713\ : LocalMux
    port map (
            O => \N__27163\,
            I => \N__27138\
        );

    \I__5712\ : InMux
    port map (
            O => \N__27162\,
            I => \N__27133\
        );

    \I__5711\ : InMux
    port map (
            O => \N__27159\,
            I => \N__27133\
        );

    \I__5710\ : Span4Mux_h
    port map (
            O => \N__27156\,
            I => \N__27130\
        );

    \I__5709\ : InMux
    port map (
            O => \N__27153\,
            I => \N__27127\
        );

    \I__5708\ : Span4Mux_v
    port map (
            O => \N__27150\,
            I => \N__27122\
        );

    \I__5707\ : Span4Mux_v
    port map (
            O => \N__27147\,
            I => \N__27122\
        );

    \I__5706\ : InMux
    port map (
            O => \N__27146\,
            I => \N__27119\
        );

    \I__5705\ : Odrv12
    port map (
            O => \N__27143\,
            I => \b2v_inst9.fsm_stateZ0Z_1\
        );

    \I__5704\ : Odrv4
    port map (
            O => \N__27138\,
            I => \b2v_inst9.fsm_stateZ0Z_1\
        );

    \I__5703\ : LocalMux
    port map (
            O => \N__27133\,
            I => \b2v_inst9.fsm_stateZ0Z_1\
        );

    \I__5702\ : Odrv4
    port map (
            O => \N__27130\,
            I => \b2v_inst9.fsm_stateZ0Z_1\
        );

    \I__5701\ : LocalMux
    port map (
            O => \N__27127\,
            I => \b2v_inst9.fsm_stateZ0Z_1\
        );

    \I__5700\ : Odrv4
    port map (
            O => \N__27122\,
            I => \b2v_inst9.fsm_stateZ0Z_1\
        );

    \I__5699\ : LocalMux
    port map (
            O => \N__27119\,
            I => \b2v_inst9.fsm_stateZ0Z_1\
        );

    \I__5698\ : CascadeMux
    port map (
            O => \N__27104\,
            I => \b2v_inst9.N_84_2_cascade_\
        );

    \I__5697\ : InMux
    port map (
            O => \N__27101\,
            I => \N__27098\
        );

    \I__5696\ : LocalMux
    port map (
            O => \N__27098\,
            I => \N__27094\
        );

    \I__5695\ : InMux
    port map (
            O => \N__27097\,
            I => \N__27091\
        );

    \I__5694\ : Odrv4
    port map (
            O => \N__27094\,
            I => \b2v_inst9.N_582\
        );

    \I__5693\ : LocalMux
    port map (
            O => \N__27091\,
            I => \b2v_inst9.N_582\
        );

    \I__5692\ : InMux
    port map (
            O => \N__27086\,
            I => \N__27083\
        );

    \I__5691\ : LocalMux
    port map (
            O => \N__27083\,
            I => \N__27080\
        );

    \I__5690\ : Span4Mux_v
    port map (
            O => \N__27080\,
            I => \N__27077\
        );

    \I__5689\ : Sp12to4
    port map (
            O => \N__27077\,
            I => \N__27074\
        );

    \I__5688\ : Span12Mux_h
    port map (
            O => \N__27074\,
            I => \N__27070\
        );

    \I__5687\ : InMux
    port map (
            O => \N__27073\,
            I => \N__27067\
        );

    \I__5686\ : Odrv12
    port map (
            O => \N__27070\,
            I => \SYNTHESIZED_WIRE_5_4\
        );

    \I__5685\ : LocalMux
    port map (
            O => \N__27067\,
            I => \SYNTHESIZED_WIRE_5_4\
        );

    \I__5684\ : CascadeMux
    port map (
            O => \N__27062\,
            I => \b2v_inst.un12_pix_count_intlto7_N_2LZ0Z1_cascade_\
        );

    \I__5683\ : InMux
    port map (
            O => \N__27059\,
            I => \N__27055\
        );

    \I__5682\ : InMux
    port map (
            O => \N__27058\,
            I => \N__27052\
        );

    \I__5681\ : LocalMux
    port map (
            O => \N__27055\,
            I => \N__27049\
        );

    \I__5680\ : LocalMux
    port map (
            O => \N__27052\,
            I => \N__27046\
        );

    \I__5679\ : Span4Mux_h
    port map (
            O => \N__27049\,
            I => \N__27043\
        );

    \I__5678\ : Span4Mux_v
    port map (
            O => \N__27046\,
            I => \N__27040\
        );

    \I__5677\ : Span4Mux_v
    port map (
            O => \N__27043\,
            I => \N__27035\
        );

    \I__5676\ : Span4Mux_h
    port map (
            O => \N__27040\,
            I => \N__27035\
        );

    \I__5675\ : Odrv4
    port map (
            O => \N__27035\,
            I => \b2v_inst.un13_pix_count_int_li_0\
        );

    \I__5674\ : CascadeMux
    port map (
            O => \N__27032\,
            I => \b2v_inst.un13_pix_count_int_li_0_cascade_\
        );

    \I__5673\ : InMux
    port map (
            O => \N__27029\,
            I => \N__27026\
        );

    \I__5672\ : LocalMux
    port map (
            O => \N__27026\,
            I => \N__27023\
        );

    \I__5671\ : Span4Mux_v
    port map (
            O => \N__27023\,
            I => \N__27019\
        );

    \I__5670\ : CascadeMux
    port map (
            O => \N__27022\,
            I => \N__27015\
        );

    \I__5669\ : Sp12to4
    port map (
            O => \N__27019\,
            I => \N__27012\
        );

    \I__5668\ : InMux
    port map (
            O => \N__27018\,
            I => \N__27009\
        );

    \I__5667\ : InMux
    port map (
            O => \N__27015\,
            I => \N__27006\
        );

    \I__5666\ : Odrv12
    port map (
            O => \N__27012\,
            I => \SYNTHESIZED_WIRE_10_1\
        );

    \I__5665\ : LocalMux
    port map (
            O => \N__27009\,
            I => \SYNTHESIZED_WIRE_10_1\
        );

    \I__5664\ : LocalMux
    port map (
            O => \N__27006\,
            I => \SYNTHESIZED_WIRE_10_1\
        );

    \I__5663\ : InMux
    port map (
            O => \N__26999\,
            I => \N__26995\
        );

    \I__5662\ : InMux
    port map (
            O => \N__26998\,
            I => \N__26992\
        );

    \I__5661\ : LocalMux
    port map (
            O => \N__26995\,
            I => \SYNTHESIZED_WIRE_5_1\
        );

    \I__5660\ : LocalMux
    port map (
            O => \N__26992\,
            I => \SYNTHESIZED_WIRE_5_1\
        );

    \I__5659\ : InMux
    port map (
            O => \N__26987\,
            I => \N__26983\
        );

    \I__5658\ : CascadeMux
    port map (
            O => \N__26986\,
            I => \N__26979\
        );

    \I__5657\ : LocalMux
    port map (
            O => \N__26983\,
            I => \N__26976\
        );

    \I__5656\ : InMux
    port map (
            O => \N__26982\,
            I => \N__26971\
        );

    \I__5655\ : InMux
    port map (
            O => \N__26979\,
            I => \N__26971\
        );

    \I__5654\ : Odrv12
    port map (
            O => \N__26976\,
            I => \SYNTHESIZED_WIRE_10_2\
        );

    \I__5653\ : LocalMux
    port map (
            O => \N__26971\,
            I => \SYNTHESIZED_WIRE_10_2\
        );

    \I__5652\ : InMux
    port map (
            O => \N__26966\,
            I => \N__26962\
        );

    \I__5651\ : InMux
    port map (
            O => \N__26965\,
            I => \N__26959\
        );

    \I__5650\ : LocalMux
    port map (
            O => \N__26962\,
            I => \SYNTHESIZED_WIRE_5_2\
        );

    \I__5649\ : LocalMux
    port map (
            O => \N__26959\,
            I => \SYNTHESIZED_WIRE_5_2\
        );

    \I__5648\ : CascadeMux
    port map (
            O => \N__26954\,
            I => \N__26951\
        );

    \I__5647\ : InMux
    port map (
            O => \N__26951\,
            I => \N__26947\
        );

    \I__5646\ : InMux
    port map (
            O => \N__26950\,
            I => \N__26944\
        );

    \I__5645\ : LocalMux
    port map (
            O => \N__26947\,
            I => \N__26941\
        );

    \I__5644\ : LocalMux
    port map (
            O => \N__26944\,
            I => \N__26938\
        );

    \I__5643\ : Span4Mux_h
    port map (
            O => \N__26941\,
            I => \N__26935\
        );

    \I__5642\ : Span4Mux_h
    port map (
            O => \N__26938\,
            I => \N__26929\
        );

    \I__5641\ : Span4Mux_h
    port map (
            O => \N__26935\,
            I => \N__26929\
        );

    \I__5640\ : InMux
    port map (
            O => \N__26934\,
            I => \N__26926\
        );

    \I__5639\ : Odrv4
    port map (
            O => \N__26929\,
            I => \b2v_inst.state_fastZ0Z_19\
        );

    \I__5638\ : LocalMux
    port map (
            O => \N__26926\,
            I => \b2v_inst.state_fastZ0Z_19\
        );

    \I__5637\ : InMux
    port map (
            O => \N__26921\,
            I => \N__26918\
        );

    \I__5636\ : LocalMux
    port map (
            O => \N__26918\,
            I => \b2v_inst9.fsm_state_srsts_1_0\
        );

    \I__5635\ : CascadeMux
    port map (
            O => \N__26915\,
            I => \N__26912\
        );

    \I__5634\ : InMux
    port map (
            O => \N__26912\,
            I => \N__26909\
        );

    \I__5633\ : LocalMux
    port map (
            O => \N__26909\,
            I => \b2v_inst9.N_522\
        );

    \I__5632\ : CascadeMux
    port map (
            O => \N__26906\,
            I => \b2v_inst9.N_522_cascade_\
        );

    \I__5631\ : InMux
    port map (
            O => \N__26903\,
            I => \N__26894\
        );

    \I__5630\ : InMux
    port map (
            O => \N__26902\,
            I => \N__26891\
        );

    \I__5629\ : InMux
    port map (
            O => \N__26901\,
            I => \N__26886\
        );

    \I__5628\ : InMux
    port map (
            O => \N__26900\,
            I => \N__26886\
        );

    \I__5627\ : InMux
    port map (
            O => \N__26899\,
            I => \N__26878\
        );

    \I__5626\ : InMux
    port map (
            O => \N__26898\,
            I => \N__26875\
        );

    \I__5625\ : InMux
    port map (
            O => \N__26897\,
            I => \N__26871\
        );

    \I__5624\ : LocalMux
    port map (
            O => \N__26894\,
            I => \N__26866\
        );

    \I__5623\ : LocalMux
    port map (
            O => \N__26891\,
            I => \N__26866\
        );

    \I__5622\ : LocalMux
    port map (
            O => \N__26886\,
            I => \N__26863\
        );

    \I__5621\ : InMux
    port map (
            O => \N__26885\,
            I => \N__26856\
        );

    \I__5620\ : InMux
    port map (
            O => \N__26884\,
            I => \N__26856\
        );

    \I__5619\ : InMux
    port map (
            O => \N__26883\,
            I => \N__26856\
        );

    \I__5618\ : InMux
    port map (
            O => \N__26882\,
            I => \N__26851\
        );

    \I__5617\ : InMux
    port map (
            O => \N__26881\,
            I => \N__26851\
        );

    \I__5616\ : LocalMux
    port map (
            O => \N__26878\,
            I => \N__26848\
        );

    \I__5615\ : LocalMux
    port map (
            O => \N__26875\,
            I => \N__26845\
        );

    \I__5614\ : InMux
    port map (
            O => \N__26874\,
            I => \N__26842\
        );

    \I__5613\ : LocalMux
    port map (
            O => \N__26871\,
            I => \N__26837\
        );

    \I__5612\ : Span4Mux_v
    port map (
            O => \N__26866\,
            I => \N__26837\
        );

    \I__5611\ : Span4Mux_v
    port map (
            O => \N__26863\,
            I => \N__26828\
        );

    \I__5610\ : LocalMux
    port map (
            O => \N__26856\,
            I => \N__26828\
        );

    \I__5609\ : LocalMux
    port map (
            O => \N__26851\,
            I => \N__26828\
        );

    \I__5608\ : Span4Mux_h
    port map (
            O => \N__26848\,
            I => \N__26828\
        );

    \I__5607\ : Odrv4
    port map (
            O => \N__26845\,
            I => \b2v_inst9.fsm_stateZ0Z_0\
        );

    \I__5606\ : LocalMux
    port map (
            O => \N__26842\,
            I => \b2v_inst9.fsm_stateZ0Z_0\
        );

    \I__5605\ : Odrv4
    port map (
            O => \N__26837\,
            I => \b2v_inst9.fsm_stateZ0Z_0\
        );

    \I__5604\ : Odrv4
    port map (
            O => \N__26828\,
            I => \b2v_inst9.fsm_stateZ0Z_0\
        );

    \I__5603\ : InMux
    port map (
            O => \N__26819\,
            I => \N__26816\
        );

    \I__5602\ : LocalMux
    port map (
            O => \N__26816\,
            I => \b2v_inst.N_268\
        );

    \I__5601\ : InMux
    port map (
            O => \N__26813\,
            I => \N__26810\
        );

    \I__5600\ : LocalMux
    port map (
            O => \N__26810\,
            I => \b2v_inst.un1_reg_anterior_iv_0_1_10\
        );

    \I__5599\ : InMux
    port map (
            O => \N__26807\,
            I => \N__26804\
        );

    \I__5598\ : LocalMux
    port map (
            O => \N__26804\,
            I => \N__26801\
        );

    \I__5597\ : Span4Mux_h
    port map (
            O => \N__26801\,
            I => \N__26797\
        );

    \I__5596\ : CascadeMux
    port map (
            O => \N__26800\,
            I => \N__26793\
        );

    \I__5595\ : Span4Mux_h
    port map (
            O => \N__26797\,
            I => \N__26790\
        );

    \I__5594\ : InMux
    port map (
            O => \N__26796\,
            I => \N__26785\
        );

    \I__5593\ : InMux
    port map (
            O => \N__26793\,
            I => \N__26785\
        );

    \I__5592\ : Odrv4
    port map (
            O => \N__26790\,
            I => \SYNTHESIZED_WIRE_10_3\
        );

    \I__5591\ : LocalMux
    port map (
            O => \N__26785\,
            I => \SYNTHESIZED_WIRE_10_3\
        );

    \I__5590\ : InMux
    port map (
            O => \N__26780\,
            I => \N__26777\
        );

    \I__5589\ : LocalMux
    port map (
            O => \N__26777\,
            I => \N__26774\
        );

    \I__5588\ : Span12Mux_h
    port map (
            O => \N__26774\,
            I => \N__26770\
        );

    \I__5587\ : InMux
    port map (
            O => \N__26773\,
            I => \N__26767\
        );

    \I__5586\ : Odrv12
    port map (
            O => \N__26770\,
            I => \SYNTHESIZED_WIRE_10_4\
        );

    \I__5585\ : LocalMux
    port map (
            O => \N__26767\,
            I => \SYNTHESIZED_WIRE_10_4\
        );

    \I__5584\ : InMux
    port map (
            O => \N__26762\,
            I => \N__26758\
        );

    \I__5583\ : CascadeMux
    port map (
            O => \N__26761\,
            I => \N__26755\
        );

    \I__5582\ : LocalMux
    port map (
            O => \N__26758\,
            I => \N__26752\
        );

    \I__5581\ : InMux
    port map (
            O => \N__26755\,
            I => \N__26749\
        );

    \I__5580\ : Odrv12
    port map (
            O => \N__26752\,
            I => \SYNTHESIZED_WIRE_10_6\
        );

    \I__5579\ : LocalMux
    port map (
            O => \N__26749\,
            I => \SYNTHESIZED_WIRE_10_6\
        );

    \I__5578\ : InMux
    port map (
            O => \N__26744\,
            I => \N__26741\
        );

    \I__5577\ : LocalMux
    port map (
            O => \N__26741\,
            I => \N__26738\
        );

    \I__5576\ : Span4Mux_h
    port map (
            O => \N__26738\,
            I => \N__26734\
        );

    \I__5575\ : CascadeMux
    port map (
            O => \N__26737\,
            I => \N__26731\
        );

    \I__5574\ : Span4Mux_h
    port map (
            O => \N__26734\,
            I => \N__26728\
        );

    \I__5573\ : InMux
    port map (
            O => \N__26731\,
            I => \N__26725\
        );

    \I__5572\ : Odrv4
    port map (
            O => \N__26728\,
            I => \SYNTHESIZED_WIRE_10_7\
        );

    \I__5571\ : LocalMux
    port map (
            O => \N__26725\,
            I => \SYNTHESIZED_WIRE_10_7\
        );

    \I__5570\ : InMux
    port map (
            O => \N__26720\,
            I => \N__26717\
        );

    \I__5569\ : LocalMux
    port map (
            O => \N__26717\,
            I => \N__26713\
        );

    \I__5568\ : CascadeMux
    port map (
            O => \N__26716\,
            I => \N__26709\
        );

    \I__5567\ : Sp12to4
    port map (
            O => \N__26713\,
            I => \N__26706\
        );

    \I__5566\ : InMux
    port map (
            O => \N__26712\,
            I => \N__26703\
        );

    \I__5565\ : InMux
    port map (
            O => \N__26709\,
            I => \N__26700\
        );

    \I__5564\ : Span12Mux_v
    port map (
            O => \N__26706\,
            I => \N__26697\
        );

    \I__5563\ : LocalMux
    port map (
            O => \N__26703\,
            I => \SYNTHESIZED_WIRE_10_0\
        );

    \I__5562\ : LocalMux
    port map (
            O => \N__26700\,
            I => \SYNTHESIZED_WIRE_10_0\
        );

    \I__5561\ : Odrv12
    port map (
            O => \N__26697\,
            I => \SYNTHESIZED_WIRE_10_0\
        );

    \I__5560\ : InMux
    port map (
            O => \N__26690\,
            I => \N__26686\
        );

    \I__5559\ : InMux
    port map (
            O => \N__26689\,
            I => \N__26683\
        );

    \I__5558\ : LocalMux
    port map (
            O => \N__26686\,
            I => \SYNTHESIZED_WIRE_5_0\
        );

    \I__5557\ : LocalMux
    port map (
            O => \N__26683\,
            I => \SYNTHESIZED_WIRE_5_0\
        );

    \I__5556\ : InMux
    port map (
            O => \N__26678\,
            I => \N__26675\
        );

    \I__5555\ : LocalMux
    port map (
            O => \N__26675\,
            I => \N__26671\
        );

    \I__5554\ : InMux
    port map (
            O => \N__26674\,
            I => \N__26668\
        );

    \I__5553\ : Span4Mux_h
    port map (
            O => \N__26671\,
            I => \N__26665\
        );

    \I__5552\ : LocalMux
    port map (
            O => \N__26668\,
            I => \b2v_inst.eventosZ0Z_6\
        );

    \I__5551\ : Odrv4
    port map (
            O => \N__26665\,
            I => \b2v_inst.eventosZ0Z_6\
        );

    \I__5550\ : CascadeMux
    port map (
            O => \N__26660\,
            I => \b2v_inst.un1_reg_anterior_iv_0_0_6_cascade_\
        );

    \I__5549\ : InMux
    port map (
            O => \N__26657\,
            I => \N__26654\
        );

    \I__5548\ : LocalMux
    port map (
            O => \N__26654\,
            I => \b2v_inst.N_272\
        );

    \I__5547\ : CEMux
    port map (
            O => \N__26651\,
            I => \N__26648\
        );

    \I__5546\ : LocalMux
    port map (
            O => \N__26648\,
            I => \N__26644\
        );

    \I__5545\ : CEMux
    port map (
            O => \N__26647\,
            I => \N__26641\
        );

    \I__5544\ : Span4Mux_h
    port map (
            O => \N__26644\,
            I => \N__26638\
        );

    \I__5543\ : LocalMux
    port map (
            O => \N__26641\,
            I => \N__26635\
        );

    \I__5542\ : Odrv4
    port map (
            O => \N__26638\,
            I => \b2v_inst.data_a_escribir_1_sqmuxa\
        );

    \I__5541\ : Odrv12
    port map (
            O => \N__26635\,
            I => \b2v_inst.data_a_escribir_1_sqmuxa\
        );

    \I__5540\ : InMux
    port map (
            O => \N__26630\,
            I => \N__26627\
        );

    \I__5539\ : LocalMux
    port map (
            O => \N__26627\,
            I => \N__26624\
        );

    \I__5538\ : Span4Mux_h
    port map (
            O => \N__26624\,
            I => \N__26621\
        );

    \I__5537\ : Odrv4
    port map (
            O => \N__26621\,
            I => \b2v_inst.data_a_escribir11_1_and\
        );

    \I__5536\ : InMux
    port map (
            O => \N__26618\,
            I => \N__26614\
        );

    \I__5535\ : InMux
    port map (
            O => \N__26617\,
            I => \N__26611\
        );

    \I__5534\ : LocalMux
    port map (
            O => \N__26614\,
            I => \N__26608\
        );

    \I__5533\ : LocalMux
    port map (
            O => \N__26611\,
            I => \b2v_inst.eventosZ0Z_4\
        );

    \I__5532\ : Odrv4
    port map (
            O => \N__26608\,
            I => \b2v_inst.eventosZ0Z_4\
        );

    \I__5531\ : CascadeMux
    port map (
            O => \N__26603\,
            I => \b2v_inst.un1_reg_anterior_iv_0_0_4_cascade_\
        );

    \I__5530\ : CascadeMux
    port map (
            O => \N__26600\,
            I => \b2v_inst.un1_reg_anterior_iv_0_1_4_cascade_\
        );

    \I__5529\ : InMux
    port map (
            O => \N__26597\,
            I => \N__26594\
        );

    \I__5528\ : LocalMux
    port map (
            O => \N__26594\,
            I => \b2v_inst.N_274\
        );

    \I__5527\ : InMux
    port map (
            O => \N__26591\,
            I => \N__26587\
        );

    \I__5526\ : InMux
    port map (
            O => \N__26590\,
            I => \N__26584\
        );

    \I__5525\ : LocalMux
    port map (
            O => \N__26587\,
            I => \b2v_inst.eventosZ0Z_0\
        );

    \I__5524\ : LocalMux
    port map (
            O => \N__26584\,
            I => \b2v_inst.eventosZ0Z_0\
        );

    \I__5523\ : CascadeMux
    port map (
            O => \N__26579\,
            I => \b2v_inst.data_a_escribir_RNO_2Z0Z_0_cascade_\
        );

    \I__5522\ : CascadeMux
    port map (
            O => \N__26576\,
            I => \b2v_inst.un1_reg_anterior_0_i_1_0_cascade_\
        );

    \I__5521\ : InMux
    port map (
            O => \N__26573\,
            I => \N__26570\
        );

    \I__5520\ : LocalMux
    port map (
            O => \N__26570\,
            I => \N__26566\
        );

    \I__5519\ : InMux
    port map (
            O => \N__26569\,
            I => \N__26563\
        );

    \I__5518\ : Odrv4
    port map (
            O => \N__26566\,
            I => \b2v_inst.eventosZ0Z_1\
        );

    \I__5517\ : LocalMux
    port map (
            O => \N__26563\,
            I => \b2v_inst.eventosZ0Z_1\
        );

    \I__5516\ : CascadeMux
    port map (
            O => \N__26558\,
            I => \b2v_inst.data_a_escribir_RNO_2Z0Z_1_cascade_\
        );

    \I__5515\ : CascadeMux
    port map (
            O => \N__26555\,
            I => \b2v_inst.un1_reg_anterior_0_i_1_1_cascade_\
        );

    \I__5514\ : InMux
    port map (
            O => \N__26552\,
            I => \N__26548\
        );

    \I__5513\ : InMux
    port map (
            O => \N__26551\,
            I => \N__26545\
        );

    \I__5512\ : LocalMux
    port map (
            O => \N__26548\,
            I => \b2v_inst.eventosZ0Z_10\
        );

    \I__5511\ : LocalMux
    port map (
            O => \N__26545\,
            I => \b2v_inst.eventosZ0Z_10\
        );

    \I__5510\ : InMux
    port map (
            O => \N__26540\,
            I => \N__26537\
        );

    \I__5509\ : LocalMux
    port map (
            O => \N__26537\,
            I => \b2v_inst.N_269\
        );

    \I__5508\ : CascadeMux
    port map (
            O => \N__26534\,
            I => \b2v_inst.un1_reg_anterior_iv_0_0_10_cascade_\
        );

    \I__5507\ : InMux
    port map (
            O => \N__26531\,
            I => \b2v_inst.un2_valor_max1\
        );

    \I__5506\ : InMux
    port map (
            O => \N__26528\,
            I => \N__26503\
        );

    \I__5505\ : InMux
    port map (
            O => \N__26527\,
            I => \N__26503\
        );

    \I__5504\ : InMux
    port map (
            O => \N__26526\,
            I => \N__26503\
        );

    \I__5503\ : InMux
    port map (
            O => \N__26525\,
            I => \N__26503\
        );

    \I__5502\ : InMux
    port map (
            O => \N__26524\,
            I => \N__26503\
        );

    \I__5501\ : InMux
    port map (
            O => \N__26523\,
            I => \N__26503\
        );

    \I__5500\ : InMux
    port map (
            O => \N__26522\,
            I => \N__26503\
        );

    \I__5499\ : InMux
    port map (
            O => \N__26521\,
            I => \N__26500\
        );

    \I__5498\ : InMux
    port map (
            O => \N__26520\,
            I => \N__26493\
        );

    \I__5497\ : InMux
    port map (
            O => \N__26519\,
            I => \N__26493\
        );

    \I__5496\ : InMux
    port map (
            O => \N__26518\,
            I => \N__26493\
        );

    \I__5495\ : LocalMux
    port map (
            O => \N__26503\,
            I => \N__26490\
        );

    \I__5494\ : LocalMux
    port map (
            O => \N__26500\,
            I => \N__26485\
        );

    \I__5493\ : LocalMux
    port map (
            O => \N__26493\,
            I => \N__26485\
        );

    \I__5492\ : Span4Mux_v
    port map (
            O => \N__26490\,
            I => \N__26482\
        );

    \I__5491\ : Span4Mux_h
    port map (
            O => \N__26485\,
            I => \N__26479\
        );

    \I__5490\ : Sp12to4
    port map (
            O => \N__26482\,
            I => \N__26476\
        );

    \I__5489\ : Span4Mux_h
    port map (
            O => \N__26479\,
            I => \N__26473\
        );

    \I__5488\ : Span12Mux_h
    port map (
            O => \N__26476\,
            I => \N__26470\
        );

    \I__5487\ : Span4Mux_h
    port map (
            O => \N__26473\,
            I => \N__26467\
        );

    \I__5486\ : Odrv12
    port map (
            O => \N__26470\,
            I => \b2v_inst.ignorar_anchoZ0Z_1\
        );

    \I__5485\ : Odrv4
    port map (
            O => \N__26467\,
            I => \b2v_inst.ignorar_anchoZ0Z_1\
        );

    \I__5484\ : CEMux
    port map (
            O => \N__26462\,
            I => \N__26459\
        );

    \I__5483\ : LocalMux
    port map (
            O => \N__26459\,
            I => \N__26455\
        );

    \I__5482\ : CEMux
    port map (
            O => \N__26458\,
            I => \N__26452\
        );

    \I__5481\ : Span4Mux_h
    port map (
            O => \N__26455\,
            I => \N__26446\
        );

    \I__5480\ : LocalMux
    port map (
            O => \N__26452\,
            I => \N__26443\
        );

    \I__5479\ : InMux
    port map (
            O => \N__26451\,
            I => \N__26436\
        );

    \I__5478\ : InMux
    port map (
            O => \N__26450\,
            I => \N__26436\
        );

    \I__5477\ : InMux
    port map (
            O => \N__26449\,
            I => \N__26433\
        );

    \I__5476\ : Span4Mux_v
    port map (
            O => \N__26446\,
            I => \N__26430\
        );

    \I__5475\ : Span4Mux_h
    port map (
            O => \N__26443\,
            I => \N__26427\
        );

    \I__5474\ : InMux
    port map (
            O => \N__26442\,
            I => \N__26422\
        );

    \I__5473\ : InMux
    port map (
            O => \N__26441\,
            I => \N__26422\
        );

    \I__5472\ : LocalMux
    port map (
            O => \N__26436\,
            I => \N__26417\
        );

    \I__5471\ : LocalMux
    port map (
            O => \N__26433\,
            I => \N__26417\
        );

    \I__5470\ : Odrv4
    port map (
            O => \N__26430\,
            I => \b2v_inst.stateZ0Z_25\
        );

    \I__5469\ : Odrv4
    port map (
            O => \N__26427\,
            I => \b2v_inst.stateZ0Z_25\
        );

    \I__5468\ : LocalMux
    port map (
            O => \N__26422\,
            I => \b2v_inst.stateZ0Z_25\
        );

    \I__5467\ : Odrv4
    port map (
            O => \N__26417\,
            I => \b2v_inst.stateZ0Z_25\
        );

    \I__5466\ : InMux
    port map (
            O => \N__26408\,
            I => \N__26405\
        );

    \I__5465\ : LocalMux
    port map (
            O => \N__26405\,
            I => \N__26402\
        );

    \I__5464\ : Odrv4
    port map (
            O => \N__26402\,
            I => \b2v_inst.data_a_escribir11_0_and\
        );

    \I__5463\ : CascadeMux
    port map (
            O => \N__26399\,
            I => \N__26396\
        );

    \I__5462\ : InMux
    port map (
            O => \N__26396\,
            I => \N__26393\
        );

    \I__5461\ : LocalMux
    port map (
            O => \N__26393\,
            I => \b2v_inst.reg_ancho_1_i_3\
        );

    \I__5460\ : CascadeMux
    port map (
            O => \N__26390\,
            I => \N__26387\
        );

    \I__5459\ : InMux
    port map (
            O => \N__26387\,
            I => \N__26384\
        );

    \I__5458\ : LocalMux
    port map (
            O => \N__26384\,
            I => \b2v_inst.reg_ancho_1_i_4\
        );

    \I__5457\ : CascadeMux
    port map (
            O => \N__26381\,
            I => \N__26378\
        );

    \I__5456\ : InMux
    port map (
            O => \N__26378\,
            I => \N__26375\
        );

    \I__5455\ : LocalMux
    port map (
            O => \N__26375\,
            I => \b2v_inst.reg_ancho_1_i_5\
        );

    \I__5454\ : CascadeMux
    port map (
            O => \N__26372\,
            I => \N__26369\
        );

    \I__5453\ : InMux
    port map (
            O => \N__26369\,
            I => \N__26366\
        );

    \I__5452\ : LocalMux
    port map (
            O => \N__26366\,
            I => \b2v_inst.reg_ancho_1_i_6\
        );

    \I__5451\ : CascadeMux
    port map (
            O => \N__26363\,
            I => \N__26360\
        );

    \I__5450\ : InMux
    port map (
            O => \N__26360\,
            I => \N__26357\
        );

    \I__5449\ : LocalMux
    port map (
            O => \N__26357\,
            I => \b2v_inst.reg_ancho_1_i_7\
        );

    \I__5448\ : CascadeMux
    port map (
            O => \N__26354\,
            I => \N__26351\
        );

    \I__5447\ : InMux
    port map (
            O => \N__26351\,
            I => \N__26348\
        );

    \I__5446\ : LocalMux
    port map (
            O => \N__26348\,
            I => \b2v_inst.reg_ancho_1_i_8\
        );

    \I__5445\ : CascadeMux
    port map (
            O => \N__26345\,
            I => \N__26342\
        );

    \I__5444\ : InMux
    port map (
            O => \N__26342\,
            I => \N__26339\
        );

    \I__5443\ : LocalMux
    port map (
            O => \N__26339\,
            I => \b2v_inst.reg_ancho_1_i_9\
        );

    \I__5442\ : CascadeMux
    port map (
            O => \N__26336\,
            I => \N__26333\
        );

    \I__5441\ : InMux
    port map (
            O => \N__26333\,
            I => \N__26330\
        );

    \I__5440\ : LocalMux
    port map (
            O => \N__26330\,
            I => \b2v_inst.reg_ancho_1_i_10\
        );

    \I__5439\ : CascadeMux
    port map (
            O => \N__26327\,
            I => \N__26324\
        );

    \I__5438\ : InMux
    port map (
            O => \N__26324\,
            I => \N__26321\
        );

    \I__5437\ : LocalMux
    port map (
            O => \N__26321\,
            I => \b2v_inst.reg_ancho_1_i_0\
        );

    \I__5436\ : CascadeMux
    port map (
            O => \N__26318\,
            I => \N__26315\
        );

    \I__5435\ : InMux
    port map (
            O => \N__26315\,
            I => \N__26312\
        );

    \I__5434\ : LocalMux
    port map (
            O => \N__26312\,
            I => \b2v_inst.reg_ancho_1_i_1\
        );

    \I__5433\ : CascadeMux
    port map (
            O => \N__26309\,
            I => \N__26306\
        );

    \I__5432\ : InMux
    port map (
            O => \N__26306\,
            I => \N__26303\
        );

    \I__5431\ : LocalMux
    port map (
            O => \N__26303\,
            I => \b2v_inst.reg_ancho_1_i_2\
        );

    \I__5430\ : InMux
    port map (
            O => \N__26300\,
            I => \N__26297\
        );

    \I__5429\ : LocalMux
    port map (
            O => \N__26297\,
            I => \b2v_inst.pix_data_regZ0Z_2\
        );

    \I__5428\ : CascadeMux
    port map (
            O => \N__26294\,
            I => \N__26291\
        );

    \I__5427\ : InMux
    port map (
            O => \N__26291\,
            I => \N__26288\
        );

    \I__5426\ : LocalMux
    port map (
            O => \N__26288\,
            I => \b2v_inst.pix_data_regZ0Z_5\
        );

    \I__5425\ : InMux
    port map (
            O => \N__26285\,
            I => \N__26282\
        );

    \I__5424\ : LocalMux
    port map (
            O => \N__26282\,
            I => \b2v_inst.pix_data_regZ0Z_6\
        );

    \I__5423\ : InMux
    port map (
            O => \N__26279\,
            I => \N__26276\
        );

    \I__5422\ : LocalMux
    port map (
            O => \N__26276\,
            I => \b2v_inst.pix_data_regZ0Z_7\
        );

    \I__5421\ : InMux
    port map (
            O => \N__26273\,
            I => \N__26270\
        );

    \I__5420\ : LocalMux
    port map (
            O => \N__26270\,
            I => \N__26267\
        );

    \I__5419\ : Span4Mux_v
    port map (
            O => \N__26267\,
            I => \N__26264\
        );

    \I__5418\ : Odrv4
    port map (
            O => \N__26264\,
            I => \b2v_inst9.N_583\
        );

    \I__5417\ : IoInMux
    port map (
            O => \N__26261\,
            I => \N__26257\
        );

    \I__5416\ : InMux
    port map (
            O => \N__26260\,
            I => \N__26254\
        );

    \I__5415\ : LocalMux
    port map (
            O => \N__26257\,
            I => \N__26251\
        );

    \I__5414\ : LocalMux
    port map (
            O => \N__26254\,
            I => \N__26248\
        );

    \I__5413\ : IoSpan4Mux
    port map (
            O => \N__26251\,
            I => \N__26245\
        );

    \I__5412\ : Span4Mux_h
    port map (
            O => \N__26248\,
            I => \N__26242\
        );

    \I__5411\ : Span4Mux_s3_h
    port map (
            O => \N__26245\,
            I => \N__26239\
        );

    \I__5410\ : Span4Mux_h
    port map (
            O => \N__26242\,
            I => \N__26236\
        );

    \I__5409\ : Span4Mux_h
    port map (
            O => \N__26239\,
            I => \N__26233\
        );

    \I__5408\ : Span4Mux_h
    port map (
            O => \N__26236\,
            I => \N__26230\
        );

    \I__5407\ : Odrv4
    port map (
            O => \N__26233\,
            I => leds_c_9
        );

    \I__5406\ : Odrv4
    port map (
            O => \N__26230\,
            I => leds_c_9
        );

    \I__5405\ : InMux
    port map (
            O => \N__26225\,
            I => \N__26222\
        );

    \I__5404\ : LocalMux
    port map (
            O => \N__26222\,
            I => \N__26218\
        );

    \I__5403\ : InMux
    port map (
            O => \N__26221\,
            I => \N__26215\
        );

    \I__5402\ : Span4Mux_h
    port map (
            O => \N__26218\,
            I => \N__26210\
        );

    \I__5401\ : LocalMux
    port map (
            O => \N__26215\,
            I => \N__26210\
        );

    \I__5400\ : Odrv4
    port map (
            O => \N__26210\,
            I => b2v_inst_energia_temp_9
        );

    \I__5399\ : CEMux
    port map (
            O => \N__26207\,
            I => \N__26202\
        );

    \I__5398\ : CEMux
    port map (
            O => \N__26206\,
            I => \N__26199\
        );

    \I__5397\ : CEMux
    port map (
            O => \N__26205\,
            I => \N__26194\
        );

    \I__5396\ : LocalMux
    port map (
            O => \N__26202\,
            I => \N__26191\
        );

    \I__5395\ : LocalMux
    port map (
            O => \N__26199\,
            I => \N__26187\
        );

    \I__5394\ : CEMux
    port map (
            O => \N__26198\,
            I => \N__26184\
        );

    \I__5393\ : CEMux
    port map (
            O => \N__26197\,
            I => \N__26181\
        );

    \I__5392\ : LocalMux
    port map (
            O => \N__26194\,
            I => \N__26177\
        );

    \I__5391\ : Span4Mux_v
    port map (
            O => \N__26191\,
            I => \N__26174\
        );

    \I__5390\ : CEMux
    port map (
            O => \N__26190\,
            I => \N__26171\
        );

    \I__5389\ : Span4Mux_v
    port map (
            O => \N__26187\,
            I => \N__26168\
        );

    \I__5388\ : LocalMux
    port map (
            O => \N__26184\,
            I => \N__26163\
        );

    \I__5387\ : LocalMux
    port map (
            O => \N__26181\,
            I => \N__26163\
        );

    \I__5386\ : CEMux
    port map (
            O => \N__26180\,
            I => \N__26160\
        );

    \I__5385\ : Span4Mux_v
    port map (
            O => \N__26177\,
            I => \N__26153\
        );

    \I__5384\ : Span4Mux_h
    port map (
            O => \N__26174\,
            I => \N__26153\
        );

    \I__5383\ : LocalMux
    port map (
            O => \N__26171\,
            I => \N__26153\
        );

    \I__5382\ : Span4Mux_h
    port map (
            O => \N__26168\,
            I => \N__26150\
        );

    \I__5381\ : Span4Mux_h
    port map (
            O => \N__26163\,
            I => \N__26145\
        );

    \I__5380\ : LocalMux
    port map (
            O => \N__26160\,
            I => \N__26145\
        );

    \I__5379\ : Span4Mux_v
    port map (
            O => \N__26153\,
            I => \N__26141\
        );

    \I__5378\ : Span4Mux_v
    port map (
            O => \N__26150\,
            I => \N__26136\
        );

    \I__5377\ : Span4Mux_v
    port map (
            O => \N__26145\,
            I => \N__26136\
        );

    \I__5376\ : CEMux
    port map (
            O => \N__26144\,
            I => \N__26133\
        );

    \I__5375\ : Span4Mux_v
    port map (
            O => \N__26141\,
            I => \N__26130\
        );

    \I__5374\ : Span4Mux_v
    port map (
            O => \N__26136\,
            I => \N__26127\
        );

    \I__5373\ : LocalMux
    port map (
            O => \N__26133\,
            I => \N__26124\
        );

    \I__5372\ : Span4Mux_h
    port map (
            O => \N__26130\,
            I => \N__26121\
        );

    \I__5371\ : Span4Mux_h
    port map (
            O => \N__26127\,
            I => \N__26116\
        );

    \I__5370\ : Span4Mux_v
    port map (
            O => \N__26124\,
            I => \N__26116\
        );

    \I__5369\ : Odrv4
    port map (
            O => \N__26121\,
            I => \b2v_inst.N_577_i\
        );

    \I__5368\ : Odrv4
    port map (
            O => \N__26116\,
            I => \b2v_inst.N_577_i\
        );

    \I__5367\ : InMux
    port map (
            O => \N__26111\,
            I => \N__26108\
        );

    \I__5366\ : LocalMux
    port map (
            O => \N__26108\,
            I => \N__26105\
        );

    \I__5365\ : Span4Mux_v
    port map (
            O => \N__26105\,
            I => \N__26102\
        );

    \I__5364\ : Odrv4
    port map (
            O => \N__26102\,
            I => \b2v_inst9.data_to_sendZ0Z_0\
        );

    \I__5363\ : IoInMux
    port map (
            O => \N__26099\,
            I => \N__26096\
        );

    \I__5362\ : LocalMux
    port map (
            O => \N__26096\,
            I => \N__26093\
        );

    \I__5361\ : IoSpan4Mux
    port map (
            O => \N__26093\,
            I => \N__26090\
        );

    \I__5360\ : Span4Mux_s2_v
    port map (
            O => \N__26090\,
            I => \N__26087\
        );

    \I__5359\ : Sp12to4
    port map (
            O => \N__26087\,
            I => \N__26084\
        );

    \I__5358\ : Span12Mux_s10_v
    port map (
            O => \N__26084\,
            I => \N__26081\
        );

    \I__5357\ : Span12Mux_h
    port map (
            O => \N__26081\,
            I => \N__26078\
        );

    \I__5356\ : Odrv12
    port map (
            O => \N__26078\,
            I => uart_tx_o_c
        );

    \I__5355\ : InMux
    port map (
            O => \N__26075\,
            I => \N__26071\
        );

    \I__5354\ : InMux
    port map (
            O => \N__26074\,
            I => \N__26068\
        );

    \I__5353\ : LocalMux
    port map (
            O => \N__26071\,
            I => \N__26062\
        );

    \I__5352\ : LocalMux
    port map (
            O => \N__26068\,
            I => \N__26062\
        );

    \I__5351\ : InMux
    port map (
            O => \N__26067\,
            I => \N__26057\
        );

    \I__5350\ : Span4Mux_h
    port map (
            O => \N__26062\,
            I => \N__26054\
        );

    \I__5349\ : InMux
    port map (
            O => \N__26061\,
            I => \N__26051\
        );

    \I__5348\ : InMux
    port map (
            O => \N__26060\,
            I => \N__26048\
        );

    \I__5347\ : LocalMux
    port map (
            O => \N__26057\,
            I => \N__26045\
        );

    \I__5346\ : Span4Mux_h
    port map (
            O => \N__26054\,
            I => \N__26042\
        );

    \I__5345\ : LocalMux
    port map (
            O => \N__26051\,
            I => b2v_inst_state_2
        );

    \I__5344\ : LocalMux
    port map (
            O => \N__26048\,
            I => b2v_inst_state_2
        );

    \I__5343\ : Odrv4
    port map (
            O => \N__26045\,
            I => b2v_inst_state_2
        );

    \I__5342\ : Odrv4
    port map (
            O => \N__26042\,
            I => b2v_inst_state_2
        );

    \I__5341\ : CascadeMux
    port map (
            O => \N__26033\,
            I => \N__26028\
        );

    \I__5340\ : InMux
    port map (
            O => \N__26032\,
            I => \N__26025\
        );

    \I__5339\ : CascadeMux
    port map (
            O => \N__26031\,
            I => \N__26022\
        );

    \I__5338\ : InMux
    port map (
            O => \N__26028\,
            I => \N__26018\
        );

    \I__5337\ : LocalMux
    port map (
            O => \N__26025\,
            I => \N__26015\
        );

    \I__5336\ : InMux
    port map (
            O => \N__26022\,
            I => \N__26011\
        );

    \I__5335\ : CascadeMux
    port map (
            O => \N__26021\,
            I => \N__26008\
        );

    \I__5334\ : LocalMux
    port map (
            O => \N__26018\,
            I => \N__26005\
        );

    \I__5333\ : Span4Mux_v
    port map (
            O => \N__26015\,
            I => \N__26001\
        );

    \I__5332\ : InMux
    port map (
            O => \N__26014\,
            I => \N__25998\
        );

    \I__5331\ : LocalMux
    port map (
            O => \N__26011\,
            I => \N__25995\
        );

    \I__5330\ : InMux
    port map (
            O => \N__26008\,
            I => \N__25992\
        );

    \I__5329\ : Span4Mux_v
    port map (
            O => \N__26005\,
            I => \N__25989\
        );

    \I__5328\ : InMux
    port map (
            O => \N__26004\,
            I => \N__25986\
        );

    \I__5327\ : Span4Mux_v
    port map (
            O => \N__26001\,
            I => \N__25981\
        );

    \I__5326\ : LocalMux
    port map (
            O => \N__25998\,
            I => \N__25981\
        );

    \I__5325\ : Span4Mux_v
    port map (
            O => \N__25995\,
            I => \N__25978\
        );

    \I__5324\ : LocalMux
    port map (
            O => \N__25992\,
            I => \N__25975\
        );

    \I__5323\ : Sp12to4
    port map (
            O => \N__25989\,
            I => \N__25970\
        );

    \I__5322\ : LocalMux
    port map (
            O => \N__25986\,
            I => \N__25970\
        );

    \I__5321\ : Span4Mux_h
    port map (
            O => \N__25981\,
            I => \N__25963\
        );

    \I__5320\ : Span4Mux_v
    port map (
            O => \N__25978\,
            I => \N__25963\
        );

    \I__5319\ : Span4Mux_h
    port map (
            O => \N__25975\,
            I => \N__25963\
        );

    \I__5318\ : Odrv12
    port map (
            O => \N__25970\,
            I => \b2v_inst.stateZ0Z_11\
        );

    \I__5317\ : Odrv4
    port map (
            O => \N__25963\,
            I => \b2v_inst.stateZ0Z_11\
        );

    \I__5316\ : InMux
    port map (
            O => \N__25958\,
            I => \N__25942\
        );

    \I__5315\ : InMux
    port map (
            O => \N__25957\,
            I => \N__25942\
        );

    \I__5314\ : InMux
    port map (
            O => \N__25956\,
            I => \N__25942\
        );

    \I__5313\ : InMux
    port map (
            O => \N__25955\,
            I => \N__25942\
        );

    \I__5312\ : InMux
    port map (
            O => \N__25954\,
            I => \N__25939\
        );

    \I__5311\ : InMux
    port map (
            O => \N__25953\,
            I => \N__25936\
        );

    \I__5310\ : InMux
    port map (
            O => \N__25952\,
            I => \N__25930\
        );

    \I__5309\ : CascadeMux
    port map (
            O => \N__25951\,
            I => \N__25927\
        );

    \I__5308\ : LocalMux
    port map (
            O => \N__25942\,
            I => \N__25922\
        );

    \I__5307\ : LocalMux
    port map (
            O => \N__25939\,
            I => \N__25922\
        );

    \I__5306\ : LocalMux
    port map (
            O => \N__25936\,
            I => \N__25919\
        );

    \I__5305\ : CascadeMux
    port map (
            O => \N__25935\,
            I => \N__25916\
        );

    \I__5304\ : CascadeMux
    port map (
            O => \N__25934\,
            I => \N__25913\
        );

    \I__5303\ : CascadeMux
    port map (
            O => \N__25933\,
            I => \N__25906\
        );

    \I__5302\ : LocalMux
    port map (
            O => \N__25930\,
            I => \N__25903\
        );

    \I__5301\ : InMux
    port map (
            O => \N__25927\,
            I => \N__25900\
        );

    \I__5300\ : Span4Mux_h
    port map (
            O => \N__25922\,
            I => \N__25896\
        );

    \I__5299\ : Span4Mux_v
    port map (
            O => \N__25919\,
            I => \N__25893\
        );

    \I__5298\ : InMux
    port map (
            O => \N__25916\,
            I => \N__25890\
        );

    \I__5297\ : InMux
    port map (
            O => \N__25913\,
            I => \N__25887\
        );

    \I__5296\ : InMux
    port map (
            O => \N__25912\,
            I => \N__25876\
        );

    \I__5295\ : InMux
    port map (
            O => \N__25911\,
            I => \N__25876\
        );

    \I__5294\ : InMux
    port map (
            O => \N__25910\,
            I => \N__25876\
        );

    \I__5293\ : InMux
    port map (
            O => \N__25909\,
            I => \N__25876\
        );

    \I__5292\ : InMux
    port map (
            O => \N__25906\,
            I => \N__25876\
        );

    \I__5291\ : Span4Mux_h
    port map (
            O => \N__25903\,
            I => \N__25873\
        );

    \I__5290\ : LocalMux
    port map (
            O => \N__25900\,
            I => \N__25870\
        );

    \I__5289\ : CascadeMux
    port map (
            O => \N__25899\,
            I => \N__25867\
        );

    \I__5288\ : Span4Mux_v
    port map (
            O => \N__25896\,
            I => \N__25864\
        );

    \I__5287\ : Span4Mux_v
    port map (
            O => \N__25893\,
            I => \N__25861\
        );

    \I__5286\ : LocalMux
    port map (
            O => \N__25890\,
            I => \N__25858\
        );

    \I__5285\ : LocalMux
    port map (
            O => \N__25887\,
            I => \N__25853\
        );

    \I__5284\ : LocalMux
    port map (
            O => \N__25876\,
            I => \N__25853\
        );

    \I__5283\ : Span4Mux_v
    port map (
            O => \N__25873\,
            I => \N__25850\
        );

    \I__5282\ : Span12Mux_v
    port map (
            O => \N__25870\,
            I => \N__25847\
        );

    \I__5281\ : InMux
    port map (
            O => \N__25867\,
            I => \N__25844\
        );

    \I__5280\ : Odrv4
    port map (
            O => \N__25864\,
            I => \b2v_inst.stateZ0Z_32\
        );

    \I__5279\ : Odrv4
    port map (
            O => \N__25861\,
            I => \b2v_inst.stateZ0Z_32\
        );

    \I__5278\ : Odrv4
    port map (
            O => \N__25858\,
            I => \b2v_inst.stateZ0Z_32\
        );

    \I__5277\ : Odrv4
    port map (
            O => \N__25853\,
            I => \b2v_inst.stateZ0Z_32\
        );

    \I__5276\ : Odrv4
    port map (
            O => \N__25850\,
            I => \b2v_inst.stateZ0Z_32\
        );

    \I__5275\ : Odrv12
    port map (
            O => \N__25847\,
            I => \b2v_inst.stateZ0Z_32\
        );

    \I__5274\ : LocalMux
    port map (
            O => \N__25844\,
            I => \b2v_inst.stateZ0Z_32\
        );

    \I__5273\ : InMux
    port map (
            O => \N__25829\,
            I => \N__25824\
        );

    \I__5272\ : InMux
    port map (
            O => \N__25828\,
            I => \N__25821\
        );

    \I__5271\ : InMux
    port map (
            O => \N__25827\,
            I => \N__25818\
        );

    \I__5270\ : LocalMux
    port map (
            O => \N__25824\,
            I => \N__25807\
        );

    \I__5269\ : LocalMux
    port map (
            O => \N__25821\,
            I => \N__25807\
        );

    \I__5268\ : LocalMux
    port map (
            O => \N__25818\,
            I => \N__25807\
        );

    \I__5267\ : InMux
    port map (
            O => \N__25817\,
            I => \N__25804\
        );

    \I__5266\ : InMux
    port map (
            O => \N__25816\,
            I => \N__25799\
        );

    \I__5265\ : InMux
    port map (
            O => \N__25815\,
            I => \N__25799\
        );

    \I__5264\ : InMux
    port map (
            O => \N__25814\,
            I => \N__25796\
        );

    \I__5263\ : Span4Mux_h
    port map (
            O => \N__25807\,
            I => \N__25793\
        );

    \I__5262\ : LocalMux
    port map (
            O => \N__25804\,
            I => b2v_inst_state_14
        );

    \I__5261\ : LocalMux
    port map (
            O => \N__25799\,
            I => b2v_inst_state_14
        );

    \I__5260\ : LocalMux
    port map (
            O => \N__25796\,
            I => b2v_inst_state_14
        );

    \I__5259\ : Odrv4
    port map (
            O => \N__25793\,
            I => b2v_inst_state_14
        );

    \I__5258\ : InMux
    port map (
            O => \N__25784\,
            I => \N__25781\
        );

    \I__5257\ : LocalMux
    port map (
            O => \N__25781\,
            I => \b2v_inst.state_ns_a3_i_0_a2_6_1\
        );

    \I__5256\ : CascadeMux
    port map (
            O => \N__25778\,
            I => \b2v_inst9.fsm_state_ns_i_0_i_0_1_cascade_\
        );

    \I__5255\ : InMux
    port map (
            O => \N__25775\,
            I => \N__25771\
        );

    \I__5254\ : InMux
    port map (
            O => \N__25774\,
            I => \N__25768\
        );

    \I__5253\ : LocalMux
    port map (
            O => \N__25771\,
            I => \b2v_inst9.N_832\
        );

    \I__5252\ : LocalMux
    port map (
            O => \N__25768\,
            I => \b2v_inst9.N_832\
        );

    \I__5251\ : CascadeMux
    port map (
            O => \N__25763\,
            I => \N__25760\
        );

    \I__5250\ : InMux
    port map (
            O => \N__25760\,
            I => \N__25757\
        );

    \I__5249\ : LocalMux
    port map (
            O => \N__25757\,
            I => \N__25754\
        );

    \I__5248\ : Span4Mux_h
    port map (
            O => \N__25754\,
            I => \N__25751\
        );

    \I__5247\ : Odrv4
    port map (
            O => \N__25751\,
            I => \b2v_inst9.data_to_sendZ0Z_3\
        );

    \I__5246\ : InMux
    port map (
            O => \N__25748\,
            I => \N__25745\
        );

    \I__5245\ : LocalMux
    port map (
            O => \N__25745\,
            I => \b2v_inst9.data_to_send_10_0_0_0_2\
        );

    \I__5244\ : CascadeMux
    port map (
            O => \N__25742\,
            I => \N__25739\
        );

    \I__5243\ : InMux
    port map (
            O => \N__25739\,
            I => \N__25735\
        );

    \I__5242\ : InMux
    port map (
            O => \N__25738\,
            I => \N__25732\
        );

    \I__5241\ : LocalMux
    port map (
            O => \N__25735\,
            I => \N__25728\
        );

    \I__5240\ : LocalMux
    port map (
            O => \N__25732\,
            I => \N__25725\
        );

    \I__5239\ : CascadeMux
    port map (
            O => \N__25731\,
            I => \N__25718\
        );

    \I__5238\ : Span4Mux_h
    port map (
            O => \N__25728\,
            I => \N__25713\
        );

    \I__5237\ : Span4Mux_h
    port map (
            O => \N__25725\,
            I => \N__25713\
        );

    \I__5236\ : InMux
    port map (
            O => \N__25724\,
            I => \N__25708\
        );

    \I__5235\ : InMux
    port map (
            O => \N__25723\,
            I => \N__25708\
        );

    \I__5234\ : InMux
    port map (
            O => \N__25722\,
            I => \N__25701\
        );

    \I__5233\ : InMux
    port map (
            O => \N__25721\,
            I => \N__25701\
        );

    \I__5232\ : InMux
    port map (
            O => \N__25718\,
            I => \N__25701\
        );

    \I__5231\ : Span4Mux_h
    port map (
            O => \N__25713\,
            I => \N__25698\
        );

    \I__5230\ : LocalMux
    port map (
            O => \N__25708\,
            I => b2v_inst_state_12
        );

    \I__5229\ : LocalMux
    port map (
            O => \N__25701\,
            I => b2v_inst_state_12
        );

    \I__5228\ : Odrv4
    port map (
            O => \N__25698\,
            I => b2v_inst_state_12
        );

    \I__5227\ : InMux
    port map (
            O => \N__25691\,
            I => \N__25688\
        );

    \I__5226\ : LocalMux
    port map (
            O => \N__25688\,
            I => \N__25682\
        );

    \I__5225\ : InMux
    port map (
            O => \N__25687\,
            I => \N__25679\
        );

    \I__5224\ : InMux
    port map (
            O => \N__25686\,
            I => \N__25676\
        );

    \I__5223\ : InMux
    port map (
            O => \N__25685\,
            I => \N__25673\
        );

    \I__5222\ : Span4Mux_v
    port map (
            O => \N__25682\,
            I => \N__25667\
        );

    \I__5221\ : LocalMux
    port map (
            O => \N__25679\,
            I => \N__25667\
        );

    \I__5220\ : LocalMux
    port map (
            O => \N__25676\,
            I => \N__25664\
        );

    \I__5219\ : LocalMux
    port map (
            O => \N__25673\,
            I => \N__25661\
        );

    \I__5218\ : CascadeMux
    port map (
            O => \N__25672\,
            I => \N__25658\
        );

    \I__5217\ : Span4Mux_h
    port map (
            O => \N__25667\,
            I => \N__25655\
        );

    \I__5216\ : Span4Mux_h
    port map (
            O => \N__25664\,
            I => \N__25650\
        );

    \I__5215\ : Span4Mux_h
    port map (
            O => \N__25661\,
            I => \N__25650\
        );

    \I__5214\ : InMux
    port map (
            O => \N__25658\,
            I => \N__25647\
        );

    \I__5213\ : Odrv4
    port map (
            O => \N__25655\,
            I => b2v_inst_state_13
        );

    \I__5212\ : Odrv4
    port map (
            O => \N__25650\,
            I => b2v_inst_state_13
        );

    \I__5211\ : LocalMux
    port map (
            O => \N__25647\,
            I => b2v_inst_state_13
        );

    \I__5210\ : InMux
    port map (
            O => \N__25640\,
            I => \N__25636\
        );

    \I__5209\ : CascadeMux
    port map (
            O => \N__25639\,
            I => \N__25629\
        );

    \I__5208\ : LocalMux
    port map (
            O => \N__25636\,
            I => \N__25625\
        );

    \I__5207\ : InMux
    port map (
            O => \N__25635\,
            I => \N__25617\
        );

    \I__5206\ : InMux
    port map (
            O => \N__25634\,
            I => \N__25617\
        );

    \I__5205\ : InMux
    port map (
            O => \N__25633\,
            I => \N__25617\
        );

    \I__5204\ : InMux
    port map (
            O => \N__25632\,
            I => \N__25614\
        );

    \I__5203\ : InMux
    port map (
            O => \N__25629\,
            I => \N__25609\
        );

    \I__5202\ : InMux
    port map (
            O => \N__25628\,
            I => \N__25609\
        );

    \I__5201\ : Span4Mux_h
    port map (
            O => \N__25625\,
            I => \N__25606\
        );

    \I__5200\ : InMux
    port map (
            O => \N__25624\,
            I => \N__25603\
        );

    \I__5199\ : LocalMux
    port map (
            O => \N__25617\,
            I => \N__25598\
        );

    \I__5198\ : LocalMux
    port map (
            O => \N__25614\,
            I => \N__25598\
        );

    \I__5197\ : LocalMux
    port map (
            O => \N__25609\,
            I => \N__25595\
        );

    \I__5196\ : Span4Mux_v
    port map (
            O => \N__25606\,
            I => \N__25590\
        );

    \I__5195\ : LocalMux
    port map (
            O => \N__25603\,
            I => \N__25590\
        );

    \I__5194\ : Span4Mux_h
    port map (
            O => \N__25598\,
            I => \N__25587\
        );

    \I__5193\ : Span4Mux_h
    port map (
            O => \N__25595\,
            I => \N__25584\
        );

    \I__5192\ : Odrv4
    port map (
            O => \N__25590\,
            I => \b2v_inst9.N_739\
        );

    \I__5191\ : Odrv4
    port map (
            O => \N__25587\,
            I => \b2v_inst9.N_739\
        );

    \I__5190\ : Odrv4
    port map (
            O => \N__25584\,
            I => \b2v_inst9.N_739\
        );

    \I__5189\ : InMux
    port map (
            O => \N__25577\,
            I => \N__25574\
        );

    \I__5188\ : LocalMux
    port map (
            O => \N__25574\,
            I => \b2v_inst.pix_data_regZ0Z_0\
        );

    \I__5187\ : InMux
    port map (
            O => \N__25571\,
            I => \N__25568\
        );

    \I__5186\ : LocalMux
    port map (
            O => \N__25568\,
            I => \b2v_inst.pix_data_regZ0Z_1\
        );

    \I__5185\ : InMux
    port map (
            O => \N__25565\,
            I => \b2v_inst.eventos_cry_6\
        );

    \I__5184\ : InMux
    port map (
            O => \N__25562\,
            I => \bfn_15_11_0_\
        );

    \I__5183\ : InMux
    port map (
            O => \N__25559\,
            I => \b2v_inst.eventos_cry_8\
        );

    \I__5182\ : InMux
    port map (
            O => \N__25556\,
            I => \b2v_inst.eventos_cry_9\
        );

    \I__5181\ : InMux
    port map (
            O => \N__25553\,
            I => \N__25550\
        );

    \I__5180\ : LocalMux
    port map (
            O => \N__25550\,
            I => \N__25547\
        );

    \I__5179\ : Span4Mux_h
    port map (
            O => \N__25547\,
            I => \N__25544\
        );

    \I__5178\ : Odrv4
    port map (
            O => \N__25544\,
            I => \b2v_inst.state_ns_a3_i_0_a2_5_1\
        );

    \I__5177\ : CascadeMux
    port map (
            O => \N__25541\,
            I => \b2v_inst.state_ns_a3_i_0_a2_4_1_cascade_\
        );

    \I__5176\ : InMux
    port map (
            O => \N__25538\,
            I => \N__25532\
        );

    \I__5175\ : InMux
    port map (
            O => \N__25537\,
            I => \N__25532\
        );

    \I__5174\ : LocalMux
    port map (
            O => \N__25532\,
            I => \N__25525\
        );

    \I__5173\ : CascadeMux
    port map (
            O => \N__25531\,
            I => \N__25521\
        );

    \I__5172\ : InMux
    port map (
            O => \N__25530\,
            I => \N__25516\
        );

    \I__5171\ : InMux
    port map (
            O => \N__25529\,
            I => \N__25516\
        );

    \I__5170\ : InMux
    port map (
            O => \N__25528\,
            I => \N__25513\
        );

    \I__5169\ : Span4Mux_v
    port map (
            O => \N__25525\,
            I => \N__25510\
        );

    \I__5168\ : InMux
    port map (
            O => \N__25524\,
            I => \N__25505\
        );

    \I__5167\ : InMux
    port map (
            O => \N__25521\,
            I => \N__25505\
        );

    \I__5166\ : LocalMux
    port map (
            O => \N__25516\,
            I => \N__25502\
        );

    \I__5165\ : LocalMux
    port map (
            O => \N__25513\,
            I => \N__25495\
        );

    \I__5164\ : Span4Mux_h
    port map (
            O => \N__25510\,
            I => \N__25495\
        );

    \I__5163\ : LocalMux
    port map (
            O => \N__25505\,
            I => \N__25495\
        );

    \I__5162\ : Span4Mux_h
    port map (
            O => \N__25502\,
            I => \N__25492\
        );

    \I__5161\ : Span4Mux_h
    port map (
            O => \N__25495\,
            I => \N__25489\
        );

    \I__5160\ : Odrv4
    port map (
            O => \N__25492\,
            I => \b2v_inst.stateZ0Z_31\
        );

    \I__5159\ : Odrv4
    port map (
            O => \N__25489\,
            I => \b2v_inst.stateZ0Z_31\
        );

    \I__5158\ : InMux
    port map (
            O => \N__25484\,
            I => \N__25480\
        );

    \I__5157\ : CascadeMux
    port map (
            O => \N__25483\,
            I => \N__25477\
        );

    \I__5156\ : LocalMux
    port map (
            O => \N__25480\,
            I => \N__25474\
        );

    \I__5155\ : InMux
    port map (
            O => \N__25477\,
            I => \N__25471\
        );

    \I__5154\ : Span4Mux_h
    port map (
            O => \N__25474\,
            I => \N__25464\
        );

    \I__5153\ : LocalMux
    port map (
            O => \N__25471\,
            I => \N__25464\
        );

    \I__5152\ : InMux
    port map (
            O => \N__25470\,
            I => \N__25459\
        );

    \I__5151\ : InMux
    port map (
            O => \N__25469\,
            I => \N__25459\
        );

    \I__5150\ : Span4Mux_h
    port map (
            O => \N__25464\,
            I => \N__25454\
        );

    \I__5149\ : LocalMux
    port map (
            O => \N__25459\,
            I => \N__25451\
        );

    \I__5148\ : InMux
    port map (
            O => \N__25458\,
            I => \N__25446\
        );

    \I__5147\ : InMux
    port map (
            O => \N__25457\,
            I => \N__25446\
        );

    \I__5146\ : Odrv4
    port map (
            O => \N__25454\,
            I => b2v_inst_state_7
        );

    \I__5145\ : Odrv12
    port map (
            O => \N__25451\,
            I => b2v_inst_state_7
        );

    \I__5144\ : LocalMux
    port map (
            O => \N__25446\,
            I => b2v_inst_state_7
        );

    \I__5143\ : InMux
    port map (
            O => \N__25439\,
            I => \N__25434\
        );

    \I__5142\ : InMux
    port map (
            O => \N__25438\,
            I => \N__25431\
        );

    \I__5141\ : InMux
    port map (
            O => \N__25437\,
            I => \N__25428\
        );

    \I__5140\ : LocalMux
    port map (
            O => \N__25434\,
            I => \N__25423\
        );

    \I__5139\ : LocalMux
    port map (
            O => \N__25431\,
            I => \N__25423\
        );

    \I__5138\ : LocalMux
    port map (
            O => \N__25428\,
            I => \N__25420\
        );

    \I__5137\ : Span4Mux_h
    port map (
            O => \N__25423\,
            I => \N__25413\
        );

    \I__5136\ : Span4Mux_v
    port map (
            O => \N__25420\,
            I => \N__25410\
        );

    \I__5135\ : InMux
    port map (
            O => \N__25419\,
            I => \N__25407\
        );

    \I__5134\ : InMux
    port map (
            O => \N__25418\,
            I => \N__25400\
        );

    \I__5133\ : InMux
    port map (
            O => \N__25417\,
            I => \N__25400\
        );

    \I__5132\ : InMux
    port map (
            O => \N__25416\,
            I => \N__25400\
        );

    \I__5131\ : Span4Mux_h
    port map (
            O => \N__25413\,
            I => \N__25397\
        );

    \I__5130\ : Odrv4
    port map (
            O => \N__25410\,
            I => b2v_inst_state_1
        );

    \I__5129\ : LocalMux
    port map (
            O => \N__25407\,
            I => b2v_inst_state_1
        );

    \I__5128\ : LocalMux
    port map (
            O => \N__25400\,
            I => b2v_inst_state_1
        );

    \I__5127\ : Odrv4
    port map (
            O => \N__25397\,
            I => b2v_inst_state_1
        );

    \I__5126\ : InMux
    port map (
            O => \N__25388\,
            I => \N__25385\
        );

    \I__5125\ : LocalMux
    port map (
            O => \N__25385\,
            I => \b2v_inst.data_a_escribir11_8_and\
        );

    \I__5124\ : InMux
    port map (
            O => \N__25382\,
            I => \N__25379\
        );

    \I__5123\ : LocalMux
    port map (
            O => \N__25379\,
            I => \N__25376\
        );

    \I__5122\ : Span4Mux_h
    port map (
            O => \N__25376\,
            I => \N__25373\
        );

    \I__5121\ : Span4Mux_h
    port map (
            O => \N__25373\,
            I => \N__25370\
        );

    \I__5120\ : Odrv4
    port map (
            O => \N__25370\,
            I => \b2v_inst.dir_mem_1Z0Z_10\
        );

    \I__5119\ : InMux
    port map (
            O => \N__25367\,
            I => \N__25360\
        );

    \I__5118\ : CascadeMux
    port map (
            O => \N__25366\,
            I => \N__25355\
        );

    \I__5117\ : InMux
    port map (
            O => \N__25365\,
            I => \N__25350\
        );

    \I__5116\ : InMux
    port map (
            O => \N__25364\,
            I => \N__25350\
        );

    \I__5115\ : CascadeMux
    port map (
            O => \N__25363\,
            I => \N__25344\
        );

    \I__5114\ : LocalMux
    port map (
            O => \N__25360\,
            I => \N__25341\
        );

    \I__5113\ : InMux
    port map (
            O => \N__25359\,
            I => \N__25336\
        );

    \I__5112\ : InMux
    port map (
            O => \N__25358\,
            I => \N__25333\
        );

    \I__5111\ : InMux
    port map (
            O => \N__25355\,
            I => \N__25330\
        );

    \I__5110\ : LocalMux
    port map (
            O => \N__25350\,
            I => \N__25327\
        );

    \I__5109\ : InMux
    port map (
            O => \N__25349\,
            I => \N__25324\
        );

    \I__5108\ : InMux
    port map (
            O => \N__25348\,
            I => \N__25321\
        );

    \I__5107\ : InMux
    port map (
            O => \N__25347\,
            I => \N__25316\
        );

    \I__5106\ : InMux
    port map (
            O => \N__25344\,
            I => \N__25316\
        );

    \I__5105\ : Span4Mux_h
    port map (
            O => \N__25341\,
            I => \N__25313\
        );

    \I__5104\ : InMux
    port map (
            O => \N__25340\,
            I => \N__25308\
        );

    \I__5103\ : InMux
    port map (
            O => \N__25339\,
            I => \N__25308\
        );

    \I__5102\ : LocalMux
    port map (
            O => \N__25336\,
            I => \N__25301\
        );

    \I__5101\ : LocalMux
    port map (
            O => \N__25333\,
            I => \N__25301\
        );

    \I__5100\ : LocalMux
    port map (
            O => \N__25330\,
            I => \N__25301\
        );

    \I__5099\ : Odrv4
    port map (
            O => \N__25327\,
            I => \b2v_inst.N_490\
        );

    \I__5098\ : LocalMux
    port map (
            O => \N__25324\,
            I => \b2v_inst.N_490\
        );

    \I__5097\ : LocalMux
    port map (
            O => \N__25321\,
            I => \b2v_inst.N_490\
        );

    \I__5096\ : LocalMux
    port map (
            O => \N__25316\,
            I => \b2v_inst.N_490\
        );

    \I__5095\ : Odrv4
    port map (
            O => \N__25313\,
            I => \b2v_inst.N_490\
        );

    \I__5094\ : LocalMux
    port map (
            O => \N__25308\,
            I => \b2v_inst.N_490\
        );

    \I__5093\ : Odrv4
    port map (
            O => \N__25301\,
            I => \b2v_inst.N_490\
        );

    \I__5092\ : CascadeMux
    port map (
            O => \N__25286\,
            I => \N__25283\
        );

    \I__5091\ : InMux
    port map (
            O => \N__25283\,
            I => \N__25280\
        );

    \I__5090\ : LocalMux
    port map (
            O => \N__25280\,
            I => \N__25277\
        );

    \I__5089\ : Span4Mux_v
    port map (
            O => \N__25277\,
            I => \N__25274\
        );

    \I__5088\ : Span4Mux_h
    port map (
            O => \N__25274\,
            I => \N__25271\
        );

    \I__5087\ : Odrv4
    port map (
            O => \N__25271\,
            I => \b2v_inst.dir_mem_3Z0Z_10\
        );

    \I__5086\ : InMux
    port map (
            O => \N__25268\,
            I => \N__25264\
        );

    \I__5085\ : InMux
    port map (
            O => \N__25267\,
            I => \N__25261\
        );

    \I__5084\ : LocalMux
    port map (
            O => \N__25264\,
            I => \N__25250\
        );

    \I__5083\ : LocalMux
    port map (
            O => \N__25261\,
            I => \N__25245\
        );

    \I__5082\ : InMux
    port map (
            O => \N__25260\,
            I => \N__25242\
        );

    \I__5081\ : InMux
    port map (
            O => \N__25259\,
            I => \N__25237\
        );

    \I__5080\ : InMux
    port map (
            O => \N__25258\,
            I => \N__25237\
        );

    \I__5079\ : InMux
    port map (
            O => \N__25257\,
            I => \N__25234\
        );

    \I__5078\ : InMux
    port map (
            O => \N__25256\,
            I => \N__25231\
        );

    \I__5077\ : InMux
    port map (
            O => \N__25255\,
            I => \N__25228\
        );

    \I__5076\ : InMux
    port map (
            O => \N__25254\,
            I => \N__25225\
        );

    \I__5075\ : InMux
    port map (
            O => \N__25253\,
            I => \N__25222\
        );

    \I__5074\ : Span4Mux_h
    port map (
            O => \N__25250\,
            I => \N__25219\
        );

    \I__5073\ : InMux
    port map (
            O => \N__25249\,
            I => \N__25214\
        );

    \I__5072\ : InMux
    port map (
            O => \N__25248\,
            I => \N__25214\
        );

    \I__5071\ : Span4Mux_h
    port map (
            O => \N__25245\,
            I => \N__25207\
        );

    \I__5070\ : LocalMux
    port map (
            O => \N__25242\,
            I => \N__25207\
        );

    \I__5069\ : LocalMux
    port map (
            O => \N__25237\,
            I => \N__25207\
        );

    \I__5068\ : LocalMux
    port map (
            O => \N__25234\,
            I => \N__25202\
        );

    \I__5067\ : LocalMux
    port map (
            O => \N__25231\,
            I => \N__25202\
        );

    \I__5066\ : LocalMux
    port map (
            O => \N__25228\,
            I => \b2v_inst.N_488\
        );

    \I__5065\ : LocalMux
    port map (
            O => \N__25225\,
            I => \b2v_inst.N_488\
        );

    \I__5064\ : LocalMux
    port map (
            O => \N__25222\,
            I => \b2v_inst.N_488\
        );

    \I__5063\ : Odrv4
    port map (
            O => \N__25219\,
            I => \b2v_inst.N_488\
        );

    \I__5062\ : LocalMux
    port map (
            O => \N__25214\,
            I => \b2v_inst.N_488\
        );

    \I__5061\ : Odrv4
    port map (
            O => \N__25207\,
            I => \b2v_inst.N_488\
        );

    \I__5060\ : Odrv4
    port map (
            O => \N__25202\,
            I => \b2v_inst.N_488\
        );

    \I__5059\ : InMux
    port map (
            O => \N__25187\,
            I => \bfn_15_10_0_\
        );

    \I__5058\ : InMux
    port map (
            O => \N__25184\,
            I => \b2v_inst.eventos_cry_0\
        );

    \I__5057\ : InMux
    port map (
            O => \N__25181\,
            I => \b2v_inst.eventos_cry_1\
        );

    \I__5056\ : InMux
    port map (
            O => \N__25178\,
            I => \b2v_inst.eventos_cry_2\
        );

    \I__5055\ : InMux
    port map (
            O => \N__25175\,
            I => \b2v_inst.eventos_cry_3\
        );

    \I__5054\ : InMux
    port map (
            O => \N__25172\,
            I => \b2v_inst.eventos_cry_4\
        );

    \I__5053\ : InMux
    port map (
            O => \N__25169\,
            I => \b2v_inst.eventos_cry_5\
        );

    \I__5052\ : InMux
    port map (
            O => \N__25166\,
            I => \N__25163\
        );

    \I__5051\ : LocalMux
    port map (
            O => \N__25163\,
            I => \b2v_inst.data_a_escribir11_4_and\
        );

    \I__5050\ : InMux
    port map (
            O => \N__25160\,
            I => \b2v_inst.data_a_escribir12\
        );

    \I__5049\ : InMux
    port map (
            O => \N__25157\,
            I => \N__25154\
        );

    \I__5048\ : LocalMux
    port map (
            O => \N__25154\,
            I => \b2v_inst.data_a_escribir11_9_and\
        );

    \I__5047\ : InMux
    port map (
            O => \N__25151\,
            I => \N__25148\
        );

    \I__5046\ : LocalMux
    port map (
            O => \N__25148\,
            I => \b2v_inst.data_a_escribir11_2_and\
        );

    \I__5045\ : CascadeMux
    port map (
            O => \N__25145\,
            I => \N__25142\
        );

    \I__5044\ : InMux
    port map (
            O => \N__25142\,
            I => \N__25138\
        );

    \I__5043\ : InMux
    port map (
            O => \N__25141\,
            I => \N__25135\
        );

    \I__5042\ : LocalMux
    port map (
            O => \N__25138\,
            I => \N__25132\
        );

    \I__5041\ : LocalMux
    port map (
            O => \N__25135\,
            I => \N__25129\
        );

    \I__5040\ : Span4Mux_v
    port map (
            O => \N__25132\,
            I => \N__25126\
        );

    \I__5039\ : Span4Mux_h
    port map (
            O => \N__25129\,
            I => \N__25123\
        );

    \I__5038\ : Span4Mux_h
    port map (
            O => \N__25126\,
            I => \N__25120\
        );

    \I__5037\ : Span4Mux_h
    port map (
            O => \N__25123\,
            I => \N__25117\
        );

    \I__5036\ : Odrv4
    port map (
            O => \N__25120\,
            I => b2v_inst_energia_temp_10
        );

    \I__5035\ : Odrv4
    port map (
            O => \N__25117\,
            I => b2v_inst_energia_temp_10
        );

    \I__5034\ : InMux
    port map (
            O => \N__25112\,
            I => \b2v_inst.un14_data_ram_energia_o_cry_9\
        );

    \I__5033\ : InMux
    port map (
            O => \N__25109\,
            I => \N__25106\
        );

    \I__5032\ : LocalMux
    port map (
            O => \N__25106\,
            I => \N__25102\
        );

    \I__5031\ : InMux
    port map (
            O => \N__25105\,
            I => \N__25099\
        );

    \I__5030\ : Span4Mux_v
    port map (
            O => \N__25102\,
            I => \N__25096\
        );

    \I__5029\ : LocalMux
    port map (
            O => \N__25099\,
            I => \N__25093\
        );

    \I__5028\ : Span4Mux_v
    port map (
            O => \N__25096\,
            I => \N__25088\
        );

    \I__5027\ : Span4Mux_h
    port map (
            O => \N__25093\,
            I => \N__25088\
        );

    \I__5026\ : Span4Mux_h
    port map (
            O => \N__25088\,
            I => \N__25085\
        );

    \I__5025\ : Odrv4
    port map (
            O => \N__25085\,
            I => b2v_inst_energia_temp_11
        );

    \I__5024\ : InMux
    port map (
            O => \N__25082\,
            I => \N__25079\
        );

    \I__5023\ : LocalMux
    port map (
            O => \N__25079\,
            I => \N__25076\
        );

    \I__5022\ : Span4Mux_v
    port map (
            O => \N__25076\,
            I => \N__25073\
        );

    \I__5021\ : Span4Mux_h
    port map (
            O => \N__25073\,
            I => \N__25070\
        );

    \I__5020\ : Span4Mux_h
    port map (
            O => \N__25070\,
            I => \N__25067\
        );

    \I__5019\ : Odrv4
    port map (
            O => \N__25067\,
            I => \SYNTHESIZED_WIRE_13_11\
        );

    \I__5018\ : InMux
    port map (
            O => \N__25064\,
            I => \b2v_inst.un14_data_ram_energia_o_cry_10\
        );

    \I__5017\ : InMux
    port map (
            O => \N__25061\,
            I => \N__25058\
        );

    \I__5016\ : LocalMux
    port map (
            O => \N__25058\,
            I => \N__25054\
        );

    \I__5015\ : InMux
    port map (
            O => \N__25057\,
            I => \N__25051\
        );

    \I__5014\ : Span4Mux_h
    port map (
            O => \N__25054\,
            I => \N__25048\
        );

    \I__5013\ : LocalMux
    port map (
            O => \N__25051\,
            I => \N__25045\
        );

    \I__5012\ : Span4Mux_v
    port map (
            O => \N__25048\,
            I => \N__25042\
        );

    \I__5011\ : Span4Mux_h
    port map (
            O => \N__25045\,
            I => \N__25039\
        );

    \I__5010\ : Odrv4
    port map (
            O => \N__25042\,
            I => b2v_inst_energia_temp_12
        );

    \I__5009\ : Odrv4
    port map (
            O => \N__25039\,
            I => b2v_inst_energia_temp_12
        );

    \I__5008\ : InMux
    port map (
            O => \N__25034\,
            I => \N__25031\
        );

    \I__5007\ : LocalMux
    port map (
            O => \N__25031\,
            I => \N__25028\
        );

    \I__5006\ : Span4Mux_v
    port map (
            O => \N__25028\,
            I => \N__25025\
        );

    \I__5005\ : Span4Mux_v
    port map (
            O => \N__25025\,
            I => \N__25022\
        );

    \I__5004\ : Sp12to4
    port map (
            O => \N__25022\,
            I => \N__25019\
        );

    \I__5003\ : Odrv12
    port map (
            O => \N__25019\,
            I => \SYNTHESIZED_WIRE_13_12\
        );

    \I__5002\ : InMux
    port map (
            O => \N__25016\,
            I => \b2v_inst.un14_data_ram_energia_o_cry_11\
        );

    \I__5001\ : InMux
    port map (
            O => \N__25013\,
            I => \N__25010\
        );

    \I__5000\ : LocalMux
    port map (
            O => \N__25010\,
            I => \N__25006\
        );

    \I__4999\ : InMux
    port map (
            O => \N__25009\,
            I => \N__25003\
        );

    \I__4998\ : Span4Mux_h
    port map (
            O => \N__25006\,
            I => \N__25000\
        );

    \I__4997\ : LocalMux
    port map (
            O => \N__25003\,
            I => b2v_inst_energia_temp_13
        );

    \I__4996\ : Odrv4
    port map (
            O => \N__25000\,
            I => b2v_inst_energia_temp_13
        );

    \I__4995\ : InMux
    port map (
            O => \N__24995\,
            I => \b2v_inst.un14_data_ram_energia_o_cry_12\
        );

    \I__4994\ : InMux
    port map (
            O => \N__24992\,
            I => \N__24989\
        );

    \I__4993\ : LocalMux
    port map (
            O => \N__24989\,
            I => \N__24986\
        );

    \I__4992\ : Span4Mux_v
    port map (
            O => \N__24986\,
            I => \N__24983\
        );

    \I__4991\ : Sp12to4
    port map (
            O => \N__24983\,
            I => \N__24980\
        );

    \I__4990\ : Odrv12
    port map (
            O => \N__24980\,
            I => \SYNTHESIZED_WIRE_13_13\
        );

    \I__4989\ : IoInMux
    port map (
            O => \N__24977\,
            I => \N__24973\
        );

    \I__4988\ : InMux
    port map (
            O => \N__24976\,
            I => \N__24970\
        );

    \I__4987\ : LocalMux
    port map (
            O => \N__24973\,
            I => \N__24967\
        );

    \I__4986\ : LocalMux
    port map (
            O => \N__24970\,
            I => \N__24964\
        );

    \I__4985\ : Span4Mux_s3_h
    port map (
            O => \N__24967\,
            I => \N__24961\
        );

    \I__4984\ : Span4Mux_v
    port map (
            O => \N__24964\,
            I => \N__24958\
        );

    \I__4983\ : Span4Mux_h
    port map (
            O => \N__24961\,
            I => \N__24955\
        );

    \I__4982\ : Sp12to4
    port map (
            O => \N__24958\,
            I => \N__24952\
        );

    \I__4981\ : Odrv4
    port map (
            O => \N__24955\,
            I => leds_c_8
        );

    \I__4980\ : Odrv12
    port map (
            O => \N__24952\,
            I => leds_c_8
        );

    \I__4979\ : InMux
    port map (
            O => \N__24947\,
            I => \N__24944\
        );

    \I__4978\ : LocalMux
    port map (
            O => \N__24944\,
            I => \N__24940\
        );

    \I__4977\ : InMux
    port map (
            O => \N__24943\,
            I => \N__24937\
        );

    \I__4976\ : Odrv4
    port map (
            O => \N__24940\,
            I => b2v_inst_energia_temp_8
        );

    \I__4975\ : LocalMux
    port map (
            O => \N__24937\,
            I => b2v_inst_energia_temp_8
        );

    \I__4974\ : InMux
    port map (
            O => \N__24932\,
            I => \N__24929\
        );

    \I__4973\ : LocalMux
    port map (
            O => \N__24929\,
            I => \b2v_inst.un14_data_ram_energia_o_cry_9_c_RNI28GBZ0\
        );

    \I__4972\ : InMux
    port map (
            O => \N__24926\,
            I => \N__24923\
        );

    \I__4971\ : LocalMux
    port map (
            O => \N__24923\,
            I => \N__24920\
        );

    \I__4970\ : Span4Mux_h
    port map (
            O => \N__24920\,
            I => \N__24917\
        );

    \I__4969\ : Span4Mux_h
    port map (
            O => \N__24917\,
            I => \N__24914\
        );

    \I__4968\ : Span4Mux_h
    port map (
            O => \N__24914\,
            I => \N__24911\
        );

    \I__4967\ : Odrv4
    port map (
            O => \N__24911\,
            I => \N_461_i\
        );

    \I__4966\ : CascadeMux
    port map (
            O => \N__24908\,
            I => \N__24904\
        );

    \I__4965\ : InMux
    port map (
            O => \N__24907\,
            I => \N__24901\
        );

    \I__4964\ : InMux
    port map (
            O => \N__24904\,
            I => \N__24898\
        );

    \I__4963\ : LocalMux
    port map (
            O => \N__24901\,
            I => b2v_inst_energia_temp_2
        );

    \I__4962\ : LocalMux
    port map (
            O => \N__24898\,
            I => b2v_inst_energia_temp_2
        );

    \I__4961\ : InMux
    port map (
            O => \N__24893\,
            I => \N__24890\
        );

    \I__4960\ : LocalMux
    port map (
            O => \N__24890\,
            I => \N__24887\
        );

    \I__4959\ : Odrv4
    port map (
            O => \N__24887\,
            I => \b2v_inst.un14_data_ram_energia_o_cry_1_c_RNIHM5MZ0\
        );

    \I__4958\ : InMux
    port map (
            O => \N__24884\,
            I => \b2v_inst.un14_data_ram_energia_o_cry_1\
        );

    \I__4957\ : CascadeMux
    port map (
            O => \N__24881\,
            I => \N__24877\
        );

    \I__4956\ : InMux
    port map (
            O => \N__24880\,
            I => \N__24874\
        );

    \I__4955\ : InMux
    port map (
            O => \N__24877\,
            I => \N__24871\
        );

    \I__4954\ : LocalMux
    port map (
            O => \N__24874\,
            I => b2v_inst_energia_temp_3
        );

    \I__4953\ : LocalMux
    port map (
            O => \N__24871\,
            I => b2v_inst_energia_temp_3
        );

    \I__4952\ : InMux
    port map (
            O => \N__24866\,
            I => \N__24863\
        );

    \I__4951\ : LocalMux
    port map (
            O => \N__24863\,
            I => \N__24860\
        );

    \I__4950\ : Odrv4
    port map (
            O => \N__24860\,
            I => \b2v_inst.un14_data_ram_energia_o_cry_2_c_RNIKQ6MZ0\
        );

    \I__4949\ : InMux
    port map (
            O => \N__24857\,
            I => \b2v_inst.un14_data_ram_energia_o_cry_2\
        );

    \I__4948\ : InMux
    port map (
            O => \N__24854\,
            I => \N__24851\
        );

    \I__4947\ : LocalMux
    port map (
            O => \N__24851\,
            I => \N__24848\
        );

    \I__4946\ : Span4Mux_v
    port map (
            O => \N__24848\,
            I => \N__24845\
        );

    \I__4945\ : Span4Mux_h
    port map (
            O => \N__24845\,
            I => \N__24842\
        );

    \I__4944\ : Span4Mux_h
    port map (
            O => \N__24842\,
            I => \N__24839\
        );

    \I__4943\ : Odrv4
    port map (
            O => \N__24839\,
            I => \b2v_inst.pix_data_regZ0Z_4\
        );

    \I__4942\ : CascadeMux
    port map (
            O => \N__24836\,
            I => \N__24832\
        );

    \I__4941\ : InMux
    port map (
            O => \N__24835\,
            I => \N__24829\
        );

    \I__4940\ : InMux
    port map (
            O => \N__24832\,
            I => \N__24826\
        );

    \I__4939\ : LocalMux
    port map (
            O => \N__24829\,
            I => \N__24823\
        );

    \I__4938\ : LocalMux
    port map (
            O => \N__24826\,
            I => \N__24820\
        );

    \I__4937\ : Span4Mux_v
    port map (
            O => \N__24823\,
            I => \N__24815\
        );

    \I__4936\ : Span4Mux_v
    port map (
            O => \N__24820\,
            I => \N__24815\
        );

    \I__4935\ : Span4Mux_h
    port map (
            O => \N__24815\,
            I => \N__24812\
        );

    \I__4934\ : Span4Mux_v
    port map (
            O => \N__24812\,
            I => \N__24809\
        );

    \I__4933\ : Odrv4
    port map (
            O => \N__24809\,
            I => b2v_inst_energia_temp_4
        );

    \I__4932\ : InMux
    port map (
            O => \N__24806\,
            I => \N__24803\
        );

    \I__4931\ : LocalMux
    port map (
            O => \N__24803\,
            I => \N__24800\
        );

    \I__4930\ : Span4Mux_h
    port map (
            O => \N__24800\,
            I => \N__24797\
        );

    \I__4929\ : Odrv4
    port map (
            O => \N__24797\,
            I => \b2v_inst.un14_data_ram_energia_o_cry_3_c_RNINU7MZ0\
        );

    \I__4928\ : InMux
    port map (
            O => \N__24794\,
            I => \b2v_inst.un14_data_ram_energia_o_cry_3\
        );

    \I__4927\ : InMux
    port map (
            O => \N__24791\,
            I => \N__24787\
        );

    \I__4926\ : InMux
    port map (
            O => \N__24790\,
            I => \N__24784\
        );

    \I__4925\ : LocalMux
    port map (
            O => \N__24787\,
            I => \N__24779\
        );

    \I__4924\ : LocalMux
    port map (
            O => \N__24784\,
            I => \N__24779\
        );

    \I__4923\ : Span12Mux_v
    port map (
            O => \N__24779\,
            I => \N__24776\
        );

    \I__4922\ : Odrv12
    port map (
            O => \N__24776\,
            I => b2v_inst_energia_temp_5
        );

    \I__4921\ : InMux
    port map (
            O => \N__24773\,
            I => \N__24770\
        );

    \I__4920\ : LocalMux
    port map (
            O => \N__24770\,
            I => \b2v_inst.un14_data_ram_energia_o_cry_4_c_RNIQ29MZ0\
        );

    \I__4919\ : InMux
    port map (
            O => \N__24767\,
            I => \b2v_inst.un14_data_ram_energia_o_cry_4\
        );

    \I__4918\ : InMux
    port map (
            O => \N__24764\,
            I => \N__24760\
        );

    \I__4917\ : CascadeMux
    port map (
            O => \N__24763\,
            I => \N__24757\
        );

    \I__4916\ : LocalMux
    port map (
            O => \N__24760\,
            I => \N__24754\
        );

    \I__4915\ : InMux
    port map (
            O => \N__24757\,
            I => \N__24751\
        );

    \I__4914\ : Span4Mux_v
    port map (
            O => \N__24754\,
            I => \N__24746\
        );

    \I__4913\ : LocalMux
    port map (
            O => \N__24751\,
            I => \N__24746\
        );

    \I__4912\ : Span4Mux_h
    port map (
            O => \N__24746\,
            I => \N__24743\
        );

    \I__4911\ : Odrv4
    port map (
            O => \N__24743\,
            I => b2v_inst_energia_temp_6
        );

    \I__4910\ : InMux
    port map (
            O => \N__24740\,
            I => \N__24737\
        );

    \I__4909\ : LocalMux
    port map (
            O => \N__24737\,
            I => \N__24734\
        );

    \I__4908\ : Odrv12
    port map (
            O => \N__24734\,
            I => \b2v_inst.un14_data_ram_energia_o_cry_5_c_RNIT6AMZ0\
        );

    \I__4907\ : InMux
    port map (
            O => \N__24731\,
            I => \b2v_inst.un14_data_ram_energia_o_cry_5\
        );

    \I__4906\ : InMux
    port map (
            O => \N__24728\,
            I => \N__24724\
        );

    \I__4905\ : CascadeMux
    port map (
            O => \N__24727\,
            I => \N__24721\
        );

    \I__4904\ : LocalMux
    port map (
            O => \N__24724\,
            I => \N__24718\
        );

    \I__4903\ : InMux
    port map (
            O => \N__24721\,
            I => \N__24715\
        );

    \I__4902\ : Span4Mux_v
    port map (
            O => \N__24718\,
            I => \N__24710\
        );

    \I__4901\ : LocalMux
    port map (
            O => \N__24715\,
            I => \N__24710\
        );

    \I__4900\ : Span4Mux_v
    port map (
            O => \N__24710\,
            I => \N__24707\
        );

    \I__4899\ : Span4Mux_h
    port map (
            O => \N__24707\,
            I => \N__24704\
        );

    \I__4898\ : Odrv4
    port map (
            O => \N__24704\,
            I => b2v_inst_energia_temp_7
        );

    \I__4897\ : InMux
    port map (
            O => \N__24701\,
            I => \N__24698\
        );

    \I__4896\ : LocalMux
    port map (
            O => \N__24698\,
            I => \b2v_inst.un14_data_ram_energia_o_cry_6_c_RNI0BBMZ0\
        );

    \I__4895\ : InMux
    port map (
            O => \N__24695\,
            I => \b2v_inst.un14_data_ram_energia_o_cry_6\
        );

    \I__4894\ : InMux
    port map (
            O => \N__24692\,
            I => \N__24689\
        );

    \I__4893\ : LocalMux
    port map (
            O => \N__24689\,
            I => \N__24686\
        );

    \I__4892\ : Span4Mux_h
    port map (
            O => \N__24686\,
            I => \N__24683\
        );

    \I__4891\ : Odrv4
    port map (
            O => \N__24683\,
            I => \b2v_inst.un14_data_ram_energia_o_cry_7_c_RNIN84CZ0\
        );

    \I__4890\ : InMux
    port map (
            O => \N__24680\,
            I => \bfn_14_15_0_\
        );

    \I__4889\ : InMux
    port map (
            O => \N__24677\,
            I => \N__24674\
        );

    \I__4888\ : LocalMux
    port map (
            O => \N__24674\,
            I => \N__24671\
        );

    \I__4887\ : Span4Mux_h
    port map (
            O => \N__24671\,
            I => \N__24668\
        );

    \I__4886\ : Odrv4
    port map (
            O => \N__24668\,
            I => \b2v_inst.un14_data_ram_energia_o_cry_8_c_RNIPB5CZ0\
        );

    \I__4885\ : InMux
    port map (
            O => \N__24665\,
            I => \b2v_inst.un14_data_ram_energia_o_cry_8\
        );

    \I__4884\ : InMux
    port map (
            O => \N__24662\,
            I => \N__24653\
        );

    \I__4883\ : InMux
    port map (
            O => \N__24661\,
            I => \N__24653\
        );

    \I__4882\ : InMux
    port map (
            O => \N__24660\,
            I => \N__24650\
        );

    \I__4881\ : InMux
    port map (
            O => \N__24659\,
            I => \N__24647\
        );

    \I__4880\ : InMux
    port map (
            O => \N__24658\,
            I => \N__24644\
        );

    \I__4879\ : LocalMux
    port map (
            O => \N__24653\,
            I => \N__24639\
        );

    \I__4878\ : LocalMux
    port map (
            O => \N__24650\,
            I => \N__24639\
        );

    \I__4877\ : LocalMux
    port map (
            O => \N__24647\,
            I => \N__24634\
        );

    \I__4876\ : LocalMux
    port map (
            O => \N__24644\,
            I => \N__24634\
        );

    \I__4875\ : Span4Mux_h
    port map (
            O => \N__24639\,
            I => \N__24629\
        );

    \I__4874\ : Span4Mux_h
    port map (
            O => \N__24634\,
            I => \N__24629\
        );

    \I__4873\ : Odrv4
    port map (
            O => \N__24629\,
            I => b2v_inst_state_15
        );

    \I__4872\ : CascadeMux
    port map (
            O => \N__24626\,
            I => \b2v_inst9.N_832_cascade_\
        );

    \I__4871\ : InMux
    port map (
            O => \N__24623\,
            I => \N__24620\
        );

    \I__4870\ : LocalMux
    port map (
            O => \N__24620\,
            I => \N__24617\
        );

    \I__4869\ : Odrv12
    port map (
            O => \N__24617\,
            I => \b2v_inst9.data_to_send_10_0_0_0_1\
        );

    \I__4868\ : InMux
    port map (
            O => \N__24614\,
            I => \N__24611\
        );

    \I__4867\ : LocalMux
    port map (
            O => \N__24611\,
            I => \N__24608\
        );

    \I__4866\ : Odrv12
    port map (
            O => \N__24608\,
            I => \b2v_inst9.data_to_send_10_0_0_1_1\
        );

    \I__4865\ : CascadeMux
    port map (
            O => \N__24605\,
            I => \b2v_inst9.data_to_send_10_0_0_2_2_cascade_\
        );

    \I__4864\ : InMux
    port map (
            O => \N__24602\,
            I => \N__24599\
        );

    \I__4863\ : LocalMux
    port map (
            O => \N__24599\,
            I => \N__24596\
        );

    \I__4862\ : Odrv4
    port map (
            O => \N__24596\,
            I => \b2v_inst9.data_to_sendZ0Z_2\
        );

    \I__4861\ : CEMux
    port map (
            O => \N__24593\,
            I => \N__24587\
        );

    \I__4860\ : CEMux
    port map (
            O => \N__24592\,
            I => \N__24584\
        );

    \I__4859\ : CEMux
    port map (
            O => \N__24591\,
            I => \N__24581\
        );

    \I__4858\ : CEMux
    port map (
            O => \N__24590\,
            I => \N__24578\
        );

    \I__4857\ : LocalMux
    port map (
            O => \N__24587\,
            I => \N__24575\
        );

    \I__4856\ : LocalMux
    port map (
            O => \N__24584\,
            I => \N__24570\
        );

    \I__4855\ : LocalMux
    port map (
            O => \N__24581\,
            I => \N__24570\
        );

    \I__4854\ : LocalMux
    port map (
            O => \N__24578\,
            I => \N__24567\
        );

    \I__4853\ : Odrv4
    port map (
            O => \N__24575\,
            I => \b2v_inst9.un2_n_fsm_state_0_sqmuxa_2_0_i_0\
        );

    \I__4852\ : Odrv4
    port map (
            O => \N__24570\,
            I => \b2v_inst9.un2_n_fsm_state_0_sqmuxa_2_0_i_0\
        );

    \I__4851\ : Odrv4
    port map (
            O => \N__24567\,
            I => \b2v_inst9.un2_n_fsm_state_0_sqmuxa_2_0_i_0\
        );

    \I__4850\ : InMux
    port map (
            O => \N__24560\,
            I => \N__24551\
        );

    \I__4849\ : InMux
    port map (
            O => \N__24559\,
            I => \N__24551\
        );

    \I__4848\ : InMux
    port map (
            O => \N__24558\,
            I => \N__24551\
        );

    \I__4847\ : LocalMux
    port map (
            O => \N__24551\,
            I => \N__24545\
        );

    \I__4846\ : InMux
    port map (
            O => \N__24550\,
            I => \N__24540\
        );

    \I__4845\ : InMux
    port map (
            O => \N__24549\,
            I => \N__24540\
        );

    \I__4844\ : InMux
    port map (
            O => \N__24548\,
            I => \N__24537\
        );

    \I__4843\ : Odrv12
    port map (
            O => \N__24545\,
            I => \b2v_inst9.N_740\
        );

    \I__4842\ : LocalMux
    port map (
            O => \N__24540\,
            I => \b2v_inst9.N_740\
        );

    \I__4841\ : LocalMux
    port map (
            O => \N__24537\,
            I => \b2v_inst9.N_740\
        );

    \I__4840\ : InMux
    port map (
            O => \N__24530\,
            I => \N__24527\
        );

    \I__4839\ : LocalMux
    port map (
            O => \N__24527\,
            I => \b2v_inst9.data_to_send_10_0_0_1_2\
        );

    \I__4838\ : InMux
    port map (
            O => \N__24524\,
            I => \N__24516\
        );

    \I__4837\ : InMux
    port map (
            O => \N__24523\,
            I => \N__24516\
        );

    \I__4836\ : InMux
    port map (
            O => \N__24522\,
            I => \N__24508\
        );

    \I__4835\ : InMux
    port map (
            O => \N__24521\,
            I => \N__24508\
        );

    \I__4834\ : LocalMux
    port map (
            O => \N__24516\,
            I => \N__24505\
        );

    \I__4833\ : InMux
    port map (
            O => \N__24515\,
            I => \N__24500\
        );

    \I__4832\ : InMux
    port map (
            O => \N__24514\,
            I => \N__24500\
        );

    \I__4831\ : InMux
    port map (
            O => \N__24513\,
            I => \N__24497\
        );

    \I__4830\ : LocalMux
    port map (
            O => \N__24508\,
            I => \b2v_inst9.N_738\
        );

    \I__4829\ : Odrv4
    port map (
            O => \N__24505\,
            I => \b2v_inst9.N_738\
        );

    \I__4828\ : LocalMux
    port map (
            O => \N__24500\,
            I => \b2v_inst9.N_738\
        );

    \I__4827\ : LocalMux
    port map (
            O => \N__24497\,
            I => \b2v_inst9.N_738\
        );

    \I__4826\ : CascadeMux
    port map (
            O => \N__24488\,
            I => \N__24484\
        );

    \I__4825\ : InMux
    port map (
            O => \N__24487\,
            I => \N__24481\
        );

    \I__4824\ : InMux
    port map (
            O => \N__24484\,
            I => \N__24478\
        );

    \I__4823\ : LocalMux
    port map (
            O => \N__24481\,
            I => \N__24470\
        );

    \I__4822\ : LocalMux
    port map (
            O => \N__24478\,
            I => \N__24470\
        );

    \I__4821\ : CascadeMux
    port map (
            O => \N__24477\,
            I => \N__24467\
        );

    \I__4820\ : CascadeMux
    port map (
            O => \N__24476\,
            I => \N__24463\
        );

    \I__4819\ : CascadeMux
    port map (
            O => \N__24475\,
            I => \N__24460\
        );

    \I__4818\ : Span4Mux_h
    port map (
            O => \N__24470\,
            I => \N__24457\
        );

    \I__4817\ : InMux
    port map (
            O => \N__24467\,
            I => \N__24452\
        );

    \I__4816\ : InMux
    port map (
            O => \N__24466\,
            I => \N__24452\
        );

    \I__4815\ : InMux
    port map (
            O => \N__24463\,
            I => \N__24449\
        );

    \I__4814\ : InMux
    port map (
            O => \N__24460\,
            I => \N__24446\
        );

    \I__4813\ : Odrv4
    port map (
            O => \N__24457\,
            I => \b2v_inst9.N_741\
        );

    \I__4812\ : LocalMux
    port map (
            O => \N__24452\,
            I => \b2v_inst9.N_741\
        );

    \I__4811\ : LocalMux
    port map (
            O => \N__24449\,
            I => \b2v_inst9.N_741\
        );

    \I__4810\ : LocalMux
    port map (
            O => \N__24446\,
            I => \b2v_inst9.N_741\
        );

    \I__4809\ : InMux
    port map (
            O => \N__24437\,
            I => \N__24434\
        );

    \I__4808\ : LocalMux
    port map (
            O => \N__24434\,
            I => \N__24431\
        );

    \I__4807\ : Span4Mux_h
    port map (
            O => \N__24431\,
            I => \N__24428\
        );

    \I__4806\ : Odrv4
    port map (
            O => \N__24428\,
            I => \b2v_inst9.data_to_send_10_0_0_1_3\
        );

    \I__4805\ : InMux
    port map (
            O => \N__24425\,
            I => \N__24422\
        );

    \I__4804\ : LocalMux
    port map (
            O => \N__24422\,
            I => \N__24418\
        );

    \I__4803\ : CascadeMux
    port map (
            O => \N__24421\,
            I => \N__24415\
        );

    \I__4802\ : Span4Mux_h
    port map (
            O => \N__24418\,
            I => \N__24412\
        );

    \I__4801\ : InMux
    port map (
            O => \N__24415\,
            I => \N__24409\
        );

    \I__4800\ : Odrv4
    port map (
            O => \N__24412\,
            I => b2v_inst_energia_temp_0
        );

    \I__4799\ : LocalMux
    port map (
            O => \N__24409\,
            I => b2v_inst_energia_temp_0
        );

    \I__4798\ : InMux
    port map (
            O => \N__24404\,
            I => \N__24401\
        );

    \I__4797\ : LocalMux
    port map (
            O => \N__24401\,
            I => \N__24398\
        );

    \I__4796\ : Span4Mux_h
    port map (
            O => \N__24398\,
            I => \N__24395\
        );

    \I__4795\ : Span4Mux_v
    port map (
            O => \N__24395\,
            I => \N__24392\
        );

    \I__4794\ : Odrv4
    port map (
            O => \N__24392\,
            I => \b2v_inst.un14_data_ram_energia_o_axb_0\
        );

    \I__4793\ : InMux
    port map (
            O => \N__24389\,
            I => \N__24385\
        );

    \I__4792\ : CascadeMux
    port map (
            O => \N__24388\,
            I => \N__24382\
        );

    \I__4791\ : LocalMux
    port map (
            O => \N__24385\,
            I => \N__24379\
        );

    \I__4790\ : InMux
    port map (
            O => \N__24382\,
            I => \N__24376\
        );

    \I__4789\ : Odrv4
    port map (
            O => \N__24379\,
            I => b2v_inst_energia_temp_1
        );

    \I__4788\ : LocalMux
    port map (
            O => \N__24376\,
            I => b2v_inst_energia_temp_1
        );

    \I__4787\ : InMux
    port map (
            O => \N__24371\,
            I => \N__24368\
        );

    \I__4786\ : LocalMux
    port map (
            O => \N__24368\,
            I => \N__24365\
        );

    \I__4785\ : Span4Mux_v
    port map (
            O => \N__24365\,
            I => \N__24362\
        );

    \I__4784\ : Span4Mux_v
    port map (
            O => \N__24362\,
            I => \N__24359\
        );

    \I__4783\ : Odrv4
    port map (
            O => \N__24359\,
            I => \b2v_inst.un14_data_ram_energia_o_cry_0_c_RNIEI4MZ0\
        );

    \I__4782\ : InMux
    port map (
            O => \N__24356\,
            I => \b2v_inst.un14_data_ram_energia_o_cry_0\
        );

    \I__4781\ : InMux
    port map (
            O => \N__24353\,
            I => \N__24350\
        );

    \I__4780\ : LocalMux
    port map (
            O => \N__24350\,
            I => \b2v_inst9.data_to_send_10_0_0_0_6\
        );

    \I__4779\ : CascadeMux
    port map (
            O => \N__24347\,
            I => \b2v_inst9.data_to_send_10_0_0_0_7_cascade_\
        );

    \I__4778\ : CascadeMux
    port map (
            O => \N__24344\,
            I => \N__24340\
        );

    \I__4777\ : InMux
    port map (
            O => \N__24343\,
            I => \N__24335\
        );

    \I__4776\ : InMux
    port map (
            O => \N__24340\,
            I => \N__24335\
        );

    \I__4775\ : LocalMux
    port map (
            O => \N__24335\,
            I => \b2v_inst9.data_to_sendZ0Z_7\
        );

    \I__4774\ : InMux
    port map (
            O => \N__24332\,
            I => \N__24329\
        );

    \I__4773\ : LocalMux
    port map (
            O => \N__24329\,
            I => \b2v_inst9.data_to_send_10_0_0_2_0\
        );

    \I__4772\ : InMux
    port map (
            O => \N__24326\,
            I => \N__24323\
        );

    \I__4771\ : LocalMux
    port map (
            O => \N__24323\,
            I => \N__24320\
        );

    \I__4770\ : Span4Mux_v
    port map (
            O => \N__24320\,
            I => \N__24317\
        );

    \I__4769\ : Odrv4
    port map (
            O => \N__24317\,
            I => \b2v_inst9.data_to_send_10_0_0_1_0\
        );

    \I__4768\ : CascadeMux
    port map (
            O => \N__24314\,
            I => \b2v_inst9.N_738_cascade_\
        );

    \I__4767\ : InMux
    port map (
            O => \N__24311\,
            I => \N__24308\
        );

    \I__4766\ : LocalMux
    port map (
            O => \N__24308\,
            I => \N__24305\
        );

    \I__4765\ : Odrv4
    port map (
            O => \N__24305\,
            I => \b2v_inst9.data_to_send_10_0_0_2_1\
        );

    \I__4764\ : InMux
    port map (
            O => \N__24302\,
            I => \N__24299\
        );

    \I__4763\ : LocalMux
    port map (
            O => \N__24299\,
            I => \N__24296\
        );

    \I__4762\ : Span4Mux_v
    port map (
            O => \N__24296\,
            I => \N__24293\
        );

    \I__4761\ : Odrv4
    port map (
            O => \N__24293\,
            I => \b2v_inst9.data_to_sendZ0Z_1\
        );

    \I__4760\ : CascadeMux
    port map (
            O => \N__24290\,
            I => \N_478_cascade_\
        );

    \I__4759\ : InMux
    port map (
            O => \N__24287\,
            I => \N__24284\
        );

    \I__4758\ : LocalMux
    port map (
            O => \N__24284\,
            I => \b2v_inst9.data_to_send_10_0_0_0_0\
        );

    \I__4757\ : InMux
    port map (
            O => \N__24281\,
            I => \N__24277\
        );

    \I__4756\ : InMux
    port map (
            O => \N__24280\,
            I => \N__24270\
        );

    \I__4755\ : LocalMux
    port map (
            O => \N__24277\,
            I => \N__24267\
        );

    \I__4754\ : InMux
    port map (
            O => \N__24276\,
            I => \N__24258\
        );

    \I__4753\ : InMux
    port map (
            O => \N__24275\,
            I => \N__24258\
        );

    \I__4752\ : InMux
    port map (
            O => \N__24274\,
            I => \N__24258\
        );

    \I__4751\ : InMux
    port map (
            O => \N__24273\,
            I => \N__24258\
        );

    \I__4750\ : LocalMux
    port map (
            O => \N__24270\,
            I => \N__24251\
        );

    \I__4749\ : Span4Mux_h
    port map (
            O => \N__24267\,
            I => \N__24246\
        );

    \I__4748\ : LocalMux
    port map (
            O => \N__24258\,
            I => \N__24246\
        );

    \I__4747\ : InMux
    port map (
            O => \N__24257\,
            I => \N__24237\
        );

    \I__4746\ : InMux
    port map (
            O => \N__24256\,
            I => \N__24237\
        );

    \I__4745\ : InMux
    port map (
            O => \N__24255\,
            I => \N__24237\
        );

    \I__4744\ : InMux
    port map (
            O => \N__24254\,
            I => \N__24237\
        );

    \I__4743\ : Odrv4
    port map (
            O => \N__24251\,
            I => \b2v_inst.N_655\
        );

    \I__4742\ : Odrv4
    port map (
            O => \N__24246\,
            I => \b2v_inst.N_655\
        );

    \I__4741\ : LocalMux
    port map (
            O => \N__24237\,
            I => \b2v_inst.N_655\
        );

    \I__4740\ : InMux
    port map (
            O => \N__24230\,
            I => \N__24227\
        );

    \I__4739\ : LocalMux
    port map (
            O => \N__24227\,
            I => \N__24223\
        );

    \I__4738\ : CascadeMux
    port map (
            O => \N__24226\,
            I => \N__24220\
        );

    \I__4737\ : Span4Mux_h
    port map (
            O => \N__24223\,
            I => \N__24217\
        );

    \I__4736\ : InMux
    port map (
            O => \N__24220\,
            I => \N__24214\
        );

    \I__4735\ : Odrv4
    port map (
            O => \N__24217\,
            I => \b2v_inst.un4_cuenta_cry_4_c_RNIFZ0Z888\
        );

    \I__4734\ : LocalMux
    port map (
            O => \N__24214\,
            I => \b2v_inst.un4_cuenta_cry_4_c_RNIFZ0Z888\
        );

    \I__4733\ : CascadeMux
    port map (
            O => \N__24209\,
            I => \N__24206\
        );

    \I__4732\ : InMux
    port map (
            O => \N__24206\,
            I => \N__24202\
        );

    \I__4731\ : InMux
    port map (
            O => \N__24205\,
            I => \N__24199\
        );

    \I__4730\ : LocalMux
    port map (
            O => \N__24202\,
            I => \N__24196\
        );

    \I__4729\ : LocalMux
    port map (
            O => \N__24199\,
            I => \N__24193\
        );

    \I__4728\ : Span4Mux_h
    port map (
            O => \N__24196\,
            I => \N__24188\
        );

    \I__4727\ : Span4Mux_v
    port map (
            O => \N__24193\,
            I => \N__24188\
        );

    \I__4726\ : Odrv4
    port map (
            O => \N__24188\,
            I => \b2v_inst.cuentaZ0Z_5\
        );

    \I__4725\ : CEMux
    port map (
            O => \N__24185\,
            I => \N__24182\
        );

    \I__4724\ : LocalMux
    port map (
            O => \N__24182\,
            I => \N__24176\
        );

    \I__4723\ : CEMux
    port map (
            O => \N__24181\,
            I => \N__24173\
        );

    \I__4722\ : CEMux
    port map (
            O => \N__24180\,
            I => \N__24170\
        );

    \I__4721\ : CEMux
    port map (
            O => \N__24179\,
            I => \N__24167\
        );

    \I__4720\ : Span4Mux_v
    port map (
            O => \N__24176\,
            I => \N__24162\
        );

    \I__4719\ : LocalMux
    port map (
            O => \N__24173\,
            I => \N__24162\
        );

    \I__4718\ : LocalMux
    port map (
            O => \N__24170\,
            I => \N__24159\
        );

    \I__4717\ : LocalMux
    port map (
            O => \N__24167\,
            I => \N__24156\
        );

    \I__4716\ : Span4Mux_v
    port map (
            O => \N__24162\,
            I => \N__24153\
        );

    \I__4715\ : Span4Mux_v
    port map (
            O => \N__24159\,
            I => \N__24150\
        );

    \I__4714\ : Span4Mux_h
    port map (
            O => \N__24156\,
            I => \N__24147\
        );

    \I__4713\ : Span4Mux_h
    port map (
            O => \N__24153\,
            I => \N__24144\
        );

    \I__4712\ : Odrv4
    port map (
            O => \N__24150\,
            I => \b2v_inst.N_547_i_0\
        );

    \I__4711\ : Odrv4
    port map (
            O => \N__24147\,
            I => \b2v_inst.N_547_i_0\
        );

    \I__4710\ : Odrv4
    port map (
            O => \N__24144\,
            I => \b2v_inst.N_547_i_0\
        );

    \I__4709\ : InMux
    port map (
            O => \N__24137\,
            I => \N__24134\
        );

    \I__4708\ : LocalMux
    port map (
            O => \N__24134\,
            I => \N__24131\
        );

    \I__4707\ : Odrv4
    port map (
            O => \N__24131\,
            I => \b2v_inst9.data_to_send_10_0_0_0_4\
        );

    \I__4706\ : CascadeMux
    port map (
            O => \N__24128\,
            I => \N__24125\
        );

    \I__4705\ : InMux
    port map (
            O => \N__24125\,
            I => \N__24122\
        );

    \I__4704\ : LocalMux
    port map (
            O => \N__24122\,
            I => \b2v_inst9.data_to_sendZ0Z_4\
        );

    \I__4703\ : InMux
    port map (
            O => \N__24119\,
            I => \N__24116\
        );

    \I__4702\ : LocalMux
    port map (
            O => \N__24116\,
            I => \b2v_inst9.data_to_send_10_0_0_1_4\
        );

    \I__4701\ : InMux
    port map (
            O => \N__24113\,
            I => \N__24110\
        );

    \I__4700\ : LocalMux
    port map (
            O => \N__24110\,
            I => \N__24107\
        );

    \I__4699\ : Odrv4
    port map (
            O => \N__24107\,
            I => \b2v_inst9.data_to_send_10_0_0_1_5\
        );

    \I__4698\ : InMux
    port map (
            O => \N__24104\,
            I => \N__24101\
        );

    \I__4697\ : LocalMux
    port map (
            O => \N__24101\,
            I => \N__24098\
        );

    \I__4696\ : Span4Mux_h
    port map (
            O => \N__24098\,
            I => \N__24095\
        );

    \I__4695\ : Odrv4
    port map (
            O => \N__24095\,
            I => \b2v_inst9.fsm_state_ns_i_i_0_a2_2_2Z0Z_0\
        );

    \I__4694\ : CascadeMux
    port map (
            O => \N__24092\,
            I => \b2v_inst9.N_583_cascade_\
        );

    \I__4693\ : InMux
    port map (
            O => \N__24089\,
            I => \N__24085\
        );

    \I__4692\ : IoInMux
    port map (
            O => \N__24088\,
            I => \N__24082\
        );

    \I__4691\ : LocalMux
    port map (
            O => \N__24085\,
            I => \N__24079\
        );

    \I__4690\ : LocalMux
    port map (
            O => \N__24082\,
            I => \N__24076\
        );

    \I__4689\ : Span12Mux_v
    port map (
            O => \N__24079\,
            I => \N__24073\
        );

    \I__4688\ : Span4Mux_s3_h
    port map (
            O => \N__24076\,
            I => \N__24070\
        );

    \I__4687\ : Span12Mux_h
    port map (
            O => \N__24073\,
            I => \N__24067\
        );

    \I__4686\ : Span4Mux_v
    port map (
            O => \N__24070\,
            I => \N__24064\
        );

    \I__4685\ : Odrv12
    port map (
            O => \N__24067\,
            I => reset_c_i
        );

    \I__4684\ : Odrv4
    port map (
            O => \N__24064\,
            I => reset_c_i
        );

    \I__4683\ : CascadeMux
    port map (
            O => \N__24059\,
            I => \b2v_inst9.un2_n_fsm_state_0_sqmuxa_2_0_i_cascade_\
        );

    \I__4682\ : InMux
    port map (
            O => \N__24056\,
            I => \N__24053\
        );

    \I__4681\ : LocalMux
    port map (
            O => \N__24053\,
            I => \N__24050\
        );

    \I__4680\ : Span4Mux_h
    port map (
            O => \N__24050\,
            I => \N__24047\
        );

    \I__4679\ : Odrv4
    port map (
            O => \N__24047\,
            I => \b2v_inst.dir_energia_s_6\
        );

    \I__4678\ : InMux
    port map (
            O => \N__24044\,
            I => \b2v_inst.dir_energia_cry_5\
        );

    \I__4677\ : InMux
    port map (
            O => \N__24041\,
            I => \N__24038\
        );

    \I__4676\ : LocalMux
    port map (
            O => \N__24038\,
            I => \N__24035\
        );

    \I__4675\ : Span4Mux_h
    port map (
            O => \N__24035\,
            I => \N__24032\
        );

    \I__4674\ : Odrv4
    port map (
            O => \N__24032\,
            I => \b2v_inst.dir_energia_s_7\
        );

    \I__4673\ : InMux
    port map (
            O => \N__24029\,
            I => \b2v_inst.dir_energia_cry_6\
        );

    \I__4672\ : InMux
    port map (
            O => \N__24026\,
            I => \N__24023\
        );

    \I__4671\ : LocalMux
    port map (
            O => \N__24023\,
            I => \N__24020\
        );

    \I__4670\ : Span4Mux_h
    port map (
            O => \N__24020\,
            I => \N__24017\
        );

    \I__4669\ : Odrv4
    port map (
            O => \N__24017\,
            I => \b2v_inst.dir_energia_s_8\
        );

    \I__4668\ : InMux
    port map (
            O => \N__24014\,
            I => \bfn_13_17_0_\
        );

    \I__4667\ : InMux
    port map (
            O => \N__24011\,
            I => \N__24008\
        );

    \I__4666\ : LocalMux
    port map (
            O => \N__24008\,
            I => \N__24005\
        );

    \I__4665\ : Span4Mux_h
    port map (
            O => \N__24005\,
            I => \N__24002\
        );

    \I__4664\ : Odrv4
    port map (
            O => \N__24002\,
            I => \b2v_inst.dir_energia_s_9\
        );

    \I__4663\ : InMux
    port map (
            O => \N__23999\,
            I => \b2v_inst.dir_energia_cry_8\
        );

    \I__4662\ : InMux
    port map (
            O => \N__23996\,
            I => \N__23993\
        );

    \I__4661\ : LocalMux
    port map (
            O => \N__23993\,
            I => \N__23990\
        );

    \I__4660\ : Span4Mux_v
    port map (
            O => \N__23990\,
            I => \N__23987\
        );

    \I__4659\ : Span4Mux_h
    port map (
            O => \N__23987\,
            I => \N__23984\
        );

    \I__4658\ : Odrv4
    port map (
            O => \N__23984\,
            I => \b2v_inst.dir_energia_s_10\
        );

    \I__4657\ : InMux
    port map (
            O => \N__23981\,
            I => \b2v_inst.dir_energia_cry_9\
        );

    \I__4656\ : InMux
    port map (
            O => \N__23978\,
            I => \N__23973\
        );

    \I__4655\ : CascadeMux
    port map (
            O => \N__23977\,
            I => \N__23970\
        );

    \I__4654\ : CascadeMux
    port map (
            O => \N__23976\,
            I => \N__23963\
        );

    \I__4653\ : LocalMux
    port map (
            O => \N__23973\,
            I => \N__23960\
        );

    \I__4652\ : InMux
    port map (
            O => \N__23970\,
            I => \N__23951\
        );

    \I__4651\ : InMux
    port map (
            O => \N__23969\,
            I => \N__23951\
        );

    \I__4650\ : InMux
    port map (
            O => \N__23968\,
            I => \N__23951\
        );

    \I__4649\ : InMux
    port map (
            O => \N__23967\,
            I => \N__23951\
        );

    \I__4648\ : InMux
    port map (
            O => \N__23966\,
            I => \N__23945\
        );

    \I__4647\ : InMux
    port map (
            O => \N__23963\,
            I => \N__23942\
        );

    \I__4646\ : Span4Mux_v
    port map (
            O => \N__23960\,
            I => \N__23939\
        );

    \I__4645\ : LocalMux
    port map (
            O => \N__23951\,
            I => \N__23936\
        );

    \I__4644\ : InMux
    port map (
            O => \N__23950\,
            I => \N__23929\
        );

    \I__4643\ : InMux
    port map (
            O => \N__23949\,
            I => \N__23929\
        );

    \I__4642\ : InMux
    port map (
            O => \N__23948\,
            I => \N__23929\
        );

    \I__4641\ : LocalMux
    port map (
            O => \N__23945\,
            I => \N__23926\
        );

    \I__4640\ : LocalMux
    port map (
            O => \N__23942\,
            I => \N__23921\
        );

    \I__4639\ : Span4Mux_h
    port map (
            O => \N__23939\,
            I => \N__23921\
        );

    \I__4638\ : Span4Mux_v
    port map (
            O => \N__23936\,
            I => \N__23916\
        );

    \I__4637\ : LocalMux
    port map (
            O => \N__23929\,
            I => \N__23916\
        );

    \I__4636\ : Span4Mux_v
    port map (
            O => \N__23926\,
            I => \N__23909\
        );

    \I__4635\ : Span4Mux_v
    port map (
            O => \N__23921\,
            I => \N__23904\
        );

    \I__4634\ : Span4Mux_v
    port map (
            O => \N__23916\,
            I => \N__23904\
        );

    \I__4633\ : InMux
    port map (
            O => \N__23915\,
            I => \N__23899\
        );

    \I__4632\ : InMux
    port map (
            O => \N__23914\,
            I => \N__23899\
        );

    \I__4631\ : InMux
    port map (
            O => \N__23913\,
            I => \N__23894\
        );

    \I__4630\ : InMux
    port map (
            O => \N__23912\,
            I => \N__23894\
        );

    \I__4629\ : Sp12to4
    port map (
            O => \N__23909\,
            I => \N__23885\
        );

    \I__4628\ : Sp12to4
    port map (
            O => \N__23904\,
            I => \N__23885\
        );

    \I__4627\ : LocalMux
    port map (
            O => \N__23899\,
            I => \N__23885\
        );

    \I__4626\ : LocalMux
    port map (
            O => \N__23894\,
            I => \N__23885\
        );

    \I__4625\ : Odrv12
    port map (
            O => \N__23885\,
            I => \b2v_inst.stateZ0Z_19\
        );

    \I__4624\ : CascadeMux
    port map (
            O => \N__23882\,
            I => \N__23879\
        );

    \I__4623\ : InMux
    port map (
            O => \N__23879\,
            I => \N__23876\
        );

    \I__4622\ : LocalMux
    port map (
            O => \N__23876\,
            I => \N__23862\
        );

    \I__4621\ : InMux
    port map (
            O => \N__23875\,
            I => \N__23847\
        );

    \I__4620\ : InMux
    port map (
            O => \N__23874\,
            I => \N__23847\
        );

    \I__4619\ : InMux
    port map (
            O => \N__23873\,
            I => \N__23847\
        );

    \I__4618\ : InMux
    port map (
            O => \N__23872\,
            I => \N__23847\
        );

    \I__4617\ : InMux
    port map (
            O => \N__23871\,
            I => \N__23847\
        );

    \I__4616\ : InMux
    port map (
            O => \N__23870\,
            I => \N__23847\
        );

    \I__4615\ : InMux
    port map (
            O => \N__23869\,
            I => \N__23847\
        );

    \I__4614\ : InMux
    port map (
            O => \N__23868\,
            I => \N__23838\
        );

    \I__4613\ : InMux
    port map (
            O => \N__23867\,
            I => \N__23838\
        );

    \I__4612\ : InMux
    port map (
            O => \N__23866\,
            I => \N__23838\
        );

    \I__4611\ : InMux
    port map (
            O => \N__23865\,
            I => \N__23838\
        );

    \I__4610\ : Span4Mux_v
    port map (
            O => \N__23862\,
            I => \N__23835\
        );

    \I__4609\ : LocalMux
    port map (
            O => \N__23847\,
            I => \b2v_inst.N_352_0\
        );

    \I__4608\ : LocalMux
    port map (
            O => \N__23838\,
            I => \b2v_inst.N_352_0\
        );

    \I__4607\ : Odrv4
    port map (
            O => \N__23835\,
            I => \b2v_inst.N_352_0\
        );

    \I__4606\ : InMux
    port map (
            O => \N__23828\,
            I => \b2v_inst.dir_energia_cry_10\
        );

    \I__4605\ : CascadeMux
    port map (
            O => \N__23825\,
            I => \N__23822\
        );

    \I__4604\ : InMux
    port map (
            O => \N__23822\,
            I => \N__23819\
        );

    \I__4603\ : LocalMux
    port map (
            O => \N__23819\,
            I => \N__23815\
        );

    \I__4602\ : InMux
    port map (
            O => \N__23818\,
            I => \N__23812\
        );

    \I__4601\ : Span4Mux_h
    port map (
            O => \N__23815\,
            I => \N__23809\
        );

    \I__4600\ : LocalMux
    port map (
            O => \N__23812\,
            I => \b2v_inst.dir_energiaZ0Z_11\
        );

    \I__4599\ : Odrv4
    port map (
            O => \N__23809\,
            I => \b2v_inst.dir_energiaZ0Z_11\
        );

    \I__4598\ : CEMux
    port map (
            O => \N__23804\,
            I => \N__23801\
        );

    \I__4597\ : LocalMux
    port map (
            O => \N__23801\,
            I => \N__23796\
        );

    \I__4596\ : CEMux
    port map (
            O => \N__23800\,
            I => \N__23793\
        );

    \I__4595\ : CEMux
    port map (
            O => \N__23799\,
            I => \N__23790\
        );

    \I__4594\ : Span4Mux_v
    port map (
            O => \N__23796\,
            I => \N__23785\
        );

    \I__4593\ : LocalMux
    port map (
            O => \N__23793\,
            I => \N__23785\
        );

    \I__4592\ : LocalMux
    port map (
            O => \N__23790\,
            I => \N__23782\
        );

    \I__4591\ : Span4Mux_h
    port map (
            O => \N__23785\,
            I => \N__23779\
        );

    \I__4590\ : Odrv4
    port map (
            O => \N__23782\,
            I => \b2v_inst.N_430_i\
        );

    \I__4589\ : Odrv4
    port map (
            O => \N__23779\,
            I => \b2v_inst.N_430_i\
        );

    \I__4588\ : InMux
    port map (
            O => \N__23774\,
            I => \N__23771\
        );

    \I__4587\ : LocalMux
    port map (
            O => \N__23771\,
            I => \N__23768\
        );

    \I__4586\ : Odrv4
    port map (
            O => \N__23768\,
            I => \b2v_inst.N_648_5\
        );

    \I__4585\ : InMux
    port map (
            O => \N__23765\,
            I => \N__23756\
        );

    \I__4584\ : InMux
    port map (
            O => \N__23764\,
            I => \N__23756\
        );

    \I__4583\ : InMux
    port map (
            O => \N__23763\,
            I => \N__23756\
        );

    \I__4582\ : LocalMux
    port map (
            O => \N__23756\,
            I => \N__23753\
        );

    \I__4581\ : Span4Mux_h
    port map (
            O => \N__23753\,
            I => \N__23750\
        );

    \I__4580\ : Span4Mux_v
    port map (
            O => \N__23750\,
            I => \N__23745\
        );

    \I__4579\ : InMux
    port map (
            O => \N__23749\,
            I => \N__23742\
        );

    \I__4578\ : InMux
    port map (
            O => \N__23748\,
            I => \N__23739\
        );

    \I__4577\ : Span4Mux_v
    port map (
            O => \N__23745\,
            I => \N__23736\
        );

    \I__4576\ : LocalMux
    port map (
            O => \N__23742\,
            I => \N__23733\
        );

    \I__4575\ : LocalMux
    port map (
            O => \N__23739\,
            I => \b2v_inst.un9_indice_0_a2_5_1\
        );

    \I__4574\ : Odrv4
    port map (
            O => \N__23736\,
            I => \b2v_inst.un9_indice_0_a2_5_1\
        );

    \I__4573\ : Odrv4
    port map (
            O => \N__23733\,
            I => \b2v_inst.un9_indice_0_a2_5_1\
        );

    \I__4572\ : InMux
    port map (
            O => \N__23726\,
            I => \N__23723\
        );

    \I__4571\ : LocalMux
    port map (
            O => \N__23723\,
            I => \N__23720\
        );

    \I__4570\ : Span4Mux_v
    port map (
            O => \N__23720\,
            I => \N__23715\
        );

    \I__4569\ : InMux
    port map (
            O => \N__23719\,
            I => \N__23710\
        );

    \I__4568\ : InMux
    port map (
            O => \N__23718\,
            I => \N__23710\
        );

    \I__4567\ : Odrv4
    port map (
            O => \N__23715\,
            I => \b2v_inst.un4_cuenta_cry_9_c_RNI01TZ0Z9\
        );

    \I__4566\ : LocalMux
    port map (
            O => \N__23710\,
            I => \b2v_inst.un4_cuenta_cry_9_c_RNI01TZ0Z9\
        );

    \I__4565\ : InMux
    port map (
            O => \N__23705\,
            I => \N__23701\
        );

    \I__4564\ : CascadeMux
    port map (
            O => \N__23704\,
            I => \N__23698\
        );

    \I__4563\ : LocalMux
    port map (
            O => \N__23701\,
            I => \N__23695\
        );

    \I__4562\ : InMux
    port map (
            O => \N__23698\,
            I => \N__23692\
        );

    \I__4561\ : Span4Mux_v
    port map (
            O => \N__23695\,
            I => \N__23687\
        );

    \I__4560\ : LocalMux
    port map (
            O => \N__23692\,
            I => \N__23687\
        );

    \I__4559\ : Span4Mux_v
    port map (
            O => \N__23687\,
            I => \N__23684\
        );

    \I__4558\ : Odrv4
    port map (
            O => \N__23684\,
            I => \b2v_inst.cuentaZ0Z_10\
        );

    \I__4557\ : InMux
    port map (
            O => \N__23681\,
            I => \N__23678\
        );

    \I__4556\ : LocalMux
    port map (
            O => \N__23678\,
            I => \N__23675\
        );

    \I__4555\ : Span4Mux_h
    port map (
            O => \N__23675\,
            I => \N__23671\
        );

    \I__4554\ : IoInMux
    port map (
            O => \N__23674\,
            I => \N__23668\
        );

    \I__4553\ : Span4Mux_v
    port map (
            O => \N__23671\,
            I => \N__23665\
        );

    \I__4552\ : LocalMux
    port map (
            O => \N__23668\,
            I => \N__23662\
        );

    \I__4551\ : Span4Mux_h
    port map (
            O => \N__23665\,
            I => \N__23659\
        );

    \I__4550\ : Odrv12
    port map (
            O => \N__23662\,
            I => leds_c_2
        );

    \I__4549\ : Odrv4
    port map (
            O => \N__23659\,
            I => leds_c_2
        );

    \I__4548\ : InMux
    port map (
            O => \N__23654\,
            I => \N__23650\
        );

    \I__4547\ : IoInMux
    port map (
            O => \N__23653\,
            I => \N__23647\
        );

    \I__4546\ : LocalMux
    port map (
            O => \N__23650\,
            I => \N__23644\
        );

    \I__4545\ : LocalMux
    port map (
            O => \N__23647\,
            I => \N__23641\
        );

    \I__4544\ : Span4Mux_v
    port map (
            O => \N__23644\,
            I => \N__23638\
        );

    \I__4543\ : Span4Mux_s3_h
    port map (
            O => \N__23641\,
            I => \N__23635\
        );

    \I__4542\ : Span4Mux_h
    port map (
            O => \N__23638\,
            I => \N__23632\
        );

    \I__4541\ : Span4Mux_h
    port map (
            O => \N__23635\,
            I => \N__23629\
        );

    \I__4540\ : Span4Mux_h
    port map (
            O => \N__23632\,
            I => \N__23626\
        );

    \I__4539\ : Odrv4
    port map (
            O => \N__23629\,
            I => leds_c_3
        );

    \I__4538\ : Odrv4
    port map (
            O => \N__23626\,
            I => leds_c_3
        );

    \I__4537\ : InMux
    port map (
            O => \N__23621\,
            I => \N__23618\
        );

    \I__4536\ : LocalMux
    port map (
            O => \N__23618\,
            I => \N__23615\
        );

    \I__4535\ : Span4Mux_h
    port map (
            O => \N__23615\,
            I => \N__23612\
        );

    \I__4534\ : Span4Mux_h
    port map (
            O => \N__23612\,
            I => \N__23609\
        );

    \I__4533\ : Span4Mux_h
    port map (
            O => \N__23609\,
            I => \N__23606\
        );

    \I__4532\ : Odrv4
    port map (
            O => \N__23606\,
            I => \N_546_i\
        );

    \I__4531\ : InMux
    port map (
            O => \N__23603\,
            I => \N__23600\
        );

    \I__4530\ : LocalMux
    port map (
            O => \N__23600\,
            I => \N__23597\
        );

    \I__4529\ : Span4Mux_h
    port map (
            O => \N__23597\,
            I => \N__23594\
        );

    \I__4528\ : Odrv4
    port map (
            O => \N__23594\,
            I => \b2v_inst.dir_energia_s_1\
        );

    \I__4527\ : InMux
    port map (
            O => \N__23591\,
            I => \b2v_inst.dir_energia_cry_0\
        );

    \I__4526\ : CascadeMux
    port map (
            O => \N__23588\,
            I => \N__23585\
        );

    \I__4525\ : InMux
    port map (
            O => \N__23585\,
            I => \N__23582\
        );

    \I__4524\ : LocalMux
    port map (
            O => \N__23582\,
            I => \N__23579\
        );

    \I__4523\ : Span4Mux_v
    port map (
            O => \N__23579\,
            I => \N__23576\
        );

    \I__4522\ : Odrv4
    port map (
            O => \N__23576\,
            I => \b2v_inst.dir_energia_s_2\
        );

    \I__4521\ : InMux
    port map (
            O => \N__23573\,
            I => \b2v_inst.dir_energia_cry_1\
        );

    \I__4520\ : InMux
    port map (
            O => \N__23570\,
            I => \N__23567\
        );

    \I__4519\ : LocalMux
    port map (
            O => \N__23567\,
            I => \N__23564\
        );

    \I__4518\ : Span4Mux_v
    port map (
            O => \N__23564\,
            I => \N__23561\
        );

    \I__4517\ : Odrv4
    port map (
            O => \N__23561\,
            I => \b2v_inst.dir_energia_s_3\
        );

    \I__4516\ : InMux
    port map (
            O => \N__23558\,
            I => \b2v_inst.dir_energia_cry_2\
        );

    \I__4515\ : CascadeMux
    port map (
            O => \N__23555\,
            I => \N__23552\
        );

    \I__4514\ : InMux
    port map (
            O => \N__23552\,
            I => \N__23549\
        );

    \I__4513\ : LocalMux
    port map (
            O => \N__23549\,
            I => \N__23546\
        );

    \I__4512\ : Span4Mux_v
    port map (
            O => \N__23546\,
            I => \N__23543\
        );

    \I__4511\ : Span4Mux_h
    port map (
            O => \N__23543\,
            I => \N__23540\
        );

    \I__4510\ : Odrv4
    port map (
            O => \N__23540\,
            I => \b2v_inst.dir_energia_s_4\
        );

    \I__4509\ : InMux
    port map (
            O => \N__23537\,
            I => \b2v_inst.dir_energia_cry_3\
        );

    \I__4508\ : InMux
    port map (
            O => \N__23534\,
            I => \N__23531\
        );

    \I__4507\ : LocalMux
    port map (
            O => \N__23531\,
            I => \N__23528\
        );

    \I__4506\ : Span4Mux_h
    port map (
            O => \N__23528\,
            I => \N__23525\
        );

    \I__4505\ : Odrv4
    port map (
            O => \N__23525\,
            I => \b2v_inst.dir_energia_s_5\
        );

    \I__4504\ : InMux
    port map (
            O => \N__23522\,
            I => \b2v_inst.dir_energia_cry_4\
        );

    \I__4503\ : InMux
    port map (
            O => \N__23519\,
            I => \N__23516\
        );

    \I__4502\ : LocalMux
    port map (
            O => \N__23516\,
            I => \N__23513\
        );

    \I__4501\ : Span4Mux_v
    port map (
            O => \N__23513\,
            I => \N__23509\
        );

    \I__4500\ : InMux
    port map (
            O => \N__23512\,
            I => \N__23506\
        );

    \I__4499\ : Odrv4
    port map (
            O => \N__23509\,
            I => \b2v_inst.cuentaZ0Z_9\
        );

    \I__4498\ : LocalMux
    port map (
            O => \N__23506\,
            I => \b2v_inst.cuentaZ0Z_9\
        );

    \I__4497\ : InMux
    port map (
            O => \N__23501\,
            I => \N__23498\
        );

    \I__4496\ : LocalMux
    port map (
            O => \N__23498\,
            I => \N__23493\
        );

    \I__4495\ : InMux
    port map (
            O => \N__23497\,
            I => \N__23488\
        );

    \I__4494\ : InMux
    port map (
            O => \N__23496\,
            I => \N__23488\
        );

    \I__4493\ : Odrv12
    port map (
            O => \N__23493\,
            I => \b2v_inst.un4_cuenta_cry_8_c_RNINKCZ0Z8\
        );

    \I__4492\ : LocalMux
    port map (
            O => \N__23488\,
            I => \b2v_inst.un4_cuenta_cry_8_c_RNINKCZ0Z8\
        );

    \I__4491\ : InMux
    port map (
            O => \N__23483\,
            I => \bfn_13_13_0_\
        );

    \I__4490\ : InMux
    port map (
            O => \N__23480\,
            I => \b2v_inst.un4_cuenta_cry_9\
        );

    \I__4489\ : InMux
    port map (
            O => \N__23477\,
            I => \N__23474\
        );

    \I__4488\ : LocalMux
    port map (
            O => \N__23474\,
            I => \N__23471\
        );

    \I__4487\ : Span4Mux_h
    port map (
            O => \N__23471\,
            I => \N__23468\
        );

    \I__4486\ : Span4Mux_h
    port map (
            O => \N__23468\,
            I => \N__23465\
        );

    \I__4485\ : Odrv4
    port map (
            O => \N__23465\,
            I => \N_458_i\
        );

    \I__4484\ : InMux
    port map (
            O => \N__23462\,
            I => \N__23459\
        );

    \I__4483\ : LocalMux
    port map (
            O => \N__23459\,
            I => \N__23455\
        );

    \I__4482\ : CascadeMux
    port map (
            O => \N__23458\,
            I => \N__23452\
        );

    \I__4481\ : Span4Mux_h
    port map (
            O => \N__23455\,
            I => \N__23447\
        );

    \I__4480\ : InMux
    port map (
            O => \N__23452\,
            I => \N__23440\
        );

    \I__4479\ : InMux
    port map (
            O => \N__23451\,
            I => \N__23440\
        );

    \I__4478\ : InMux
    port map (
            O => \N__23450\,
            I => \N__23440\
        );

    \I__4477\ : Odrv4
    port map (
            O => \N__23447\,
            I => b2v_inst_state_4
        );

    \I__4476\ : LocalMux
    port map (
            O => \N__23440\,
            I => b2v_inst_state_4
        );

    \I__4475\ : InMux
    port map (
            O => \N__23435\,
            I => \N__23432\
        );

    \I__4474\ : LocalMux
    port map (
            O => \N__23432\,
            I => \N__23427\
        );

    \I__4473\ : CascadeMux
    port map (
            O => \N__23431\,
            I => \N__23424\
        );

    \I__4472\ : CascadeMux
    port map (
            O => \N__23430\,
            I => \N__23420\
        );

    \I__4471\ : Span4Mux_v
    port map (
            O => \N__23427\,
            I => \N__23417\
        );

    \I__4470\ : InMux
    port map (
            O => \N__23424\,
            I => \N__23410\
        );

    \I__4469\ : InMux
    port map (
            O => \N__23423\,
            I => \N__23410\
        );

    \I__4468\ : InMux
    port map (
            O => \N__23420\,
            I => \N__23410\
        );

    \I__4467\ : Odrv4
    port map (
            O => \N__23417\,
            I => b2v_inst_state_8
        );

    \I__4466\ : LocalMux
    port map (
            O => \N__23410\,
            I => b2v_inst_state_8
        );

    \I__4465\ : InMux
    port map (
            O => \N__23405\,
            I => \N__23401\
        );

    \I__4464\ : IoInMux
    port map (
            O => \N__23404\,
            I => \N__23398\
        );

    \I__4463\ : LocalMux
    port map (
            O => \N__23401\,
            I => \N__23395\
        );

    \I__4462\ : LocalMux
    port map (
            O => \N__23398\,
            I => \N__23392\
        );

    \I__4461\ : Span4Mux_v
    port map (
            O => \N__23395\,
            I => \N__23389\
        );

    \I__4460\ : Span12Mux_s6_v
    port map (
            O => \N__23392\,
            I => \N__23386\
        );

    \I__4459\ : Span4Mux_h
    port map (
            O => \N__23389\,
            I => \N__23383\
        );

    \I__4458\ : Span12Mux_v
    port map (
            O => \N__23386\,
            I => \N__23380\
        );

    \I__4457\ : Span4Mux_h
    port map (
            O => \N__23383\,
            I => \N__23377\
        );

    \I__4456\ : Odrv12
    port map (
            O => \N__23380\,
            I => leds_c_0
        );

    \I__4455\ : Odrv4
    port map (
            O => \N__23377\,
            I => leds_c_0
        );

    \I__4454\ : IoInMux
    port map (
            O => \N__23372\,
            I => \N__23368\
        );

    \I__4453\ : InMux
    port map (
            O => \N__23371\,
            I => \N__23365\
        );

    \I__4452\ : LocalMux
    port map (
            O => \N__23368\,
            I => \N__23362\
        );

    \I__4451\ : LocalMux
    port map (
            O => \N__23365\,
            I => \N__23359\
        );

    \I__4450\ : Span4Mux_s3_h
    port map (
            O => \N__23362\,
            I => \N__23356\
        );

    \I__4449\ : Span4Mux_h
    port map (
            O => \N__23359\,
            I => \N__23353\
        );

    \I__4448\ : Span4Mux_v
    port map (
            O => \N__23356\,
            I => \N__23350\
        );

    \I__4447\ : Span4Mux_h
    port map (
            O => \N__23353\,
            I => \N__23347\
        );

    \I__4446\ : Span4Mux_v
    port map (
            O => \N__23350\,
            I => \N__23344\
        );

    \I__4445\ : Span4Mux_h
    port map (
            O => \N__23347\,
            I => \N__23341\
        );

    \I__4444\ : Span4Mux_h
    port map (
            O => \N__23344\,
            I => \N__23336\
        );

    \I__4443\ : Span4Mux_v
    port map (
            O => \N__23341\,
            I => \N__23336\
        );

    \I__4442\ : Odrv4
    port map (
            O => \N__23336\,
            I => leds_c_1
        );

    \I__4441\ : InMux
    port map (
            O => \N__23333\,
            I => \N__23329\
        );

    \I__4440\ : IoInMux
    port map (
            O => \N__23332\,
            I => \N__23326\
        );

    \I__4439\ : LocalMux
    port map (
            O => \N__23329\,
            I => \N__23323\
        );

    \I__4438\ : LocalMux
    port map (
            O => \N__23326\,
            I => \N__23320\
        );

    \I__4437\ : Span4Mux_v
    port map (
            O => \N__23323\,
            I => \N__23317\
        );

    \I__4436\ : Span4Mux_s3_h
    port map (
            O => \N__23320\,
            I => \N__23314\
        );

    \I__4435\ : Span4Mux_h
    port map (
            O => \N__23317\,
            I => \N__23311\
        );

    \I__4434\ : Span4Mux_h
    port map (
            O => \N__23314\,
            I => \N__23308\
        );

    \I__4433\ : Span4Mux_h
    port map (
            O => \N__23311\,
            I => \N__23305\
        );

    \I__4432\ : Odrv4
    port map (
            O => \N__23308\,
            I => leds_c_13
        );

    \I__4431\ : Odrv4
    port map (
            O => \N__23305\,
            I => leds_c_13
        );

    \I__4430\ : InMux
    port map (
            O => \N__23300\,
            I => \N__23293\
        );

    \I__4429\ : InMux
    port map (
            O => \N__23299\,
            I => \N__23288\
        );

    \I__4428\ : InMux
    port map (
            O => \N__23298\,
            I => \N__23288\
        );

    \I__4427\ : InMux
    port map (
            O => \N__23297\,
            I => \N__23285\
        );

    \I__4426\ : InMux
    port map (
            O => \N__23296\,
            I => \N__23282\
        );

    \I__4425\ : LocalMux
    port map (
            O => \N__23293\,
            I => \b2v_inst.cuentaZ0Z_0\
        );

    \I__4424\ : LocalMux
    port map (
            O => \N__23288\,
            I => \b2v_inst.cuentaZ0Z_0\
        );

    \I__4423\ : LocalMux
    port map (
            O => \N__23285\,
            I => \b2v_inst.cuentaZ0Z_0\
        );

    \I__4422\ : LocalMux
    port map (
            O => \N__23282\,
            I => \b2v_inst.cuentaZ0Z_0\
        );

    \I__4421\ : InMux
    port map (
            O => \N__23273\,
            I => \N__23269\
        );

    \I__4420\ : CascadeMux
    port map (
            O => \N__23272\,
            I => \N__23265\
        );

    \I__4419\ : LocalMux
    port map (
            O => \N__23269\,
            I => \N__23262\
        );

    \I__4418\ : InMux
    port map (
            O => \N__23268\,
            I => \N__23259\
        );

    \I__4417\ : InMux
    port map (
            O => \N__23265\,
            I => \N__23256\
        );

    \I__4416\ : Odrv4
    port map (
            O => \N__23262\,
            I => \b2v_inst.cuentaZ0Z_1\
        );

    \I__4415\ : LocalMux
    port map (
            O => \N__23259\,
            I => \b2v_inst.cuentaZ0Z_1\
        );

    \I__4414\ : LocalMux
    port map (
            O => \N__23256\,
            I => \b2v_inst.cuentaZ0Z_1\
        );

    \I__4413\ : CascadeMux
    port map (
            O => \N__23249\,
            I => \N__23245\
        );

    \I__4412\ : InMux
    port map (
            O => \N__23248\,
            I => \N__23242\
        );

    \I__4411\ : InMux
    port map (
            O => \N__23245\,
            I => \N__23239\
        );

    \I__4410\ : LocalMux
    port map (
            O => \N__23242\,
            I => \b2v_inst.cuentaZ0Z_2\
        );

    \I__4409\ : LocalMux
    port map (
            O => \N__23239\,
            I => \b2v_inst.cuentaZ0Z_2\
        );

    \I__4408\ : InMux
    port map (
            O => \N__23234\,
            I => \N__23230\
        );

    \I__4407\ : InMux
    port map (
            O => \N__23233\,
            I => \N__23227\
        );

    \I__4406\ : LocalMux
    port map (
            O => \N__23230\,
            I => \N__23224\
        );

    \I__4405\ : LocalMux
    port map (
            O => \N__23227\,
            I => \b2v_inst.un4_cuenta_cry_1_c_RNI9VZ0Z48\
        );

    \I__4404\ : Odrv4
    port map (
            O => \N__23224\,
            I => \b2v_inst.un4_cuenta_cry_1_c_RNI9VZ0Z48\
        );

    \I__4403\ : InMux
    port map (
            O => \N__23219\,
            I => \b2v_inst.un4_cuenta_cry_1\
        );

    \I__4402\ : CascadeMux
    port map (
            O => \N__23216\,
            I => \N__23212\
        );

    \I__4401\ : InMux
    port map (
            O => \N__23215\,
            I => \N__23209\
        );

    \I__4400\ : InMux
    port map (
            O => \N__23212\,
            I => \N__23206\
        );

    \I__4399\ : LocalMux
    port map (
            O => \N__23209\,
            I => \b2v_inst.cuentaZ0Z_3\
        );

    \I__4398\ : LocalMux
    port map (
            O => \N__23206\,
            I => \b2v_inst.cuentaZ0Z_3\
        );

    \I__4397\ : InMux
    port map (
            O => \N__23201\,
            I => \N__23197\
        );

    \I__4396\ : InMux
    port map (
            O => \N__23200\,
            I => \N__23194\
        );

    \I__4395\ : LocalMux
    port map (
            O => \N__23197\,
            I => \b2v_inst.un4_cuenta_cry_2_c_RNIBZ0Z268\
        );

    \I__4394\ : LocalMux
    port map (
            O => \N__23194\,
            I => \b2v_inst.un4_cuenta_cry_2_c_RNIBZ0Z268\
        );

    \I__4393\ : InMux
    port map (
            O => \N__23189\,
            I => \b2v_inst.un4_cuenta_cry_2\
        );

    \I__4392\ : CascadeMux
    port map (
            O => \N__23186\,
            I => \N__23182\
        );

    \I__4391\ : InMux
    port map (
            O => \N__23185\,
            I => \N__23179\
        );

    \I__4390\ : InMux
    port map (
            O => \N__23182\,
            I => \N__23176\
        );

    \I__4389\ : LocalMux
    port map (
            O => \N__23179\,
            I => \b2v_inst.cuentaZ0Z_4\
        );

    \I__4388\ : LocalMux
    port map (
            O => \N__23176\,
            I => \b2v_inst.cuentaZ0Z_4\
        );

    \I__4387\ : InMux
    port map (
            O => \N__23171\,
            I => \N__23167\
        );

    \I__4386\ : InMux
    port map (
            O => \N__23170\,
            I => \N__23164\
        );

    \I__4385\ : LocalMux
    port map (
            O => \N__23167\,
            I => \b2v_inst.un4_cuenta_cry_3_c_RNIDZ0Z578\
        );

    \I__4384\ : LocalMux
    port map (
            O => \N__23164\,
            I => \b2v_inst.un4_cuenta_cry_3_c_RNIDZ0Z578\
        );

    \I__4383\ : InMux
    port map (
            O => \N__23159\,
            I => \b2v_inst.un4_cuenta_cry_3\
        );

    \I__4382\ : InMux
    port map (
            O => \N__23156\,
            I => \b2v_inst.un4_cuenta_cry_4\
        );

    \I__4381\ : InMux
    port map (
            O => \N__23153\,
            I => \N__23149\
        );

    \I__4380\ : InMux
    port map (
            O => \N__23152\,
            I => \N__23146\
        );

    \I__4379\ : LocalMux
    port map (
            O => \N__23149\,
            I => \N__23141\
        );

    \I__4378\ : LocalMux
    port map (
            O => \N__23146\,
            I => \N__23141\
        );

    \I__4377\ : Span4Mux_v
    port map (
            O => \N__23141\,
            I => \N__23138\
        );

    \I__4376\ : Odrv4
    port map (
            O => \N__23138\,
            I => \b2v_inst.cuentaZ0Z_6\
        );

    \I__4375\ : InMux
    port map (
            O => \N__23135\,
            I => \N__23132\
        );

    \I__4374\ : LocalMux
    port map (
            O => \N__23132\,
            I => \N__23128\
        );

    \I__4373\ : InMux
    port map (
            O => \N__23131\,
            I => \N__23125\
        );

    \I__4372\ : Odrv12
    port map (
            O => \N__23128\,
            I => \b2v_inst.un4_cuenta_cry_5_c_RNIHBZ0Z98\
        );

    \I__4371\ : LocalMux
    port map (
            O => \N__23125\,
            I => \b2v_inst.un4_cuenta_cry_5_c_RNIHBZ0Z98\
        );

    \I__4370\ : InMux
    port map (
            O => \N__23120\,
            I => \b2v_inst.un4_cuenta_cry_5\
        );

    \I__4369\ : CascadeMux
    port map (
            O => \N__23117\,
            I => \N__23113\
        );

    \I__4368\ : InMux
    port map (
            O => \N__23116\,
            I => \N__23110\
        );

    \I__4367\ : InMux
    port map (
            O => \N__23113\,
            I => \N__23107\
        );

    \I__4366\ : LocalMux
    port map (
            O => \N__23110\,
            I => \N__23104\
        );

    \I__4365\ : LocalMux
    port map (
            O => \N__23107\,
            I => \N__23099\
        );

    \I__4364\ : Span4Mux_v
    port map (
            O => \N__23104\,
            I => \N__23099\
        );

    \I__4363\ : Odrv4
    port map (
            O => \N__23099\,
            I => \b2v_inst.cuentaZ0Z_7\
        );

    \I__4362\ : InMux
    port map (
            O => \N__23096\,
            I => \N__23093\
        );

    \I__4361\ : LocalMux
    port map (
            O => \N__23093\,
            I => \N__23089\
        );

    \I__4360\ : InMux
    port map (
            O => \N__23092\,
            I => \N__23086\
        );

    \I__4359\ : Odrv12
    port map (
            O => \N__23089\,
            I => \b2v_inst.un4_cuenta_cry_6_c_RNIJEAZ0Z8\
        );

    \I__4358\ : LocalMux
    port map (
            O => \N__23086\,
            I => \b2v_inst.un4_cuenta_cry_6_c_RNIJEAZ0Z8\
        );

    \I__4357\ : InMux
    port map (
            O => \N__23081\,
            I => \b2v_inst.un4_cuenta_cry_6\
        );

    \I__4356\ : InMux
    port map (
            O => \N__23078\,
            I => \N__23075\
        );

    \I__4355\ : LocalMux
    port map (
            O => \N__23075\,
            I => \N__23071\
        );

    \I__4354\ : InMux
    port map (
            O => \N__23074\,
            I => \N__23068\
        );

    \I__4353\ : Span4Mux_v
    port map (
            O => \N__23071\,
            I => \N__23065\
        );

    \I__4352\ : LocalMux
    port map (
            O => \N__23068\,
            I => \b2v_inst.cuentaZ0Z_8\
        );

    \I__4351\ : Odrv4
    port map (
            O => \N__23065\,
            I => \b2v_inst.cuentaZ0Z_8\
        );

    \I__4350\ : InMux
    port map (
            O => \N__23060\,
            I => \N__23057\
        );

    \I__4349\ : LocalMux
    port map (
            O => \N__23057\,
            I => \N__23052\
        );

    \I__4348\ : InMux
    port map (
            O => \N__23056\,
            I => \N__23047\
        );

    \I__4347\ : InMux
    port map (
            O => \N__23055\,
            I => \N__23047\
        );

    \I__4346\ : Odrv12
    port map (
            O => \N__23052\,
            I => \b2v_inst.un4_cuenta_cry_7_c_RNILHBZ0Z8\
        );

    \I__4345\ : LocalMux
    port map (
            O => \N__23047\,
            I => \b2v_inst.un4_cuenta_cry_7_c_RNILHBZ0Z8\
        );

    \I__4344\ : InMux
    port map (
            O => \N__23042\,
            I => \b2v_inst.un4_cuenta_cry_7\
        );

    \I__4343\ : CascadeMux
    port map (
            O => \N__23039\,
            I => \b2v_inst9.data_to_send_10_0_0_0_3_cascade_\
        );

    \I__4342\ : CascadeMux
    port map (
            O => \N__23036\,
            I => \N__23033\
        );

    \I__4341\ : InMux
    port map (
            O => \N__23033\,
            I => \N__23030\
        );

    \I__4340\ : LocalMux
    port map (
            O => \N__23030\,
            I => \b2v_inst9.data_to_sendZ0Z_6\
        );

    \I__4339\ : InMux
    port map (
            O => \N__23027\,
            I => \N__23024\
        );

    \I__4338\ : LocalMux
    port map (
            O => \N__23024\,
            I => \b2v_inst.un1_data_a_escribir_0_sqmuxa_3_i_i_a2_0\
        );

    \I__4337\ : CascadeMux
    port map (
            O => \N__23021\,
            I => \b2v_inst.N_655_cascade_\
        );

    \I__4336\ : InMux
    port map (
            O => \N__23018\,
            I => \N__23011\
        );

    \I__4335\ : InMux
    port map (
            O => \N__23017\,
            I => \N__23006\
        );

    \I__4334\ : InMux
    port map (
            O => \N__23016\,
            I => \N__23006\
        );

    \I__4333\ : CascadeMux
    port map (
            O => \N__23015\,
            I => \N__23001\
        );

    \I__4332\ : CascadeMux
    port map (
            O => \N__23014\,
            I => \N__22997\
        );

    \I__4331\ : LocalMux
    port map (
            O => \N__23011\,
            I => \N__22989\
        );

    \I__4330\ : LocalMux
    port map (
            O => \N__23006\,
            I => \N__22986\
        );

    \I__4329\ : InMux
    port map (
            O => \N__23005\,
            I => \N__22979\
        );

    \I__4328\ : InMux
    port map (
            O => \N__23004\,
            I => \N__22979\
        );

    \I__4327\ : InMux
    port map (
            O => \N__23001\,
            I => \N__22979\
        );

    \I__4326\ : InMux
    port map (
            O => \N__23000\,
            I => \N__22972\
        );

    \I__4325\ : InMux
    port map (
            O => \N__22997\,
            I => \N__22972\
        );

    \I__4324\ : InMux
    port map (
            O => \N__22996\,
            I => \N__22972\
        );

    \I__4323\ : CascadeMux
    port map (
            O => \N__22995\,
            I => \N__22969\
        );

    \I__4322\ : InMux
    port map (
            O => \N__22994\,
            I => \N__22963\
        );

    \I__4321\ : InMux
    port map (
            O => \N__22993\,
            I => \N__22963\
        );

    \I__4320\ : InMux
    port map (
            O => \N__22992\,
            I => \N__22960\
        );

    \I__4319\ : Span4Mux_h
    port map (
            O => \N__22989\,
            I => \N__22951\
        );

    \I__4318\ : Span4Mux_h
    port map (
            O => \N__22986\,
            I => \N__22951\
        );

    \I__4317\ : LocalMux
    port map (
            O => \N__22979\,
            I => \N__22951\
        );

    \I__4316\ : LocalMux
    port map (
            O => \N__22972\,
            I => \N__22951\
        );

    \I__4315\ : InMux
    port map (
            O => \N__22969\,
            I => \N__22946\
        );

    \I__4314\ : InMux
    port map (
            O => \N__22968\,
            I => \N__22946\
        );

    \I__4313\ : LocalMux
    port map (
            O => \N__22963\,
            I => \b2v_inst.state18_li_0\
        );

    \I__4312\ : LocalMux
    port map (
            O => \N__22960\,
            I => \b2v_inst.state18_li_0\
        );

    \I__4311\ : Odrv4
    port map (
            O => \N__22951\,
            I => \b2v_inst.state18_li_0\
        );

    \I__4310\ : LocalMux
    port map (
            O => \N__22946\,
            I => \b2v_inst.state18_li_0\
        );

    \I__4309\ : InMux
    port map (
            O => \N__22937\,
            I => \N__22933\
        );

    \I__4308\ : InMux
    port map (
            O => \N__22936\,
            I => \N__22930\
        );

    \I__4307\ : LocalMux
    port map (
            O => \N__22933\,
            I => \b2v_inst.cuenta_RNIR03AZ0Z_1\
        );

    \I__4306\ : LocalMux
    port map (
            O => \N__22930\,
            I => \b2v_inst.cuenta_RNIR03AZ0Z_1\
        );

    \I__4305\ : CascadeMux
    port map (
            O => \N__22925\,
            I => \N__22920\
        );

    \I__4304\ : CascadeMux
    port map (
            O => \N__22924\,
            I => \N__22917\
        );

    \I__4303\ : CascadeMux
    port map (
            O => \N__22923\,
            I => \N__22912\
        );

    \I__4302\ : InMux
    port map (
            O => \N__22920\,
            I => \N__22909\
        );

    \I__4301\ : InMux
    port map (
            O => \N__22917\,
            I => \N__22904\
        );

    \I__4300\ : InMux
    port map (
            O => \N__22916\,
            I => \N__22897\
        );

    \I__4299\ : InMux
    port map (
            O => \N__22915\,
            I => \N__22897\
        );

    \I__4298\ : InMux
    port map (
            O => \N__22912\,
            I => \N__22897\
        );

    \I__4297\ : LocalMux
    port map (
            O => \N__22909\,
            I => \N__22894\
        );

    \I__4296\ : InMux
    port map (
            O => \N__22908\,
            I => \N__22890\
        );

    \I__4295\ : InMux
    port map (
            O => \N__22907\,
            I => \N__22887\
        );

    \I__4294\ : LocalMux
    port map (
            O => \N__22904\,
            I => \N__22884\
        );

    \I__4293\ : LocalMux
    port map (
            O => \N__22897\,
            I => \N__22881\
        );

    \I__4292\ : Span4Mux_v
    port map (
            O => \N__22894\,
            I => \N__22878\
        );

    \I__4291\ : InMux
    port map (
            O => \N__22893\,
            I => \N__22875\
        );

    \I__4290\ : LocalMux
    port map (
            O => \N__22890\,
            I => \N__22872\
        );

    \I__4289\ : LocalMux
    port map (
            O => \N__22887\,
            I => \N__22869\
        );

    \I__4288\ : Span4Mux_v
    port map (
            O => \N__22884\,
            I => \N__22864\
        );

    \I__4287\ : Span4Mux_h
    port map (
            O => \N__22881\,
            I => \N__22864\
        );

    \I__4286\ : Span4Mux_h
    port map (
            O => \N__22878\,
            I => \N__22859\
        );

    \I__4285\ : LocalMux
    port map (
            O => \N__22875\,
            I => \N__22856\
        );

    \I__4284\ : Span12Mux_h
    port map (
            O => \N__22872\,
            I => \N__22853\
        );

    \I__4283\ : Span4Mux_h
    port map (
            O => \N__22869\,
            I => \N__22848\
        );

    \I__4282\ : Span4Mux_h
    port map (
            O => \N__22864\,
            I => \N__22848\
        );

    \I__4281\ : InMux
    port map (
            O => \N__22863\,
            I => \N__22843\
        );

    \I__4280\ : InMux
    port map (
            O => \N__22862\,
            I => \N__22843\
        );

    \I__4279\ : Odrv4
    port map (
            O => \N__22859\,
            I => \b2v_inst1.r_SM_MainZ0Z_1\
        );

    \I__4278\ : Odrv12
    port map (
            O => \N__22856\,
            I => \b2v_inst1.r_SM_MainZ0Z_1\
        );

    \I__4277\ : Odrv12
    port map (
            O => \N__22853\,
            I => \b2v_inst1.r_SM_MainZ0Z_1\
        );

    \I__4276\ : Odrv4
    port map (
            O => \N__22848\,
            I => \b2v_inst1.r_SM_MainZ0Z_1\
        );

    \I__4275\ : LocalMux
    port map (
            O => \N__22843\,
            I => \b2v_inst1.r_SM_MainZ0Z_1\
        );

    \I__4274\ : InMux
    port map (
            O => \N__22832\,
            I => \N__22823\
        );

    \I__4273\ : InMux
    port map (
            O => \N__22831\,
            I => \N__22820\
        );

    \I__4272\ : InMux
    port map (
            O => \N__22830\,
            I => \N__22817\
        );

    \I__4271\ : InMux
    port map (
            O => \N__22829\,
            I => \N__22813\
        );

    \I__4270\ : InMux
    port map (
            O => \N__22828\,
            I => \N__22809\
        );

    \I__4269\ : InMux
    port map (
            O => \N__22827\,
            I => \N__22804\
        );

    \I__4268\ : InMux
    port map (
            O => \N__22826\,
            I => \N__22804\
        );

    \I__4267\ : LocalMux
    port map (
            O => \N__22823\,
            I => \N__22801\
        );

    \I__4266\ : LocalMux
    port map (
            O => \N__22820\,
            I => \N__22796\
        );

    \I__4265\ : LocalMux
    port map (
            O => \N__22817\,
            I => \N__22796\
        );

    \I__4264\ : InMux
    port map (
            O => \N__22816\,
            I => \N__22793\
        );

    \I__4263\ : LocalMux
    port map (
            O => \N__22813\,
            I => \N__22790\
        );

    \I__4262\ : InMux
    port map (
            O => \N__22812\,
            I => \N__22787\
        );

    \I__4261\ : LocalMux
    port map (
            O => \N__22809\,
            I => \N__22782\
        );

    \I__4260\ : LocalMux
    port map (
            O => \N__22804\,
            I => \N__22777\
        );

    \I__4259\ : Span4Mux_h
    port map (
            O => \N__22801\,
            I => \N__22777\
        );

    \I__4258\ : Span4Mux_v
    port map (
            O => \N__22796\,
            I => \N__22770\
        );

    \I__4257\ : LocalMux
    port map (
            O => \N__22793\,
            I => \N__22770\
        );

    \I__4256\ : Span4Mux_h
    port map (
            O => \N__22790\,
            I => \N__22770\
        );

    \I__4255\ : LocalMux
    port map (
            O => \N__22787\,
            I => \N__22767\
        );

    \I__4254\ : InMux
    port map (
            O => \N__22786\,
            I => \N__22762\
        );

    \I__4253\ : InMux
    port map (
            O => \N__22785\,
            I => \N__22762\
        );

    \I__4252\ : Span4Mux_h
    port map (
            O => \N__22782\,
            I => \N__22759\
        );

    \I__4251\ : Span4Mux_h
    port map (
            O => \N__22777\,
            I => \N__22756\
        );

    \I__4250\ : Span4Mux_h
    port map (
            O => \N__22770\,
            I => \N__22753\
        );

    \I__4249\ : Span12Mux_h
    port map (
            O => \N__22767\,
            I => \N__22748\
        );

    \I__4248\ : LocalMux
    port map (
            O => \N__22762\,
            I => \N__22748\
        );

    \I__4247\ : Odrv4
    port map (
            O => \N__22759\,
            I => \b2v_inst1.r_RX_DataZ0\
        );

    \I__4246\ : Odrv4
    port map (
            O => \N__22756\,
            I => \b2v_inst1.r_RX_DataZ0\
        );

    \I__4245\ : Odrv4
    port map (
            O => \N__22753\,
            I => \b2v_inst1.r_RX_DataZ0\
        );

    \I__4244\ : Odrv12
    port map (
            O => \N__22748\,
            I => \b2v_inst1.r_RX_DataZ0\
        );

    \I__4243\ : InMux
    port map (
            O => \N__22739\,
            I => \N__22734\
        );

    \I__4242\ : InMux
    port map (
            O => \N__22738\,
            I => \N__22728\
        );

    \I__4241\ : InMux
    port map (
            O => \N__22737\,
            I => \N__22728\
        );

    \I__4240\ : LocalMux
    port map (
            O => \N__22734\,
            I => \N__22725\
        );

    \I__4239\ : CascadeMux
    port map (
            O => \N__22733\,
            I => \N__22721\
        );

    \I__4238\ : LocalMux
    port map (
            O => \N__22728\,
            I => \N__22717\
        );

    \I__4237\ : Span4Mux_h
    port map (
            O => \N__22725\,
            I => \N__22714\
        );

    \I__4236\ : InMux
    port map (
            O => \N__22724\,
            I => \N__22710\
        );

    \I__4235\ : InMux
    port map (
            O => \N__22721\,
            I => \N__22707\
        );

    \I__4234\ : InMux
    port map (
            O => \N__22720\,
            I => \N__22704\
        );

    \I__4233\ : Span4Mux_v
    port map (
            O => \N__22717\,
            I => \N__22701\
        );

    \I__4232\ : Span4Mux_h
    port map (
            O => \N__22714\,
            I => \N__22698\
        );

    \I__4231\ : InMux
    port map (
            O => \N__22713\,
            I => \N__22695\
        );

    \I__4230\ : LocalMux
    port map (
            O => \N__22710\,
            I => \N__22690\
        );

    \I__4229\ : LocalMux
    port map (
            O => \N__22707\,
            I => \N__22690\
        );

    \I__4228\ : LocalMux
    port map (
            O => \N__22704\,
            I => \N__22685\
        );

    \I__4227\ : Span4Mux_h
    port map (
            O => \N__22701\,
            I => \N__22685\
        );

    \I__4226\ : Odrv4
    port map (
            O => \N__22698\,
            I => \b2v_inst1.r_SM_MainZ0Z_2\
        );

    \I__4225\ : LocalMux
    port map (
            O => \N__22695\,
            I => \b2v_inst1.r_SM_MainZ0Z_2\
        );

    \I__4224\ : Odrv4
    port map (
            O => \N__22690\,
            I => \b2v_inst1.r_SM_MainZ0Z_2\
        );

    \I__4223\ : Odrv4
    port map (
            O => \N__22685\,
            I => \b2v_inst1.r_SM_MainZ0Z_2\
        );

    \I__4222\ : InMux
    port map (
            O => \N__22676\,
            I => \N__22673\
        );

    \I__4221\ : LocalMux
    port map (
            O => \N__22673\,
            I => \N__22670\
        );

    \I__4220\ : Span4Mux_v
    port map (
            O => \N__22670\,
            I => \N__22667\
        );

    \I__4219\ : Span4Mux_h
    port map (
            O => \N__22667\,
            I => \N__22664\
        );

    \I__4218\ : Odrv4
    port map (
            O => \N__22664\,
            I => \b2v_inst1.m13_i_2\
        );

    \I__4217\ : CascadeMux
    port map (
            O => \N__22661\,
            I => \b2v_inst1.N_95_cascade_\
        );

    \I__4216\ : InMux
    port map (
            O => \N__22658\,
            I => \N__22655\
        );

    \I__4215\ : LocalMux
    port map (
            O => \N__22655\,
            I => \N__22652\
        );

    \I__4214\ : Span4Mux_v
    port map (
            O => \N__22652\,
            I => \N__22649\
        );

    \I__4213\ : Span4Mux_h
    port map (
            O => \N__22649\,
            I => \N__22646\
        );

    \I__4212\ : Odrv4
    port map (
            O => \N__22646\,
            I => \b2v_inst1.N_96\
        );

    \I__4211\ : InMux
    port map (
            O => \N__22643\,
            I => \N__22639\
        );

    \I__4210\ : InMux
    port map (
            O => \N__22642\,
            I => \N__22635\
        );

    \I__4209\ : LocalMux
    port map (
            O => \N__22639\,
            I => \N__22631\
        );

    \I__4208\ : InMux
    port map (
            O => \N__22638\,
            I => \N__22628\
        );

    \I__4207\ : LocalMux
    port map (
            O => \N__22635\,
            I => \N__22621\
        );

    \I__4206\ : InMux
    port map (
            O => \N__22634\,
            I => \N__22616\
        );

    \I__4205\ : Span4Mux_v
    port map (
            O => \N__22631\,
            I => \N__22611\
        );

    \I__4204\ : LocalMux
    port map (
            O => \N__22628\,
            I => \N__22611\
        );

    \I__4203\ : InMux
    port map (
            O => \N__22627\,
            I => \N__22608\
        );

    \I__4202\ : InMux
    port map (
            O => \N__22626\,
            I => \N__22601\
        );

    \I__4201\ : InMux
    port map (
            O => \N__22625\,
            I => \N__22601\
        );

    \I__4200\ : InMux
    port map (
            O => \N__22624\,
            I => \N__22601\
        );

    \I__4199\ : Span4Mux_h
    port map (
            O => \N__22621\,
            I => \N__22598\
        );

    \I__4198\ : InMux
    port map (
            O => \N__22620\,
            I => \N__22593\
        );

    \I__4197\ : InMux
    port map (
            O => \N__22619\,
            I => \N__22593\
        );

    \I__4196\ : LocalMux
    port map (
            O => \N__22616\,
            I => \N__22590\
        );

    \I__4195\ : Span4Mux_v
    port map (
            O => \N__22611\,
            I => \N__22583\
        );

    \I__4194\ : LocalMux
    port map (
            O => \N__22608\,
            I => \N__22583\
        );

    \I__4193\ : LocalMux
    port map (
            O => \N__22601\,
            I => \N__22583\
        );

    \I__4192\ : Span4Mux_h
    port map (
            O => \N__22598\,
            I => \N__22580\
        );

    \I__4191\ : LocalMux
    port map (
            O => \N__22593\,
            I => \N__22577\
        );

    \I__4190\ : Span4Mux_h
    port map (
            O => \N__22590\,
            I => \N__22574\
        );

    \I__4189\ : Span4Mux_v
    port map (
            O => \N__22583\,
            I => \N__22570\
        );

    \I__4188\ : Span4Mux_v
    port map (
            O => \N__22580\,
            I => \N__22567\
        );

    \I__4187\ : Span4Mux_v
    port map (
            O => \N__22577\,
            I => \N__22564\
        );

    \I__4186\ : Span4Mux_h
    port map (
            O => \N__22574\,
            I => \N__22561\
        );

    \I__4185\ : InMux
    port map (
            O => \N__22573\,
            I => \N__22558\
        );

    \I__4184\ : Span4Mux_h
    port map (
            O => \N__22570\,
            I => \N__22555\
        );

    \I__4183\ : Odrv4
    port map (
            O => \N__22567\,
            I => \b2v_inst1.r_SM_MainZ0Z_0\
        );

    \I__4182\ : Odrv4
    port map (
            O => \N__22564\,
            I => \b2v_inst1.r_SM_MainZ0Z_0\
        );

    \I__4181\ : Odrv4
    port map (
            O => \N__22561\,
            I => \b2v_inst1.r_SM_MainZ0Z_0\
        );

    \I__4180\ : LocalMux
    port map (
            O => \N__22558\,
            I => \b2v_inst1.r_SM_MainZ0Z_0\
        );

    \I__4179\ : Odrv4
    port map (
            O => \N__22555\,
            I => \b2v_inst1.r_SM_MainZ0Z_0\
        );

    \I__4178\ : InMux
    port map (
            O => \N__22544\,
            I => \N__22541\
        );

    \I__4177\ : LocalMux
    port map (
            O => \N__22541\,
            I => \N__22538\
        );

    \I__4176\ : Span4Mux_v
    port map (
            O => \N__22538\,
            I => \N__22535\
        );

    \I__4175\ : Odrv4
    port map (
            O => \N__22535\,
            I => \b2v_inst.dir_memZ0Z_5\
        );

    \I__4174\ : CascadeMux
    port map (
            O => \N__22532\,
            I => \N__22528\
        );

    \I__4173\ : InMux
    port map (
            O => \N__22531\,
            I => \N__22520\
        );

    \I__4172\ : InMux
    port map (
            O => \N__22528\,
            I => \N__22515\
        );

    \I__4171\ : InMux
    port map (
            O => \N__22527\,
            I => \N__22515\
        );

    \I__4170\ : InMux
    port map (
            O => \N__22526\,
            I => \N__22512\
        );

    \I__4169\ : InMux
    port map (
            O => \N__22525\,
            I => \N__22508\
        );

    \I__4168\ : InMux
    port map (
            O => \N__22524\,
            I => \N__22505\
        );

    \I__4167\ : InMux
    port map (
            O => \N__22523\,
            I => \N__22502\
        );

    \I__4166\ : LocalMux
    port map (
            O => \N__22520\,
            I => \N__22494\
        );

    \I__4165\ : LocalMux
    port map (
            O => \N__22515\,
            I => \N__22494\
        );

    \I__4164\ : LocalMux
    port map (
            O => \N__22512\,
            I => \N__22491\
        );

    \I__4163\ : InMux
    port map (
            O => \N__22511\,
            I => \N__22488\
        );

    \I__4162\ : LocalMux
    port map (
            O => \N__22508\,
            I => \N__22481\
        );

    \I__4161\ : LocalMux
    port map (
            O => \N__22505\,
            I => \N__22481\
        );

    \I__4160\ : LocalMux
    port map (
            O => \N__22502\,
            I => \N__22481\
        );

    \I__4159\ : InMux
    port map (
            O => \N__22501\,
            I => \N__22476\
        );

    \I__4158\ : InMux
    port map (
            O => \N__22500\,
            I => \N__22476\
        );

    \I__4157\ : InMux
    port map (
            O => \N__22499\,
            I => \N__22473\
        );

    \I__4156\ : Odrv4
    port map (
            O => \N__22494\,
            I => \b2v_inst.N_450_i_1\
        );

    \I__4155\ : Odrv4
    port map (
            O => \N__22491\,
            I => \b2v_inst.N_450_i_1\
        );

    \I__4154\ : LocalMux
    port map (
            O => \N__22488\,
            I => \b2v_inst.N_450_i_1\
        );

    \I__4153\ : Odrv4
    port map (
            O => \N__22481\,
            I => \b2v_inst.N_450_i_1\
        );

    \I__4152\ : LocalMux
    port map (
            O => \N__22476\,
            I => \b2v_inst.N_450_i_1\
        );

    \I__4151\ : LocalMux
    port map (
            O => \N__22473\,
            I => \b2v_inst.N_450_i_1\
        );

    \I__4150\ : CascadeMux
    port map (
            O => \N__22460\,
            I => \N__22457\
        );

    \I__4149\ : InMux
    port map (
            O => \N__22457\,
            I => \N__22454\
        );

    \I__4148\ : LocalMux
    port map (
            O => \N__22454\,
            I => \N__22451\
        );

    \I__4147\ : Span4Mux_h
    port map (
            O => \N__22451\,
            I => \N__22448\
        );

    \I__4146\ : Odrv4
    port map (
            O => \N__22448\,
            I => \b2v_inst.dir_mem_2Z0Z_5\
        );

    \I__4145\ : CascadeMux
    port map (
            O => \N__22445\,
            I => \N__22440\
        );

    \I__4144\ : InMux
    port map (
            O => \N__22444\,
            I => \N__22435\
        );

    \I__4143\ : InMux
    port map (
            O => \N__22443\,
            I => \N__22432\
        );

    \I__4142\ : InMux
    port map (
            O => \N__22440\,
            I => \N__22426\
        );

    \I__4141\ : InMux
    port map (
            O => \N__22439\,
            I => \N__22421\
        );

    \I__4140\ : InMux
    port map (
            O => \N__22438\,
            I => \N__22421\
        );

    \I__4139\ : LocalMux
    port map (
            O => \N__22435\,
            I => \N__22415\
        );

    \I__4138\ : LocalMux
    port map (
            O => \N__22432\,
            I => \N__22415\
        );

    \I__4137\ : InMux
    port map (
            O => \N__22431\,
            I => \N__22410\
        );

    \I__4136\ : InMux
    port map (
            O => \N__22430\,
            I => \N__22410\
        );

    \I__4135\ : InMux
    port map (
            O => \N__22429\,
            I => \N__22407\
        );

    \I__4134\ : LocalMux
    port map (
            O => \N__22426\,
            I => \N__22399\
        );

    \I__4133\ : LocalMux
    port map (
            O => \N__22421\,
            I => \N__22399\
        );

    \I__4132\ : InMux
    port map (
            O => \N__22420\,
            I => \N__22396\
        );

    \I__4131\ : Span4Mux_v
    port map (
            O => \N__22415\,
            I => \N__22389\
        );

    \I__4130\ : LocalMux
    port map (
            O => \N__22410\,
            I => \N__22389\
        );

    \I__4129\ : LocalMux
    port map (
            O => \N__22407\,
            I => \N__22389\
        );

    \I__4128\ : InMux
    port map (
            O => \N__22406\,
            I => \N__22386\
        );

    \I__4127\ : InMux
    port map (
            O => \N__22405\,
            I => \N__22381\
        );

    \I__4126\ : InMux
    port map (
            O => \N__22404\,
            I => \N__22381\
        );

    \I__4125\ : Odrv4
    port map (
            O => \N__22399\,
            I => \b2v_inst.N_489\
        );

    \I__4124\ : LocalMux
    port map (
            O => \N__22396\,
            I => \b2v_inst.N_489\
        );

    \I__4123\ : Odrv4
    port map (
            O => \N__22389\,
            I => \b2v_inst.N_489\
        );

    \I__4122\ : LocalMux
    port map (
            O => \N__22386\,
            I => \b2v_inst.N_489\
        );

    \I__4121\ : LocalMux
    port map (
            O => \N__22381\,
            I => \b2v_inst.N_489\
        );

    \I__4120\ : CascadeMux
    port map (
            O => \N__22370\,
            I => \b2v_inst9.data_to_send_10_0_0_0_5_cascade_\
        );

    \I__4119\ : CascadeMux
    port map (
            O => \N__22367\,
            I => \N__22364\
        );

    \I__4118\ : InMux
    port map (
            O => \N__22364\,
            I => \N__22361\
        );

    \I__4117\ : LocalMux
    port map (
            O => \N__22361\,
            I => \b2v_inst9.data_to_sendZ0Z_5\
        );

    \I__4116\ : CascadeMux
    port map (
            O => \N__22358\,
            I => \N__22355\
        );

    \I__4115\ : InMux
    port map (
            O => \N__22355\,
            I => \N__22352\
        );

    \I__4114\ : LocalMux
    port map (
            O => \N__22352\,
            I => \N__22349\
        );

    \I__4113\ : Odrv4
    port map (
            O => \N__22349\,
            I => \b2v_inst.dir_mem_2_RNO_0Z0Z_5\
        );

    \I__4112\ : InMux
    port map (
            O => \N__22346\,
            I => \b2v_inst.un2_dir_mem_2_cry_4\
        );

    \I__4111\ : CascadeMux
    port map (
            O => \N__22343\,
            I => \N__22340\
        );

    \I__4110\ : InMux
    port map (
            O => \N__22340\,
            I => \N__22337\
        );

    \I__4109\ : LocalMux
    port map (
            O => \N__22337\,
            I => \N__22334\
        );

    \I__4108\ : Odrv4
    port map (
            O => \N__22334\,
            I => \b2v_inst.dir_mem_2_RNO_0Z0Z_6\
        );

    \I__4107\ : InMux
    port map (
            O => \N__22331\,
            I => \b2v_inst.un2_dir_mem_2_cry_5\
        );

    \I__4106\ : CascadeMux
    port map (
            O => \N__22328\,
            I => \N__22325\
        );

    \I__4105\ : InMux
    port map (
            O => \N__22325\,
            I => \N__22322\
        );

    \I__4104\ : LocalMux
    port map (
            O => \N__22322\,
            I => \N__22319\
        );

    \I__4103\ : Odrv4
    port map (
            O => \N__22319\,
            I => \b2v_inst.dir_mem_2_RNO_0Z0Z_7\
        );

    \I__4102\ : InMux
    port map (
            O => \N__22316\,
            I => \b2v_inst.un2_dir_mem_2_cry_6\
        );

    \I__4101\ : InMux
    port map (
            O => \N__22313\,
            I => \N__22310\
        );

    \I__4100\ : LocalMux
    port map (
            O => \N__22310\,
            I => \N__22307\
        );

    \I__4099\ : Odrv4
    port map (
            O => \N__22307\,
            I => \b2v_inst.dir_mem_2_RNO_0Z0Z_8\
        );

    \I__4098\ : InMux
    port map (
            O => \N__22304\,
            I => \bfn_13_7_0_\
        );

    \I__4097\ : CascadeMux
    port map (
            O => \N__22301\,
            I => \N__22298\
        );

    \I__4096\ : InMux
    port map (
            O => \N__22298\,
            I => \N__22295\
        );

    \I__4095\ : LocalMux
    port map (
            O => \N__22295\,
            I => \b2v_inst.dir_mem_2_RNO_0Z0Z_9\
        );

    \I__4094\ : InMux
    port map (
            O => \N__22292\,
            I => \b2v_inst.un2_dir_mem_2_cry_8\
        );

    \I__4093\ : InMux
    port map (
            O => \N__22289\,
            I => \b2v_inst.un2_dir_mem_2_cry_9\
        );

    \I__4092\ : CascadeMux
    port map (
            O => \N__22286\,
            I => \N__22283\
        );

    \I__4091\ : InMux
    port map (
            O => \N__22283\,
            I => \N__22280\
        );

    \I__4090\ : LocalMux
    port map (
            O => \N__22280\,
            I => \b2v_inst.dir_mem_2_RNO_0Z0Z_10\
        );

    \I__4089\ : InMux
    port map (
            O => \N__22277\,
            I => \N__22274\
        );

    \I__4088\ : LocalMux
    port map (
            O => \N__22274\,
            I => \b2v_inst1.r_RX_Data_RZ0\
        );

    \I__4087\ : CascadeMux
    port map (
            O => \N__22271\,
            I => \N__22267\
        );

    \I__4086\ : InMux
    port map (
            O => \N__22270\,
            I => \N__22259\
        );

    \I__4085\ : InMux
    port map (
            O => \N__22267\,
            I => \N__22259\
        );

    \I__4084\ : InMux
    port map (
            O => \N__22266\,
            I => \N__22259\
        );

    \I__4083\ : LocalMux
    port map (
            O => \N__22259\,
            I => \N__22256\
        );

    \I__4082\ : Sp12to4
    port map (
            O => \N__22256\,
            I => \N__22253\
        );

    \I__4081\ : Odrv12
    port map (
            O => \N__22253\,
            I => \b2v_inst.un9_indice_0_a2_2\
        );

    \I__4080\ : CascadeMux
    port map (
            O => \N__22250\,
            I => \N__22245\
        );

    \I__4079\ : InMux
    port map (
            O => \N__22249\,
            I => \N__22238\
        );

    \I__4078\ : InMux
    port map (
            O => \N__22248\,
            I => \N__22238\
        );

    \I__4077\ : InMux
    port map (
            O => \N__22245\,
            I => \N__22238\
        );

    \I__4076\ : LocalMux
    port map (
            O => \N__22238\,
            I => \N__22234\
        );

    \I__4075\ : InMux
    port map (
            O => \N__22237\,
            I => \N__22231\
        );

    \I__4074\ : Span4Mux_h
    port map (
            O => \N__22234\,
            I => \N__22228\
        );

    \I__4073\ : LocalMux
    port map (
            O => \N__22231\,
            I => \N__22225\
        );

    \I__4072\ : Span4Mux_v
    port map (
            O => \N__22228\,
            I => \N__22222\
        );

    \I__4071\ : Span4Mux_v
    port map (
            O => \N__22225\,
            I => \N__22217\
        );

    \I__4070\ : Span4Mux_v
    port map (
            O => \N__22222\,
            I => \N__22217\
        );

    \I__4069\ : Odrv4
    port map (
            O => \N__22217\,
            I => \b2v_inst.un9_indice_0_a2_3\
        );

    \I__4068\ : InMux
    port map (
            O => \N__22214\,
            I => \N__22211\
        );

    \I__4067\ : LocalMux
    port map (
            O => \N__22211\,
            I => \N__22208\
        );

    \I__4066\ : Span4Mux_h
    port map (
            O => \N__22208\,
            I => \N__22205\
        );

    \I__4065\ : Span4Mux_h
    port map (
            O => \N__22205\,
            I => \N__22202\
        );

    \I__4064\ : Odrv4
    port map (
            O => \N__22202\,
            I => \b2v_inst.dir_mem_RNO_0Z0Z_5\
        );

    \I__4063\ : CascadeMux
    port map (
            O => \N__22199\,
            I => \b2v_inst.un9_indice_0_a2_2_cascade_\
        );

    \I__4062\ : CEMux
    port map (
            O => \N__22196\,
            I => \N__22192\
        );

    \I__4061\ : CEMux
    port map (
            O => \N__22195\,
            I => \N__22189\
        );

    \I__4060\ : LocalMux
    port map (
            O => \N__22192\,
            I => \N__22183\
        );

    \I__4059\ : LocalMux
    port map (
            O => \N__22189\,
            I => \N__22180\
        );

    \I__4058\ : CEMux
    port map (
            O => \N__22188\,
            I => \N__22177\
        );

    \I__4057\ : CEMux
    port map (
            O => \N__22187\,
            I => \N__22174\
        );

    \I__4056\ : CEMux
    port map (
            O => \N__22186\,
            I => \N__22171\
        );

    \I__4055\ : Span4Mux_v
    port map (
            O => \N__22183\,
            I => \N__22166\
        );

    \I__4054\ : Span4Mux_v
    port map (
            O => \N__22180\,
            I => \N__22163\
        );

    \I__4053\ : LocalMux
    port map (
            O => \N__22177\,
            I => \N__22160\
        );

    \I__4052\ : LocalMux
    port map (
            O => \N__22174\,
            I => \N__22157\
        );

    \I__4051\ : LocalMux
    port map (
            O => \N__22171\,
            I => \N__22154\
        );

    \I__4050\ : CEMux
    port map (
            O => \N__22170\,
            I => \N__22151\
        );

    \I__4049\ : CascadeMux
    port map (
            O => \N__22169\,
            I => \N__22146\
        );

    \I__4048\ : Span4Mux_h
    port map (
            O => \N__22166\,
            I => \N__22139\
        );

    \I__4047\ : Span4Mux_h
    port map (
            O => \N__22163\,
            I => \N__22139\
        );

    \I__4046\ : Span4Mux_h
    port map (
            O => \N__22160\,
            I => \N__22139\
        );

    \I__4045\ : Span4Mux_v
    port map (
            O => \N__22157\,
            I => \N__22136\
        );

    \I__4044\ : Span4Mux_h
    port map (
            O => \N__22154\,
            I => \N__22131\
        );

    \I__4043\ : LocalMux
    port map (
            O => \N__22151\,
            I => \N__22131\
        );

    \I__4042\ : InMux
    port map (
            O => \N__22150\,
            I => \N__22128\
        );

    \I__4041\ : InMux
    port map (
            O => \N__22149\,
            I => \N__22125\
        );

    \I__4040\ : InMux
    port map (
            O => \N__22146\,
            I => \N__22122\
        );

    \I__4039\ : Odrv4
    port map (
            O => \N__22139\,
            I => \b2v_inst.stateZ0Z_28\
        );

    \I__4038\ : Odrv4
    port map (
            O => \N__22136\,
            I => \b2v_inst.stateZ0Z_28\
        );

    \I__4037\ : Odrv4
    port map (
            O => \N__22131\,
            I => \b2v_inst.stateZ0Z_28\
        );

    \I__4036\ : LocalMux
    port map (
            O => \N__22128\,
            I => \b2v_inst.stateZ0Z_28\
        );

    \I__4035\ : LocalMux
    port map (
            O => \N__22125\,
            I => \b2v_inst.stateZ0Z_28\
        );

    \I__4034\ : LocalMux
    port map (
            O => \N__22122\,
            I => \b2v_inst.stateZ0Z_28\
        );

    \I__4033\ : InMux
    port map (
            O => \N__22109\,
            I => \N__22097\
        );

    \I__4032\ : InMux
    port map (
            O => \N__22108\,
            I => \N__22097\
        );

    \I__4031\ : InMux
    port map (
            O => \N__22107\,
            I => \N__22097\
        );

    \I__4030\ : InMux
    port map (
            O => \N__22106\,
            I => \N__22097\
        );

    \I__4029\ : LocalMux
    port map (
            O => \N__22097\,
            I => \N__22092\
        );

    \I__4028\ : InMux
    port map (
            O => \N__22096\,
            I => \N__22089\
        );

    \I__4027\ : InMux
    port map (
            O => \N__22095\,
            I => \N__22082\
        );

    \I__4026\ : Sp12to4
    port map (
            O => \N__22092\,
            I => \N__22077\
        );

    \I__4025\ : LocalMux
    port map (
            O => \N__22089\,
            I => \N__22077\
        );

    \I__4024\ : InMux
    port map (
            O => \N__22088\,
            I => \N__22070\
        );

    \I__4023\ : InMux
    port map (
            O => \N__22087\,
            I => \N__22070\
        );

    \I__4022\ : InMux
    port map (
            O => \N__22086\,
            I => \N__22070\
        );

    \I__4021\ : InMux
    port map (
            O => \N__22085\,
            I => \N__22067\
        );

    \I__4020\ : LocalMux
    port map (
            O => \N__22082\,
            I => \b2v_inst.N_432_1\
        );

    \I__4019\ : Odrv12
    port map (
            O => \N__22077\,
            I => \b2v_inst.N_432_1\
        );

    \I__4018\ : LocalMux
    port map (
            O => \N__22070\,
            I => \b2v_inst.N_432_1\
        );

    \I__4017\ : LocalMux
    port map (
            O => \N__22067\,
            I => \b2v_inst.N_432_1\
        );

    \I__4016\ : CEMux
    port map (
            O => \N__22058\,
            I => \N__22053\
        );

    \I__4015\ : CEMux
    port map (
            O => \N__22057\,
            I => \N__22050\
        );

    \I__4014\ : CEMux
    port map (
            O => \N__22056\,
            I => \N__22047\
        );

    \I__4013\ : LocalMux
    port map (
            O => \N__22053\,
            I => \N__22043\
        );

    \I__4012\ : LocalMux
    port map (
            O => \N__22050\,
            I => \N__22040\
        );

    \I__4011\ : LocalMux
    port map (
            O => \N__22047\,
            I => \N__22037\
        );

    \I__4010\ : CEMux
    port map (
            O => \N__22046\,
            I => \N__22034\
        );

    \I__4009\ : Span4Mux_h
    port map (
            O => \N__22043\,
            I => \N__22030\
        );

    \I__4008\ : Span4Mux_h
    port map (
            O => \N__22040\,
            I => \N__22027\
        );

    \I__4007\ : Span4Mux_h
    port map (
            O => \N__22037\,
            I => \N__22022\
        );

    \I__4006\ : LocalMux
    port map (
            O => \N__22034\,
            I => \N__22022\
        );

    \I__4005\ : CEMux
    port map (
            O => \N__22033\,
            I => \N__22019\
        );

    \I__4004\ : Span4Mux_h
    port map (
            O => \N__22030\,
            I => \N__22016\
        );

    \I__4003\ : Span4Mux_h
    port map (
            O => \N__22027\,
            I => \N__22011\
        );

    \I__4002\ : Span4Mux_h
    port map (
            O => \N__22022\,
            I => \N__22011\
        );

    \I__4001\ : LocalMux
    port map (
            O => \N__22019\,
            I => \N__22008\
        );

    \I__4000\ : Odrv4
    port map (
            O => \N__22016\,
            I => \b2v_inst.N_442_i\
        );

    \I__3999\ : Odrv4
    port map (
            O => \N__22011\,
            I => \b2v_inst.N_442_i\
        );

    \I__3998\ : Odrv4
    port map (
            O => \N__22008\,
            I => \b2v_inst.N_442_i\
        );

    \I__3997\ : CascadeMux
    port map (
            O => \N__22001\,
            I => \N__21998\
        );

    \I__3996\ : InMux
    port map (
            O => \N__21998\,
            I => \N__21995\
        );

    \I__3995\ : LocalMux
    port map (
            O => \N__21995\,
            I => \N__21992\
        );

    \I__3994\ : Span4Mux_h
    port map (
            O => \N__21992\,
            I => \N__21989\
        );

    \I__3993\ : Odrv4
    port map (
            O => \N__21989\,
            I => \b2v_inst.un2_dir_mem_2_cry_0_THRU_CO\
        );

    \I__3992\ : InMux
    port map (
            O => \N__21986\,
            I => \b2v_inst.un2_dir_mem_2_cry_0\
        );

    \I__3991\ : CascadeMux
    port map (
            O => \N__21983\,
            I => \N__21980\
        );

    \I__3990\ : InMux
    port map (
            O => \N__21980\,
            I => \N__21977\
        );

    \I__3989\ : LocalMux
    port map (
            O => \N__21977\,
            I => \N__21974\
        );

    \I__3988\ : Span4Mux_h
    port map (
            O => \N__21974\,
            I => \N__21971\
        );

    \I__3987\ : Odrv4
    port map (
            O => \N__21971\,
            I => \b2v_inst.dir_mem_2_RNO_0Z0Z_2\
        );

    \I__3986\ : InMux
    port map (
            O => \N__21968\,
            I => \b2v_inst.un2_dir_mem_2_cry_1\
        );

    \I__3985\ : CascadeMux
    port map (
            O => \N__21965\,
            I => \N__21962\
        );

    \I__3984\ : InMux
    port map (
            O => \N__21962\,
            I => \N__21959\
        );

    \I__3983\ : LocalMux
    port map (
            O => \N__21959\,
            I => \N__21956\
        );

    \I__3982\ : Odrv4
    port map (
            O => \N__21956\,
            I => \b2v_inst.dir_mem_2_RNO_0Z0Z_3\
        );

    \I__3981\ : InMux
    port map (
            O => \N__21953\,
            I => \b2v_inst.un2_dir_mem_2_cry_2\
        );

    \I__3980\ : CascadeMux
    port map (
            O => \N__21950\,
            I => \N__21947\
        );

    \I__3979\ : InMux
    port map (
            O => \N__21947\,
            I => \N__21944\
        );

    \I__3978\ : LocalMux
    port map (
            O => \N__21944\,
            I => \N__21941\
        );

    \I__3977\ : Odrv4
    port map (
            O => \N__21941\,
            I => \b2v_inst.dir_mem_2_RNO_0Z0Z_4\
        );

    \I__3976\ : InMux
    port map (
            O => \N__21938\,
            I => \b2v_inst.un2_dir_mem_2_cry_3\
        );

    \I__3975\ : InMux
    port map (
            O => \N__21935\,
            I => \N__21932\
        );

    \I__3974\ : LocalMux
    port map (
            O => \N__21932\,
            I => \N__21928\
        );

    \I__3973\ : InMux
    port map (
            O => \N__21931\,
            I => \N__21925\
        );

    \I__3972\ : Span4Mux_v
    port map (
            O => \N__21928\,
            I => \N__21920\
        );

    \I__3971\ : LocalMux
    port map (
            O => \N__21925\,
            I => \N__21920\
        );

    \I__3970\ : Odrv4
    port map (
            O => \N__21920\,
            I => \b2v_inst.state_ns_0_i_o2_8_23\
        );

    \I__3969\ : InMux
    port map (
            O => \N__21917\,
            I => \N__21914\
        );

    \I__3968\ : LocalMux
    port map (
            O => \N__21914\,
            I => \N__21911\
        );

    \I__3967\ : Span4Mux_h
    port map (
            O => \N__21911\,
            I => \N__21908\
        );

    \I__3966\ : Span4Mux_v
    port map (
            O => \N__21908\,
            I => \N__21905\
        );

    \I__3965\ : Span4Mux_h
    port map (
            O => \N__21905\,
            I => \N__21902\
        );

    \I__3964\ : Odrv4
    port map (
            O => \N__21902\,
            I => \N_550_i\
        );

    \I__3963\ : InMux
    port map (
            O => \N__21899\,
            I => \N__21896\
        );

    \I__3962\ : LocalMux
    port map (
            O => \N__21896\,
            I => \b2v_inst.state_fastZ0Z_32\
        );

    \I__3961\ : InMux
    port map (
            O => \N__21893\,
            I => \N__21883\
        );

    \I__3960\ : InMux
    port map (
            O => \N__21892\,
            I => \N__21883\
        );

    \I__3959\ : CascadeMux
    port map (
            O => \N__21891\,
            I => \N__21879\
        );

    \I__3958\ : InMux
    port map (
            O => \N__21890\,
            I => \N__21871\
        );

    \I__3957\ : InMux
    port map (
            O => \N__21889\,
            I => \N__21871\
        );

    \I__3956\ : InMux
    port map (
            O => \N__21888\,
            I => \N__21871\
        );

    \I__3955\ : LocalMux
    port map (
            O => \N__21883\,
            I => \N__21868\
        );

    \I__3954\ : InMux
    port map (
            O => \N__21882\,
            I => \N__21865\
        );

    \I__3953\ : InMux
    port map (
            O => \N__21879\,
            I => \N__21860\
        );

    \I__3952\ : InMux
    port map (
            O => \N__21878\,
            I => \N__21857\
        );

    \I__3951\ : LocalMux
    port map (
            O => \N__21871\,
            I => \N__21854\
        );

    \I__3950\ : Span4Mux_h
    port map (
            O => \N__21868\,
            I => \N__21851\
        );

    \I__3949\ : LocalMux
    port map (
            O => \N__21865\,
            I => \N__21848\
        );

    \I__3948\ : InMux
    port map (
            O => \N__21864\,
            I => \N__21845\
        );

    \I__3947\ : InMux
    port map (
            O => \N__21863\,
            I => \N__21842\
        );

    \I__3946\ : LocalMux
    port map (
            O => \N__21860\,
            I => \b2v_inst.stateZ0Z_5\
        );

    \I__3945\ : LocalMux
    port map (
            O => \N__21857\,
            I => \b2v_inst.stateZ0Z_5\
        );

    \I__3944\ : Odrv4
    port map (
            O => \N__21854\,
            I => \b2v_inst.stateZ0Z_5\
        );

    \I__3943\ : Odrv4
    port map (
            O => \N__21851\,
            I => \b2v_inst.stateZ0Z_5\
        );

    \I__3942\ : Odrv12
    port map (
            O => \N__21848\,
            I => \b2v_inst.stateZ0Z_5\
        );

    \I__3941\ : LocalMux
    port map (
            O => \N__21845\,
            I => \b2v_inst.stateZ0Z_5\
        );

    \I__3940\ : LocalMux
    port map (
            O => \N__21842\,
            I => \b2v_inst.stateZ0Z_5\
        );

    \I__3939\ : InMux
    port map (
            O => \N__21827\,
            I => \N__21824\
        );

    \I__3938\ : LocalMux
    port map (
            O => \N__21824\,
            I => \b2v_inst.addr_ram_energia_ss0_0_i_o2_i_o2_0\
        );

    \I__3937\ : InMux
    port map (
            O => \N__21821\,
            I => \N__21818\
        );

    \I__3936\ : LocalMux
    port map (
            O => \N__21818\,
            I => \N__21815\
        );

    \I__3935\ : Span12Mux_h
    port map (
            O => \N__21815\,
            I => \N__21812\
        );

    \I__3934\ : Odrv12
    port map (
            O => \N__21812\,
            I => \b2v_inst.dir_mem_RNO_0Z0Z_6\
        );

    \I__3933\ : InMux
    port map (
            O => \N__21809\,
            I => \N__21806\
        );

    \I__3932\ : LocalMux
    port map (
            O => \N__21806\,
            I => \N__21803\
        );

    \I__3931\ : Span4Mux_h
    port map (
            O => \N__21803\,
            I => \N__21800\
        );

    \I__3930\ : Span4Mux_v
    port map (
            O => \N__21800\,
            I => \N__21797\
        );

    \I__3929\ : Odrv4
    port map (
            O => \N__21797\,
            I => \b2v_inst.dir_memZ0Z_6\
        );

    \I__3928\ : InMux
    port map (
            O => \N__21794\,
            I => \N__21791\
        );

    \I__3927\ : LocalMux
    port map (
            O => \N__21791\,
            I => \N__21788\
        );

    \I__3926\ : Span4Mux_v
    port map (
            O => \N__21788\,
            I => \N__21785\
        );

    \I__3925\ : Span4Mux_h
    port map (
            O => \N__21785\,
            I => \N__21782\
        );

    \I__3924\ : Odrv4
    port map (
            O => \N__21782\,
            I => \b2v_inst.dir_mem_RNO_0Z0Z_8\
        );

    \I__3923\ : InMux
    port map (
            O => \N__21779\,
            I => \N__21776\
        );

    \I__3922\ : LocalMux
    port map (
            O => \N__21776\,
            I => \N__21773\
        );

    \I__3921\ : Span4Mux_v
    port map (
            O => \N__21773\,
            I => \N__21770\
        );

    \I__3920\ : Span4Mux_v
    port map (
            O => \N__21770\,
            I => \N__21767\
        );

    \I__3919\ : Odrv4
    port map (
            O => \N__21767\,
            I => \b2v_inst.dir_memZ0Z_8\
        );

    \I__3918\ : CascadeMux
    port map (
            O => \N__21764\,
            I => \N__21761\
        );

    \I__3917\ : InMux
    port map (
            O => \N__21761\,
            I => \N__21758\
        );

    \I__3916\ : LocalMux
    port map (
            O => \N__21758\,
            I => \N__21755\
        );

    \I__3915\ : Span4Mux_v
    port map (
            O => \N__21755\,
            I => \N__21752\
        );

    \I__3914\ : Span4Mux_h
    port map (
            O => \N__21752\,
            I => \N__21749\
        );

    \I__3913\ : Odrv4
    port map (
            O => \N__21749\,
            I => \b2v_inst.dir_mem_RNO_0Z0Z_9\
        );

    \I__3912\ : InMux
    port map (
            O => \N__21746\,
            I => \N__21743\
        );

    \I__3911\ : LocalMux
    port map (
            O => \N__21743\,
            I => \N__21740\
        );

    \I__3910\ : Odrv12
    port map (
            O => \N__21740\,
            I => \b2v_inst.dir_memZ0Z_9\
        );

    \I__3909\ : InMux
    port map (
            O => \N__21737\,
            I => \N__21734\
        );

    \I__3908\ : LocalMux
    port map (
            O => \N__21734\,
            I => \N__21731\
        );

    \I__3907\ : Span4Mux_v
    port map (
            O => \N__21731\,
            I => \N__21728\
        );

    \I__3906\ : Sp12to4
    port map (
            O => \N__21728\,
            I => \N__21725\
        );

    \I__3905\ : Span12Mux_h
    port map (
            O => \N__21725\,
            I => \N__21722\
        );

    \I__3904\ : Odrv12
    port map (
            O => \N__21722\,
            I => swit_c_4
        );

    \I__3903\ : InMux
    port map (
            O => \N__21719\,
            I => \N__21714\
        );

    \I__3902\ : InMux
    port map (
            O => \N__21718\,
            I => \N__21711\
        );

    \I__3901\ : InMux
    port map (
            O => \N__21717\,
            I => \N__21701\
        );

    \I__3900\ : LocalMux
    port map (
            O => \N__21714\,
            I => \N__21698\
        );

    \I__3899\ : LocalMux
    port map (
            O => \N__21711\,
            I => \N__21695\
        );

    \I__3898\ : InMux
    port map (
            O => \N__21710\,
            I => \N__21692\
        );

    \I__3897\ : InMux
    port map (
            O => \N__21709\,
            I => \N__21687\
        );

    \I__3896\ : InMux
    port map (
            O => \N__21708\,
            I => \N__21687\
        );

    \I__3895\ : InMux
    port map (
            O => \N__21707\,
            I => \N__21678\
        );

    \I__3894\ : InMux
    port map (
            O => \N__21706\,
            I => \N__21678\
        );

    \I__3893\ : InMux
    port map (
            O => \N__21705\,
            I => \N__21678\
        );

    \I__3892\ : InMux
    port map (
            O => \N__21704\,
            I => \N__21678\
        );

    \I__3891\ : LocalMux
    port map (
            O => \N__21701\,
            I => \b2v_inst.N_494\
        );

    \I__3890\ : Odrv12
    port map (
            O => \N__21698\,
            I => \b2v_inst.N_494\
        );

    \I__3889\ : Odrv4
    port map (
            O => \N__21695\,
            I => \b2v_inst.N_494\
        );

    \I__3888\ : LocalMux
    port map (
            O => \N__21692\,
            I => \b2v_inst.N_494\
        );

    \I__3887\ : LocalMux
    port map (
            O => \N__21687\,
            I => \b2v_inst.N_494\
        );

    \I__3886\ : LocalMux
    port map (
            O => \N__21678\,
            I => \b2v_inst.N_494\
        );

    \I__3885\ : InMux
    port map (
            O => \N__21665\,
            I => \N__21655\
        );

    \I__3884\ : InMux
    port map (
            O => \N__21664\,
            I => \N__21655\
        );

    \I__3883\ : InMux
    port map (
            O => \N__21663\,
            I => \N__21655\
        );

    \I__3882\ : InMux
    port map (
            O => \N__21662\,
            I => \N__21651\
        );

    \I__3881\ : LocalMux
    port map (
            O => \N__21655\,
            I => \N__21648\
        );

    \I__3880\ : InMux
    port map (
            O => \N__21654\,
            I => \N__21645\
        );

    \I__3879\ : LocalMux
    port map (
            O => \N__21651\,
            I => \N__21642\
        );

    \I__3878\ : Span4Mux_h
    port map (
            O => \N__21648\,
            I => \N__21637\
        );

    \I__3877\ : LocalMux
    port map (
            O => \N__21645\,
            I => \N__21637\
        );

    \I__3876\ : Span12Mux_h
    port map (
            O => \N__21642\,
            I => \N__21628\
        );

    \I__3875\ : Span4Mux_v
    port map (
            O => \N__21637\,
            I => \N__21625\
        );

    \I__3874\ : InMux
    port map (
            O => \N__21636\,
            I => \N__21622\
        );

    \I__3873\ : InMux
    port map (
            O => \N__21635\,
            I => \N__21619\
        );

    \I__3872\ : InMux
    port map (
            O => \N__21634\,
            I => \N__21610\
        );

    \I__3871\ : InMux
    port map (
            O => \N__21633\,
            I => \N__21610\
        );

    \I__3870\ : InMux
    port map (
            O => \N__21632\,
            I => \N__21610\
        );

    \I__3869\ : InMux
    port map (
            O => \N__21631\,
            I => \N__21610\
        );

    \I__3868\ : Odrv12
    port map (
            O => \N__21628\,
            I => \b2v_inst.N_247\
        );

    \I__3867\ : Odrv4
    port map (
            O => \N__21625\,
            I => \b2v_inst.N_247\
        );

    \I__3866\ : LocalMux
    port map (
            O => \N__21622\,
            I => \b2v_inst.N_247\
        );

    \I__3865\ : LocalMux
    port map (
            O => \N__21619\,
            I => \b2v_inst.N_247\
        );

    \I__3864\ : LocalMux
    port map (
            O => \N__21610\,
            I => \b2v_inst.N_247\
        );

    \I__3863\ : CascadeMux
    port map (
            O => \N__21599\,
            I => \b2v_inst.addr_ram_energia_m0_4_cascade_\
        );

    \I__3862\ : CascadeMux
    port map (
            O => \N__21596\,
            I => \N__21592\
        );

    \I__3861\ : CascadeMux
    port map (
            O => \N__21595\,
            I => \N__21589\
        );

    \I__3860\ : CascadeBuf
    port map (
            O => \N__21592\,
            I => \N__21586\
        );

    \I__3859\ : CascadeBuf
    port map (
            O => \N__21589\,
            I => \N__21583\
        );

    \I__3858\ : CascadeMux
    port map (
            O => \N__21586\,
            I => \N__21580\
        );

    \I__3857\ : CascadeMux
    port map (
            O => \N__21583\,
            I => \N__21577\
        );

    \I__3856\ : CascadeBuf
    port map (
            O => \N__21580\,
            I => \N__21574\
        );

    \I__3855\ : CascadeBuf
    port map (
            O => \N__21577\,
            I => \N__21571\
        );

    \I__3854\ : CascadeMux
    port map (
            O => \N__21574\,
            I => \N__21568\
        );

    \I__3853\ : CascadeMux
    port map (
            O => \N__21571\,
            I => \N__21565\
        );

    \I__3852\ : CascadeBuf
    port map (
            O => \N__21568\,
            I => \N__21562\
        );

    \I__3851\ : CascadeBuf
    port map (
            O => \N__21565\,
            I => \N__21559\
        );

    \I__3850\ : CascadeMux
    port map (
            O => \N__21562\,
            I => \N__21556\
        );

    \I__3849\ : CascadeMux
    port map (
            O => \N__21559\,
            I => \N__21553\
        );

    \I__3848\ : CascadeBuf
    port map (
            O => \N__21556\,
            I => \N__21550\
        );

    \I__3847\ : CascadeBuf
    port map (
            O => \N__21553\,
            I => \N__21547\
        );

    \I__3846\ : CascadeMux
    port map (
            O => \N__21550\,
            I => \N__21544\
        );

    \I__3845\ : CascadeMux
    port map (
            O => \N__21547\,
            I => \N__21541\
        );

    \I__3844\ : CascadeBuf
    port map (
            O => \N__21544\,
            I => \N__21538\
        );

    \I__3843\ : CascadeBuf
    port map (
            O => \N__21541\,
            I => \N__21535\
        );

    \I__3842\ : CascadeMux
    port map (
            O => \N__21538\,
            I => \N__21532\
        );

    \I__3841\ : CascadeMux
    port map (
            O => \N__21535\,
            I => \N__21529\
        );

    \I__3840\ : CascadeBuf
    port map (
            O => \N__21532\,
            I => \N__21526\
        );

    \I__3839\ : CascadeBuf
    port map (
            O => \N__21529\,
            I => \N__21523\
        );

    \I__3838\ : CascadeMux
    port map (
            O => \N__21526\,
            I => \N__21520\
        );

    \I__3837\ : CascadeMux
    port map (
            O => \N__21523\,
            I => \N__21517\
        );

    \I__3836\ : InMux
    port map (
            O => \N__21520\,
            I => \N__21514\
        );

    \I__3835\ : InMux
    port map (
            O => \N__21517\,
            I => \N__21511\
        );

    \I__3834\ : LocalMux
    port map (
            O => \N__21514\,
            I => \N__21506\
        );

    \I__3833\ : LocalMux
    port map (
            O => \N__21511\,
            I => \N__21506\
        );

    \I__3832\ : Span4Mux_v
    port map (
            O => \N__21506\,
            I => \N__21503\
        );

    \I__3831\ : Span4Mux_h
    port map (
            O => \N__21503\,
            I => \N__21500\
        );

    \I__3830\ : Span4Mux_h
    port map (
            O => \N__21500\,
            I => \N__21497\
        );

    \I__3829\ : Odrv4
    port map (
            O => \N__21497\,
            I => \SYNTHESIZED_WIRE_12_4\
        );

    \I__3828\ : InMux
    port map (
            O => \N__21494\,
            I => \N__21491\
        );

    \I__3827\ : LocalMux
    port map (
            O => \N__21491\,
            I => \N__21488\
        );

    \I__3826\ : Span4Mux_h
    port map (
            O => \N__21488\,
            I => \N__21485\
        );

    \I__3825\ : Span4Mux_v
    port map (
            O => \N__21485\,
            I => \N__21482\
        );

    \I__3824\ : Span4Mux_v
    port map (
            O => \N__21482\,
            I => \N__21479\
        );

    \I__3823\ : Odrv4
    port map (
            O => \N__21479\,
            I => uart_rx_i_c
        );

    \I__3822\ : CascadeMux
    port map (
            O => \N__21476\,
            I => \b2v_inst.state18_li_0_cascade_\
        );

    \I__3821\ : CEMux
    port map (
            O => \N__21473\,
            I => \N__21470\
        );

    \I__3820\ : LocalMux
    port map (
            O => \N__21470\,
            I => \N__21464\
        );

    \I__3819\ : CEMux
    port map (
            O => \N__21469\,
            I => \N__21461\
        );

    \I__3818\ : CEMux
    port map (
            O => \N__21468\,
            I => \N__21458\
        );

    \I__3817\ : CEMux
    port map (
            O => \N__21467\,
            I => \N__21450\
        );

    \I__3816\ : Span4Mux_v
    port map (
            O => \N__21464\,
            I => \N__21440\
        );

    \I__3815\ : LocalMux
    port map (
            O => \N__21461\,
            I => \N__21440\
        );

    \I__3814\ : LocalMux
    port map (
            O => \N__21458\,
            I => \N__21440\
        );

    \I__3813\ : CEMux
    port map (
            O => \N__21457\,
            I => \N__21437\
        );

    \I__3812\ : CEMux
    port map (
            O => \N__21456\,
            I => \N__21434\
        );

    \I__3811\ : CEMux
    port map (
            O => \N__21455\,
            I => \N__21431\
        );

    \I__3810\ : CEMux
    port map (
            O => \N__21454\,
            I => \N__21428\
        );

    \I__3809\ : CEMux
    port map (
            O => \N__21453\,
            I => \N__21423\
        );

    \I__3808\ : LocalMux
    port map (
            O => \N__21450\,
            I => \N__21420\
        );

    \I__3807\ : CEMux
    port map (
            O => \N__21449\,
            I => \N__21417\
        );

    \I__3806\ : CEMux
    port map (
            O => \N__21448\,
            I => \N__21414\
        );

    \I__3805\ : CEMux
    port map (
            O => \N__21447\,
            I => \N__21411\
        );

    \I__3804\ : Span4Mux_v
    port map (
            O => \N__21440\,
            I => \N__21403\
        );

    \I__3803\ : LocalMux
    port map (
            O => \N__21437\,
            I => \N__21403\
        );

    \I__3802\ : LocalMux
    port map (
            O => \N__21434\,
            I => \N__21403\
        );

    \I__3801\ : LocalMux
    port map (
            O => \N__21431\,
            I => \N__21398\
        );

    \I__3800\ : LocalMux
    port map (
            O => \N__21428\,
            I => \N__21398\
        );

    \I__3799\ : CEMux
    port map (
            O => \N__21427\,
            I => \N__21395\
        );

    \I__3798\ : CEMux
    port map (
            O => \N__21426\,
            I => \N__21392\
        );

    \I__3797\ : LocalMux
    port map (
            O => \N__21423\,
            I => \N__21388\
        );

    \I__3796\ : Span4Mux_v
    port map (
            O => \N__21420\,
            I => \N__21381\
        );

    \I__3795\ : LocalMux
    port map (
            O => \N__21417\,
            I => \N__21381\
        );

    \I__3794\ : LocalMux
    port map (
            O => \N__21414\,
            I => \N__21381\
        );

    \I__3793\ : LocalMux
    port map (
            O => \N__21411\,
            I => \N__21378\
        );

    \I__3792\ : CEMux
    port map (
            O => \N__21410\,
            I => \N__21375\
        );

    \I__3791\ : Span4Mux_v
    port map (
            O => \N__21403\,
            I => \N__21368\
        );

    \I__3790\ : Span4Mux_v
    port map (
            O => \N__21398\,
            I => \N__21368\
        );

    \I__3789\ : LocalMux
    port map (
            O => \N__21395\,
            I => \N__21368\
        );

    \I__3788\ : LocalMux
    port map (
            O => \N__21392\,
            I => \N__21365\
        );

    \I__3787\ : CEMux
    port map (
            O => \N__21391\,
            I => \N__21362\
        );

    \I__3786\ : Span4Mux_h
    port map (
            O => \N__21388\,
            I => \N__21359\
        );

    \I__3785\ : Span4Mux_v
    port map (
            O => \N__21381\,
            I => \N__21352\
        );

    \I__3784\ : Span4Mux_v
    port map (
            O => \N__21378\,
            I => \N__21352\
        );

    \I__3783\ : LocalMux
    port map (
            O => \N__21375\,
            I => \N__21352\
        );

    \I__3782\ : Span4Mux_v
    port map (
            O => \N__21368\,
            I => \N__21349\
        );

    \I__3781\ : Span4Mux_v
    port map (
            O => \N__21365\,
            I => \N__21344\
        );

    \I__3780\ : LocalMux
    port map (
            O => \N__21362\,
            I => \N__21344\
        );

    \I__3779\ : Span4Mux_h
    port map (
            O => \N__21359\,
            I => \N__21341\
        );

    \I__3778\ : Span4Mux_h
    port map (
            O => \N__21352\,
            I => \N__21338\
        );

    \I__3777\ : Span4Mux_h
    port map (
            O => \N__21349\,
            I => \N__21335\
        );

    \I__3776\ : Span4Mux_h
    port map (
            O => \N__21344\,
            I => \N__21332\
        );

    \I__3775\ : Span4Mux_v
    port map (
            O => \N__21341\,
            I => \N__21327\
        );

    \I__3774\ : Span4Mux_h
    port map (
            O => \N__21338\,
            I => \N__21327\
        );

    \I__3773\ : Span4Mux_h
    port map (
            O => \N__21335\,
            I => \N__21324\
        );

    \I__3772\ : Span4Mux_h
    port map (
            O => \N__21332\,
            I => \N__21319\
        );

    \I__3771\ : Span4Mux_h
    port map (
            O => \N__21327\,
            I => \N__21319\
        );

    \I__3770\ : Odrv4
    port map (
            O => \N__21324\,
            I => \N_130_i\
        );

    \I__3769\ : Odrv4
    port map (
            O => \N__21319\,
            I => \N_130_i\
        );

    \I__3768\ : InMux
    port map (
            O => \N__21314\,
            I => \N__21309\
        );

    \I__3767\ : InMux
    port map (
            O => \N__21313\,
            I => \N__21304\
        );

    \I__3766\ : InMux
    port map (
            O => \N__21312\,
            I => \N__21304\
        );

    \I__3765\ : LocalMux
    port map (
            O => \N__21309\,
            I => \N__21299\
        );

    \I__3764\ : LocalMux
    port map (
            O => \N__21304\,
            I => \N__21296\
        );

    \I__3763\ : CascadeMux
    port map (
            O => \N__21303\,
            I => \N__21293\
        );

    \I__3762\ : CascadeMux
    port map (
            O => \N__21302\,
            I => \N__21290\
        );

    \I__3761\ : Span4Mux_h
    port map (
            O => \N__21299\,
            I => \N__21287\
        );

    \I__3760\ : Span4Mux_h
    port map (
            O => \N__21296\,
            I => \N__21284\
        );

    \I__3759\ : InMux
    port map (
            O => \N__21293\,
            I => \N__21281\
        );

    \I__3758\ : InMux
    port map (
            O => \N__21290\,
            I => \N__21278\
        );

    \I__3757\ : Odrv4
    port map (
            O => \N__21287\,
            I => \b2v_inst.N_512\
        );

    \I__3756\ : Odrv4
    port map (
            O => \N__21284\,
            I => \b2v_inst.N_512\
        );

    \I__3755\ : LocalMux
    port map (
            O => \N__21281\,
            I => \b2v_inst.N_512\
        );

    \I__3754\ : LocalMux
    port map (
            O => \N__21278\,
            I => \b2v_inst.N_512\
        );

    \I__3753\ : InMux
    port map (
            O => \N__21269\,
            I => \N__21266\
        );

    \I__3752\ : LocalMux
    port map (
            O => \N__21266\,
            I => \N__21262\
        );

    \I__3751\ : CascadeMux
    port map (
            O => \N__21265\,
            I => \N__21259\
        );

    \I__3750\ : Span4Mux_v
    port map (
            O => \N__21262\,
            I => \N__21255\
        );

    \I__3749\ : InMux
    port map (
            O => \N__21259\,
            I => \N__21244\
        );

    \I__3748\ : InMux
    port map (
            O => \N__21258\,
            I => \N__21244\
        );

    \I__3747\ : Span4Mux_h
    port map (
            O => \N__21255\,
            I => \N__21241\
        );

    \I__3746\ : InMux
    port map (
            O => \N__21254\,
            I => \N__21236\
        );

    \I__3745\ : InMux
    port map (
            O => \N__21253\,
            I => \N__21236\
        );

    \I__3744\ : InMux
    port map (
            O => \N__21252\,
            I => \N__21229\
        );

    \I__3743\ : InMux
    port map (
            O => \N__21251\,
            I => \N__21229\
        );

    \I__3742\ : InMux
    port map (
            O => \N__21250\,
            I => \N__21229\
        );

    \I__3741\ : InMux
    port map (
            O => \N__21249\,
            I => \N__21226\
        );

    \I__3740\ : LocalMux
    port map (
            O => \N__21244\,
            I => \N__21223\
        );

    \I__3739\ : Span4Mux_h
    port map (
            O => \N__21241\,
            I => \N__21218\
        );

    \I__3738\ : LocalMux
    port map (
            O => \N__21236\,
            I => \N__21218\
        );

    \I__3737\ : LocalMux
    port map (
            O => \N__21229\,
            I => \b2v_inst.stateZ0Z_30\
        );

    \I__3736\ : LocalMux
    port map (
            O => \N__21226\,
            I => \b2v_inst.stateZ0Z_30\
        );

    \I__3735\ : Odrv4
    port map (
            O => \N__21223\,
            I => \b2v_inst.stateZ0Z_30\
        );

    \I__3734\ : Odrv4
    port map (
            O => \N__21218\,
            I => \b2v_inst.stateZ0Z_30\
        );

    \I__3733\ : CascadeMux
    port map (
            O => \N__21209\,
            I => \b2v_inst.N_828_cascade_\
        );

    \I__3732\ : InMux
    port map (
            O => \N__21206\,
            I => \N__21203\
        );

    \I__3731\ : LocalMux
    port map (
            O => \N__21203\,
            I => \N__21200\
        );

    \I__3730\ : Span4Mux_h
    port map (
            O => \N__21200\,
            I => \N__21197\
        );

    \I__3729\ : Span4Mux_h
    port map (
            O => \N__21197\,
            I => \N__21194\
        );

    \I__3728\ : Odrv4
    port map (
            O => \N__21194\,
            I => \N_552_i\
        );

    \I__3727\ : InMux
    port map (
            O => \N__21191\,
            I => \N__21185\
        );

    \I__3726\ : InMux
    port map (
            O => \N__21190\,
            I => \N__21185\
        );

    \I__3725\ : LocalMux
    port map (
            O => \N__21185\,
            I => \N__21182\
        );

    \I__3724\ : Span4Mux_h
    port map (
            O => \N__21182\,
            I => \N__21178\
        );

    \I__3723\ : InMux
    port map (
            O => \N__21181\,
            I => \N__21175\
        );

    \I__3722\ : Odrv4
    port map (
            O => \N__21178\,
            I => \b2v_inst1.N_119\
        );

    \I__3721\ : LocalMux
    port map (
            O => \N__21175\,
            I => \b2v_inst1.N_119\
        );

    \I__3720\ : CascadeMux
    port map (
            O => \N__21170\,
            I => \b2v_inst1.r_Clk_Count_6_iv_0_a3_1_1_1_cascade_\
        );

    \I__3719\ : InMux
    port map (
            O => \N__21167\,
            I => \N__21160\
        );

    \I__3718\ : InMux
    port map (
            O => \N__21166\,
            I => \N__21160\
        );

    \I__3717\ : InMux
    port map (
            O => \N__21165\,
            I => \N__21157\
        );

    \I__3716\ : LocalMux
    port map (
            O => \N__21160\,
            I => \N__21154\
        );

    \I__3715\ : LocalMux
    port map (
            O => \N__21157\,
            I => \N__21151\
        );

    \I__3714\ : Span4Mux_v
    port map (
            O => \N__21154\,
            I => \N__21147\
        );

    \I__3713\ : Span4Mux_h
    port map (
            O => \N__21151\,
            I => \N__21142\
        );

    \I__3712\ : InMux
    port map (
            O => \N__21150\,
            I => \N__21139\
        );

    \I__3711\ : Span4Mux_h
    port map (
            O => \N__21147\,
            I => \N__21136\
        );

    \I__3710\ : InMux
    port map (
            O => \N__21146\,
            I => \N__21131\
        );

    \I__3709\ : InMux
    port map (
            O => \N__21145\,
            I => \N__21131\
        );

    \I__3708\ : Odrv4
    port map (
            O => \N__21142\,
            I => \b2v_inst1.N_43\
        );

    \I__3707\ : LocalMux
    port map (
            O => \N__21139\,
            I => \b2v_inst1.N_43\
        );

    \I__3706\ : Odrv4
    port map (
            O => \N__21136\,
            I => \b2v_inst1.N_43\
        );

    \I__3705\ : LocalMux
    port map (
            O => \N__21131\,
            I => \b2v_inst1.N_43\
        );

    \I__3704\ : CascadeMux
    port map (
            O => \N__21122\,
            I => \b2v_inst1.r_Clk_Count_6_iv_0_0_1_cascade_\
        );

    \I__3703\ : InMux
    port map (
            O => \N__21119\,
            I => \N__21116\
        );

    \I__3702\ : LocalMux
    port map (
            O => \N__21116\,
            I => \N__21113\
        );

    \I__3701\ : Span4Mux_h
    port map (
            O => \N__21113\,
            I => \N__21105\
        );

    \I__3700\ : InMux
    port map (
            O => \N__21112\,
            I => \N__21102\
        );

    \I__3699\ : InMux
    port map (
            O => \N__21111\,
            I => \N__21097\
        );

    \I__3698\ : InMux
    port map (
            O => \N__21110\,
            I => \N__21097\
        );

    \I__3697\ : InMux
    port map (
            O => \N__21109\,
            I => \N__21092\
        );

    \I__3696\ : InMux
    port map (
            O => \N__21108\,
            I => \N__21092\
        );

    \I__3695\ : Odrv4
    port map (
            O => \N__21105\,
            I => \b2v_inst1.r_Clk_CountZ0Z_0\
        );

    \I__3694\ : LocalMux
    port map (
            O => \N__21102\,
            I => \b2v_inst1.r_Clk_CountZ0Z_0\
        );

    \I__3693\ : LocalMux
    port map (
            O => \N__21097\,
            I => \b2v_inst1.r_Clk_CountZ0Z_0\
        );

    \I__3692\ : LocalMux
    port map (
            O => \N__21092\,
            I => \b2v_inst1.r_Clk_CountZ0Z_0\
        );

    \I__3691\ : CascadeMux
    port map (
            O => \N__21083\,
            I => \N__21079\
        );

    \I__3690\ : InMux
    port map (
            O => \N__21082\,
            I => \N__21073\
        );

    \I__3689\ : InMux
    port map (
            O => \N__21079\,
            I => \N__21068\
        );

    \I__3688\ : InMux
    port map (
            O => \N__21078\,
            I => \N__21068\
        );

    \I__3687\ : InMux
    port map (
            O => \N__21077\,
            I => \N__21064\
        );

    \I__3686\ : CascadeMux
    port map (
            O => \N__21076\,
            I => \N__21061\
        );

    \I__3685\ : LocalMux
    port map (
            O => \N__21073\,
            I => \N__21058\
        );

    \I__3684\ : LocalMux
    port map (
            O => \N__21068\,
            I => \N__21055\
        );

    \I__3683\ : InMux
    port map (
            O => \N__21067\,
            I => \N__21052\
        );

    \I__3682\ : LocalMux
    port map (
            O => \N__21064\,
            I => \N__21049\
        );

    \I__3681\ : InMux
    port map (
            O => \N__21061\,
            I => \N__21046\
        );

    \I__3680\ : Span4Mux_h
    port map (
            O => \N__21058\,
            I => \N__21043\
        );

    \I__3679\ : Span4Mux_h
    port map (
            O => \N__21055\,
            I => \N__21040\
        );

    \I__3678\ : LocalMux
    port map (
            O => \N__21052\,
            I => \N__21035\
        );

    \I__3677\ : Span4Mux_h
    port map (
            O => \N__21049\,
            I => \N__21035\
        );

    \I__3676\ : LocalMux
    port map (
            O => \N__21046\,
            I => \b2v_inst1.r_Clk_CountZ0Z_1\
        );

    \I__3675\ : Odrv4
    port map (
            O => \N__21043\,
            I => \b2v_inst1.r_Clk_CountZ0Z_1\
        );

    \I__3674\ : Odrv4
    port map (
            O => \N__21040\,
            I => \b2v_inst1.r_Clk_CountZ0Z_1\
        );

    \I__3673\ : Odrv4
    port map (
            O => \N__21035\,
            I => \b2v_inst1.r_Clk_CountZ0Z_1\
        );

    \I__3672\ : CascadeMux
    port map (
            O => \N__21026\,
            I => \b2v_inst.N_653_cascade_\
        );

    \I__3671\ : CascadeMux
    port map (
            O => \N__21023\,
            I => \N__21019\
        );

    \I__3670\ : InMux
    port map (
            O => \N__21022\,
            I => \N__21011\
        );

    \I__3669\ : InMux
    port map (
            O => \N__21019\,
            I => \N__21011\
        );

    \I__3668\ : InMux
    port map (
            O => \N__21018\,
            I => \N__21011\
        );

    \I__3667\ : LocalMux
    port map (
            O => \N__21011\,
            I => \b2v_inst.stateZ0Z_17\
        );

    \I__3666\ : InMux
    port map (
            O => \N__21008\,
            I => \N__21005\
        );

    \I__3665\ : LocalMux
    port map (
            O => \N__21005\,
            I => \b2v_inst.state_ns_i_a2_1_15\
        );

    \I__3664\ : CascadeMux
    port map (
            O => \N__21002\,
            I => \b2v_inst.cuenta_RNIKUJVZ0Z_0_cascade_\
        );

    \I__3663\ : CascadeMux
    port map (
            O => \N__20999\,
            I => \b2v_inst.un20_cuentalto10_5_cascade_\
        );

    \I__3662\ : InMux
    port map (
            O => \N__20996\,
            I => \N__20993\
        );

    \I__3661\ : LocalMux
    port map (
            O => \N__20993\,
            I => \b2v_inst.un20_cuentalto10_sx\
        );

    \I__3660\ : CascadeMux
    port map (
            O => \N__20990\,
            I => \b2v_inst.un20_cuentalto10_sx_cascade_\
        );

    \I__3659\ : InMux
    port map (
            O => \N__20987\,
            I => \N__20983\
        );

    \I__3658\ : InMux
    port map (
            O => \N__20986\,
            I => \N__20980\
        );

    \I__3657\ : LocalMux
    port map (
            O => \N__20983\,
            I => \b2v_inst.N_829\
        );

    \I__3656\ : LocalMux
    port map (
            O => \N__20980\,
            I => \b2v_inst.N_829\
        );

    \I__3655\ : CascadeMux
    port map (
            O => \N__20975\,
            I => \b2v_inst.un1_state_23_i_a2_0_a2_0_a2_0_cascade_\
        );

    \I__3654\ : InMux
    port map (
            O => \N__20972\,
            I => \N__20969\
        );

    \I__3653\ : LocalMux
    port map (
            O => \N__20969\,
            I => \N__20965\
        );

    \I__3652\ : InMux
    port map (
            O => \N__20968\,
            I => \N__20961\
        );

    \I__3651\ : Span4Mux_h
    port map (
            O => \N__20965\,
            I => \N__20958\
        );

    \I__3650\ : InMux
    port map (
            O => \N__20964\,
            I => \N__20955\
        );

    \I__3649\ : LocalMux
    port map (
            O => \N__20961\,
            I => \b2v_inst.stateZ0Z_22\
        );

    \I__3648\ : Odrv4
    port map (
            O => \N__20958\,
            I => \b2v_inst.stateZ0Z_22\
        );

    \I__3647\ : LocalMux
    port map (
            O => \N__20955\,
            I => \b2v_inst.stateZ0Z_22\
        );

    \I__3646\ : InMux
    port map (
            O => \N__20948\,
            I => \N__20943\
        );

    \I__3645\ : InMux
    port map (
            O => \N__20947\,
            I => \N__20939\
        );

    \I__3644\ : InMux
    port map (
            O => \N__20946\,
            I => \N__20936\
        );

    \I__3643\ : LocalMux
    port map (
            O => \N__20943\,
            I => \N__20933\
        );

    \I__3642\ : InMux
    port map (
            O => \N__20942\,
            I => \N__20930\
        );

    \I__3641\ : LocalMux
    port map (
            O => \N__20939\,
            I => \N__20927\
        );

    \I__3640\ : LocalMux
    port map (
            O => \N__20936\,
            I => \b2v_inst.stateZ0Z_26\
        );

    \I__3639\ : Odrv4
    port map (
            O => \N__20933\,
            I => \b2v_inst.stateZ0Z_26\
        );

    \I__3638\ : LocalMux
    port map (
            O => \N__20930\,
            I => \b2v_inst.stateZ0Z_26\
        );

    \I__3637\ : Odrv4
    port map (
            O => \N__20927\,
            I => \b2v_inst.stateZ0Z_26\
        );

    \I__3636\ : InMux
    port map (
            O => \N__20918\,
            I => \N__20915\
        );

    \I__3635\ : LocalMux
    port map (
            O => \N__20915\,
            I => \b2v_inst.un2_cuentalto10_i_a2_6\
        );

    \I__3634\ : InMux
    port map (
            O => \N__20912\,
            I => \N__20909\
        );

    \I__3633\ : LocalMux
    port map (
            O => \N__20909\,
            I => \N__20906\
        );

    \I__3632\ : Span4Mux_v
    port map (
            O => \N__20906\,
            I => \N__20903\
        );

    \I__3631\ : Span4Mux_h
    port map (
            O => \N__20903\,
            I => \N__20899\
        );

    \I__3630\ : InMux
    port map (
            O => \N__20902\,
            I => \N__20896\
        );

    \I__3629\ : Odrv4
    port map (
            O => \N__20899\,
            I => \b2v_inst1.m16_0_o2\
        );

    \I__3628\ : LocalMux
    port map (
            O => \N__20896\,
            I => \b2v_inst1.m16_0_o2\
        );

    \I__3627\ : CascadeMux
    port map (
            O => \N__20891\,
            I => \b2v_inst1.m16_0_a3_0_cascade_\
        );

    \I__3626\ : InMux
    port map (
            O => \N__20888\,
            I => \N__20885\
        );

    \I__3625\ : LocalMux
    port map (
            O => \N__20885\,
            I => \N__20882\
        );

    \I__3624\ : Span4Mux_h
    port map (
            O => \N__20882\,
            I => \N__20879\
        );

    \I__3623\ : Odrv4
    port map (
            O => \N__20879\,
            I => \b2v_inst.dir_mem_1Z0Z_9\
        );

    \I__3622\ : CascadeMux
    port map (
            O => \N__20876\,
            I => \N__20873\
        );

    \I__3621\ : InMux
    port map (
            O => \N__20873\,
            I => \N__20870\
        );

    \I__3620\ : LocalMux
    port map (
            O => \N__20870\,
            I => \N__20867\
        );

    \I__3619\ : Span4Mux_v
    port map (
            O => \N__20867\,
            I => \N__20864\
        );

    \I__3618\ : Span4Mux_h
    port map (
            O => \N__20864\,
            I => \N__20861\
        );

    \I__3617\ : Odrv4
    port map (
            O => \N__20861\,
            I => \b2v_inst.dir_mem_3Z0Z_9\
        );

    \I__3616\ : InMux
    port map (
            O => \N__20858\,
            I => \N__20855\
        );

    \I__3615\ : LocalMux
    port map (
            O => \N__20855\,
            I => \N__20852\
        );

    \I__3614\ : Span4Mux_h
    port map (
            O => \N__20852\,
            I => \N__20849\
        );

    \I__3613\ : Span4Mux_h
    port map (
            O => \N__20849\,
            I => \N__20846\
        );

    \I__3612\ : Odrv4
    port map (
            O => \N__20846\,
            I => \N_554_i\
        );

    \I__3611\ : InMux
    port map (
            O => \N__20843\,
            I => \N__20840\
        );

    \I__3610\ : LocalMux
    port map (
            O => \N__20840\,
            I => \N__20837\
        );

    \I__3609\ : Span4Mux_v
    port map (
            O => \N__20837\,
            I => \N__20834\
        );

    \I__3608\ : Span4Mux_h
    port map (
            O => \N__20834\,
            I => \N__20831\
        );

    \I__3607\ : Odrv4
    port map (
            O => \N__20831\,
            I => \b2v_inst.dir_mem_2Z0Z_2\
        );

    \I__3606\ : CascadeMux
    port map (
            O => \N__20828\,
            I => \N__20825\
        );

    \I__3605\ : InMux
    port map (
            O => \N__20825\,
            I => \N__20822\
        );

    \I__3604\ : LocalMux
    port map (
            O => \N__20822\,
            I => \N__20819\
        );

    \I__3603\ : Odrv12
    port map (
            O => \N__20819\,
            I => \b2v_inst.dir_memZ0Z_2\
        );

    \I__3602\ : CascadeMux
    port map (
            O => \N__20816\,
            I => \N__20813\
        );

    \I__3601\ : InMux
    port map (
            O => \N__20813\,
            I => \N__20810\
        );

    \I__3600\ : LocalMux
    port map (
            O => \N__20810\,
            I => \N__20807\
        );

    \I__3599\ : Odrv4
    port map (
            O => \N__20807\,
            I => \b2v_inst.dir_mem_2Z0Z_9\
        );

    \I__3598\ : InMux
    port map (
            O => \N__20804\,
            I => \N__20801\
        );

    \I__3597\ : LocalMux
    port map (
            O => \N__20801\,
            I => \b2v_inst.dir_mem_1Z0Z_2\
        );

    \I__3596\ : CascadeMux
    port map (
            O => \N__20798\,
            I => \N__20795\
        );

    \I__3595\ : InMux
    port map (
            O => \N__20795\,
            I => \N__20792\
        );

    \I__3594\ : LocalMux
    port map (
            O => \N__20792\,
            I => \N__20789\
        );

    \I__3593\ : Odrv12
    port map (
            O => \N__20789\,
            I => \b2v_inst.dir_mem_3Z0Z_2\
        );

    \I__3592\ : CascadeMux
    port map (
            O => \N__20786\,
            I => \b2v_inst.N_829_cascade_\
        );

    \I__3591\ : InMux
    port map (
            O => \N__20783\,
            I => \N__20780\
        );

    \I__3590\ : LocalMux
    port map (
            O => \N__20780\,
            I => \N__20776\
        );

    \I__3589\ : CascadeMux
    port map (
            O => \N__20779\,
            I => \N__20773\
        );

    \I__3588\ : Span4Mux_v
    port map (
            O => \N__20776\,
            I => \N__20770\
        );

    \I__3587\ : InMux
    port map (
            O => \N__20773\,
            I => \N__20767\
        );

    \I__3586\ : Span4Mux_h
    port map (
            O => \N__20770\,
            I => \N__20764\
        );

    \I__3585\ : LocalMux
    port map (
            O => \N__20767\,
            I => \N__20761\
        );

    \I__3584\ : Odrv4
    port map (
            O => \N__20764\,
            I => \b2v_inst.dir_mem_215lto7\
        );

    \I__3583\ : Odrv4
    port map (
            O => \N__20761\,
            I => \b2v_inst.dir_mem_215lto7\
        );

    \I__3582\ : InMux
    port map (
            O => \N__20756\,
            I => \N__20753\
        );

    \I__3581\ : LocalMux
    port map (
            O => \N__20753\,
            I => \N__20750\
        );

    \I__3580\ : Span4Mux_v
    port map (
            O => \N__20750\,
            I => \N__20747\
        );

    \I__3579\ : Span4Mux_h
    port map (
            O => \N__20747\,
            I => \N__20744\
        );

    \I__3578\ : Odrv4
    port map (
            O => \N__20744\,
            I => \b2v_inst.dir_mem_2Z0Z_7\
        );

    \I__3577\ : InMux
    port map (
            O => \N__20741\,
            I => \N__20738\
        );

    \I__3576\ : LocalMux
    port map (
            O => \N__20738\,
            I => \N__20735\
        );

    \I__3575\ : Span4Mux_v
    port map (
            O => \N__20735\,
            I => \N__20731\
        );

    \I__3574\ : InMux
    port map (
            O => \N__20734\,
            I => \N__20728\
        );

    \I__3573\ : Odrv4
    port map (
            O => \N__20731\,
            I => \b2v_inst.un8_dir_mem_2_cry_6_c_RNIINQZ0Z5\
        );

    \I__3572\ : LocalMux
    port map (
            O => \N__20728\,
            I => \b2v_inst.un8_dir_mem_2_cry_6_c_RNIINQZ0Z5\
        );

    \I__3571\ : CascadeMux
    port map (
            O => \N__20723\,
            I => \N__20720\
        );

    \I__3570\ : InMux
    port map (
            O => \N__20720\,
            I => \N__20717\
        );

    \I__3569\ : LocalMux
    port map (
            O => \N__20717\,
            I => \N__20714\
        );

    \I__3568\ : Span4Mux_v
    port map (
            O => \N__20714\,
            I => \N__20711\
        );

    \I__3567\ : Odrv4
    port map (
            O => \N__20711\,
            I => \b2v_inst.dir_mem_2Z0Z_8\
        );

    \I__3566\ : InMux
    port map (
            O => \N__20708\,
            I => \N__20705\
        );

    \I__3565\ : LocalMux
    port map (
            O => \N__20705\,
            I => \N__20702\
        );

    \I__3564\ : Span4Mux_h
    port map (
            O => \N__20702\,
            I => \N__20698\
        );

    \I__3563\ : InMux
    port map (
            O => \N__20701\,
            I => \N__20695\
        );

    \I__3562\ : Odrv4
    port map (
            O => \N__20698\,
            I => \b2v_inst.un8_dir_mem_2_cry_7_c_RNIKQRZ0Z5\
        );

    \I__3561\ : LocalMux
    port map (
            O => \N__20695\,
            I => \b2v_inst.un8_dir_mem_2_cry_7_c_RNIKQRZ0Z5\
        );

    \I__3560\ : CascadeMux
    port map (
            O => \N__20690\,
            I => \N__20686\
        );

    \I__3559\ : InMux
    port map (
            O => \N__20689\,
            I => \N__20672\
        );

    \I__3558\ : InMux
    port map (
            O => \N__20686\,
            I => \N__20672\
        );

    \I__3557\ : InMux
    port map (
            O => \N__20685\,
            I => \N__20672\
        );

    \I__3556\ : InMux
    port map (
            O => \N__20684\,
            I => \N__20659\
        );

    \I__3555\ : InMux
    port map (
            O => \N__20683\,
            I => \N__20659\
        );

    \I__3554\ : InMux
    port map (
            O => \N__20682\,
            I => \N__20659\
        );

    \I__3553\ : InMux
    port map (
            O => \N__20681\,
            I => \N__20659\
        );

    \I__3552\ : InMux
    port map (
            O => \N__20680\,
            I => \N__20659\
        );

    \I__3551\ : InMux
    port map (
            O => \N__20679\,
            I => \N__20659\
        );

    \I__3550\ : LocalMux
    port map (
            O => \N__20672\,
            I => \N__20656\
        );

    \I__3549\ : LocalMux
    port map (
            O => \N__20659\,
            I => \N__20653\
        );

    \I__3548\ : Odrv12
    port map (
            O => \N__20656\,
            I => \b2v_inst.dir_mem_215lto11_0\
        );

    \I__3547\ : Odrv4
    port map (
            O => \N__20653\,
            I => \b2v_inst.dir_mem_215lto11_0\
        );

    \I__3546\ : InMux
    port map (
            O => \N__20648\,
            I => \N__20627\
        );

    \I__3545\ : InMux
    port map (
            O => \N__20647\,
            I => \N__20627\
        );

    \I__3544\ : InMux
    port map (
            O => \N__20646\,
            I => \N__20627\
        );

    \I__3543\ : InMux
    port map (
            O => \N__20645\,
            I => \N__20627\
        );

    \I__3542\ : InMux
    port map (
            O => \N__20644\,
            I => \N__20627\
        );

    \I__3541\ : InMux
    port map (
            O => \N__20643\,
            I => \N__20614\
        );

    \I__3540\ : InMux
    port map (
            O => \N__20642\,
            I => \N__20614\
        );

    \I__3539\ : InMux
    port map (
            O => \N__20641\,
            I => \N__20614\
        );

    \I__3538\ : InMux
    port map (
            O => \N__20640\,
            I => \N__20614\
        );

    \I__3537\ : InMux
    port map (
            O => \N__20639\,
            I => \N__20614\
        );

    \I__3536\ : InMux
    port map (
            O => \N__20638\,
            I => \N__20614\
        );

    \I__3535\ : LocalMux
    port map (
            O => \N__20627\,
            I => \N__20611\
        );

    \I__3534\ : LocalMux
    port map (
            O => \N__20614\,
            I => \b2v_inst.dir_mem_215lt11\
        );

    \I__3533\ : Odrv4
    port map (
            O => \N__20611\,
            I => \b2v_inst.dir_mem_215lt11\
        );

    \I__3532\ : CEMux
    port map (
            O => \N__20606\,
            I => \N__20603\
        );

    \I__3531\ : LocalMux
    port map (
            O => \N__20603\,
            I => \N__20599\
        );

    \I__3530\ : CEMux
    port map (
            O => \N__20602\,
            I => \N__20596\
        );

    \I__3529\ : Odrv4
    port map (
            O => \N__20599\,
            I => \b2v_inst.N_463_i\
        );

    \I__3528\ : LocalMux
    port map (
            O => \N__20596\,
            I => \b2v_inst.N_463_i\
        );

    \I__3527\ : InMux
    port map (
            O => \N__20591\,
            I => \N__20588\
        );

    \I__3526\ : LocalMux
    port map (
            O => \N__20588\,
            I => \N__20585\
        );

    \I__3525\ : Odrv12
    port map (
            O => \N__20585\,
            I => \b2v_inst.indice_4_i_a2_0_7_3_1\
        );

    \I__3524\ : InMux
    port map (
            O => \N__20582\,
            I => \N__20579\
        );

    \I__3523\ : LocalMux
    port map (
            O => \N__20579\,
            I => \b2v_inst.N_432_1_tz\
        );

    \I__3522\ : InMux
    port map (
            O => \N__20576\,
            I => \N__20573\
        );

    \I__3521\ : LocalMux
    port map (
            O => \N__20573\,
            I => \N__20570\
        );

    \I__3520\ : Span4Mux_h
    port map (
            O => \N__20570\,
            I => \N__20567\
        );

    \I__3519\ : Span4Mux_h
    port map (
            O => \N__20567\,
            I => \N__20564\
        );

    \I__3518\ : Odrv4
    port map (
            O => \N__20564\,
            I => \N_556_i\
        );

    \I__3517\ : InMux
    port map (
            O => \N__20561\,
            I => \N__20558\
        );

    \I__3516\ : LocalMux
    port map (
            O => \N__20558\,
            I => \b2v_inst.indice_4_i_a2_0_7_2_1\
        );

    \I__3515\ : InMux
    port map (
            O => \N__20555\,
            I => \N__20552\
        );

    \I__3514\ : LocalMux
    port map (
            O => \N__20552\,
            I => \N__20549\
        );

    \I__3513\ : Span4Mux_h
    port map (
            O => \N__20549\,
            I => \N__20546\
        );

    \I__3512\ : Span4Mux_v
    port map (
            O => \N__20546\,
            I => \N__20543\
        );

    \I__3511\ : Span4Mux_h
    port map (
            O => \N__20543\,
            I => \N__20540\
        );

    \I__3510\ : Odrv4
    port map (
            O => \N__20540\,
            I => \N_117_i\
        );

    \I__3509\ : CascadeMux
    port map (
            O => \N__20537\,
            I => \b2v_inst.addr_ram_energia_m0_3_cascade_\
        );

    \I__3508\ : CascadeMux
    port map (
            O => \N__20534\,
            I => \N__20530\
        );

    \I__3507\ : CascadeMux
    port map (
            O => \N__20533\,
            I => \N__20527\
        );

    \I__3506\ : CascadeBuf
    port map (
            O => \N__20530\,
            I => \N__20524\
        );

    \I__3505\ : CascadeBuf
    port map (
            O => \N__20527\,
            I => \N__20521\
        );

    \I__3504\ : CascadeMux
    port map (
            O => \N__20524\,
            I => \N__20518\
        );

    \I__3503\ : CascadeMux
    port map (
            O => \N__20521\,
            I => \N__20515\
        );

    \I__3502\ : CascadeBuf
    port map (
            O => \N__20518\,
            I => \N__20512\
        );

    \I__3501\ : CascadeBuf
    port map (
            O => \N__20515\,
            I => \N__20509\
        );

    \I__3500\ : CascadeMux
    port map (
            O => \N__20512\,
            I => \N__20506\
        );

    \I__3499\ : CascadeMux
    port map (
            O => \N__20509\,
            I => \N__20503\
        );

    \I__3498\ : CascadeBuf
    port map (
            O => \N__20506\,
            I => \N__20500\
        );

    \I__3497\ : CascadeBuf
    port map (
            O => \N__20503\,
            I => \N__20497\
        );

    \I__3496\ : CascadeMux
    port map (
            O => \N__20500\,
            I => \N__20494\
        );

    \I__3495\ : CascadeMux
    port map (
            O => \N__20497\,
            I => \N__20491\
        );

    \I__3494\ : CascadeBuf
    port map (
            O => \N__20494\,
            I => \N__20488\
        );

    \I__3493\ : CascadeBuf
    port map (
            O => \N__20491\,
            I => \N__20485\
        );

    \I__3492\ : CascadeMux
    port map (
            O => \N__20488\,
            I => \N__20482\
        );

    \I__3491\ : CascadeMux
    port map (
            O => \N__20485\,
            I => \N__20479\
        );

    \I__3490\ : CascadeBuf
    port map (
            O => \N__20482\,
            I => \N__20476\
        );

    \I__3489\ : CascadeBuf
    port map (
            O => \N__20479\,
            I => \N__20473\
        );

    \I__3488\ : CascadeMux
    port map (
            O => \N__20476\,
            I => \N__20470\
        );

    \I__3487\ : CascadeMux
    port map (
            O => \N__20473\,
            I => \N__20467\
        );

    \I__3486\ : CascadeBuf
    port map (
            O => \N__20470\,
            I => \N__20464\
        );

    \I__3485\ : CascadeBuf
    port map (
            O => \N__20467\,
            I => \N__20461\
        );

    \I__3484\ : CascadeMux
    port map (
            O => \N__20464\,
            I => \N__20458\
        );

    \I__3483\ : CascadeMux
    port map (
            O => \N__20461\,
            I => \N__20455\
        );

    \I__3482\ : InMux
    port map (
            O => \N__20458\,
            I => \N__20452\
        );

    \I__3481\ : InMux
    port map (
            O => \N__20455\,
            I => \N__20449\
        );

    \I__3480\ : LocalMux
    port map (
            O => \N__20452\,
            I => \N__20444\
        );

    \I__3479\ : LocalMux
    port map (
            O => \N__20449\,
            I => \N__20444\
        );

    \I__3478\ : Span4Mux_v
    port map (
            O => \N__20444\,
            I => \N__20441\
        );

    \I__3477\ : Span4Mux_h
    port map (
            O => \N__20441\,
            I => \N__20438\
        );

    \I__3476\ : Span4Mux_h
    port map (
            O => \N__20438\,
            I => \N__20435\
        );

    \I__3475\ : Odrv4
    port map (
            O => \N__20435\,
            I => \SYNTHESIZED_WIRE_12_3\
        );

    \I__3474\ : IoInMux
    port map (
            O => \N__20432\,
            I => \N__20429\
        );

    \I__3473\ : LocalMux
    port map (
            O => \N__20429\,
            I => \N__20426\
        );

    \I__3472\ : Span4Mux_s3_h
    port map (
            O => \N__20426\,
            I => \N__20422\
        );

    \I__3471\ : InMux
    port map (
            O => \N__20425\,
            I => \N__20419\
        );

    \I__3470\ : Span4Mux_v
    port map (
            O => \N__20422\,
            I => \N__20416\
        );

    \I__3469\ : LocalMux
    port map (
            O => \N__20419\,
            I => \N__20413\
        );

    \I__3468\ : Span4Mux_h
    port map (
            O => \N__20416\,
            I => \N__20410\
        );

    \I__3467\ : Span4Mux_h
    port map (
            O => \N__20413\,
            I => \N__20407\
        );

    \I__3466\ : Sp12to4
    port map (
            O => \N__20410\,
            I => \N__20404\
        );

    \I__3465\ : Span4Mux_h
    port map (
            O => \N__20407\,
            I => \N__20401\
        );

    \I__3464\ : Odrv12
    port map (
            O => \N__20404\,
            I => leds_c_6
        );

    \I__3463\ : Odrv4
    port map (
            O => \N__20401\,
            I => leds_c_6
        );

    \I__3462\ : InMux
    port map (
            O => \N__20396\,
            I => \N__20393\
        );

    \I__3461\ : LocalMux
    port map (
            O => \N__20393\,
            I => \N__20390\
        );

    \I__3460\ : Sp12to4
    port map (
            O => \N__20390\,
            I => \N__20387\
        );

    \I__3459\ : Odrv12
    port map (
            O => \N__20387\,
            I => swit_c_0
        );

    \I__3458\ : CascadeMux
    port map (
            O => \N__20384\,
            I => \N__20381\
        );

    \I__3457\ : InMux
    port map (
            O => \N__20381\,
            I => \N__20378\
        );

    \I__3456\ : LocalMux
    port map (
            O => \N__20378\,
            I => \N__20375\
        );

    \I__3455\ : Odrv12
    port map (
            O => \N__20375\,
            I => \b2v_inst.addr_ram_energia_m0_0\
        );

    \I__3454\ : InMux
    port map (
            O => \N__20372\,
            I => \N__20369\
        );

    \I__3453\ : LocalMux
    port map (
            O => \N__20369\,
            I => \N__20366\
        );

    \I__3452\ : Span4Mux_v
    port map (
            O => \N__20366\,
            I => \N__20363\
        );

    \I__3451\ : Sp12to4
    port map (
            O => \N__20363\,
            I => \N__20360\
        );

    \I__3450\ : Odrv12
    port map (
            O => \N__20360\,
            I => \N_120_i\
        );

    \I__3449\ : CascadeMux
    port map (
            O => \N__20357\,
            I => \b2v_inst.N_432_1_cascade_\
        );

    \I__3448\ : InMux
    port map (
            O => \N__20354\,
            I => \N__20351\
        );

    \I__3447\ : LocalMux
    port map (
            O => \N__20351\,
            I => \N__20346\
        );

    \I__3446\ : InMux
    port map (
            O => \N__20350\,
            I => \N__20341\
        );

    \I__3445\ : InMux
    port map (
            O => \N__20349\,
            I => \N__20341\
        );

    \I__3444\ : Span4Mux_h
    port map (
            O => \N__20346\,
            I => \N__20338\
        );

    \I__3443\ : LocalMux
    port map (
            O => \N__20341\,
            I => \N__20334\
        );

    \I__3442\ : Span4Mux_h
    port map (
            O => \N__20338\,
            I => \N__20331\
        );

    \I__3441\ : InMux
    port map (
            O => \N__20337\,
            I => \N__20328\
        );

    \I__3440\ : Odrv4
    port map (
            O => \N__20334\,
            I => \b2v_inst.un1_indice_cry_9_c_RNILAJPZ0\
        );

    \I__3439\ : Odrv4
    port map (
            O => \N__20331\,
            I => \b2v_inst.un1_indice_cry_9_c_RNILAJPZ0\
        );

    \I__3438\ : LocalMux
    port map (
            O => \N__20328\,
            I => \b2v_inst.un1_indice_cry_9_c_RNILAJPZ0\
        );

    \I__3437\ : InMux
    port map (
            O => \N__20321\,
            I => \N__20317\
        );

    \I__3436\ : InMux
    port map (
            O => \N__20320\,
            I => \N__20314\
        );

    \I__3435\ : LocalMux
    port map (
            O => \N__20317\,
            I => \N__20311\
        );

    \I__3434\ : LocalMux
    port map (
            O => \N__20314\,
            I => \N__20307\
        );

    \I__3433\ : Span4Mux_h
    port map (
            O => \N__20311\,
            I => \N__20304\
        );

    \I__3432\ : InMux
    port map (
            O => \N__20310\,
            I => \N__20301\
        );

    \I__3431\ : Span4Mux_h
    port map (
            O => \N__20307\,
            I => \N__20298\
        );

    \I__3430\ : Span4Mux_h
    port map (
            O => \N__20304\,
            I => \N__20293\
        );

    \I__3429\ : LocalMux
    port map (
            O => \N__20301\,
            I => \N__20293\
        );

    \I__3428\ : Odrv4
    port map (
            O => \N__20298\,
            I => \b2v_inst.un1_indice_cry_7_c_RNIAFQGZ0\
        );

    \I__3427\ : Odrv4
    port map (
            O => \N__20293\,
            I => \b2v_inst.un1_indice_cry_7_c_RNIAFQGZ0\
        );

    \I__3426\ : CascadeMux
    port map (
            O => \N__20288\,
            I => \N__20285\
        );

    \I__3425\ : InMux
    port map (
            O => \N__20285\,
            I => \N__20282\
        );

    \I__3424\ : LocalMux
    port map (
            O => \N__20282\,
            I => \N__20279\
        );

    \I__3423\ : Span4Mux_h
    port map (
            O => \N__20279\,
            I => \N__20276\
        );

    \I__3422\ : Span4Mux_v
    port map (
            O => \N__20276\,
            I => \N__20273\
        );

    \I__3421\ : Odrv4
    port map (
            O => \N__20273\,
            I => \b2v_inst.dir_mem_2Z0Z_0\
        );

    \I__3420\ : CascadeMux
    port map (
            O => \N__20270\,
            I => \N__20266\
        );

    \I__3419\ : InMux
    port map (
            O => \N__20269\,
            I => \N__20261\
        );

    \I__3418\ : InMux
    port map (
            O => \N__20266\,
            I => \N__20261\
        );

    \I__3417\ : LocalMux
    port map (
            O => \N__20261\,
            I => \N__20257\
        );

    \I__3416\ : InMux
    port map (
            O => \N__20260\,
            I => \N__20254\
        );

    \I__3415\ : Odrv4
    port map (
            O => \N__20257\,
            I => \b2v_inst.un8_dir_mem_2_cry_9_THRU_CO\
        );

    \I__3414\ : LocalMux
    port map (
            O => \N__20254\,
            I => \b2v_inst.un8_dir_mem_2_cry_9_THRU_CO\
        );

    \I__3413\ : InMux
    port map (
            O => \N__20249\,
            I => \N__20245\
        );

    \I__3412\ : InMux
    port map (
            O => \N__20248\,
            I => \N__20242\
        );

    \I__3411\ : LocalMux
    port map (
            O => \N__20245\,
            I => \N__20236\
        );

    \I__3410\ : LocalMux
    port map (
            O => \N__20242\,
            I => \N__20236\
        );

    \I__3409\ : InMux
    port map (
            O => \N__20241\,
            I => \N__20233\
        );

    \I__3408\ : Odrv4
    port map (
            O => \N__20236\,
            I => \b2v_inst.un8_dir_mem_2_cry_8_c_RNITIJEZ0\
        );

    \I__3407\ : LocalMux
    port map (
            O => \N__20233\,
            I => \b2v_inst.un8_dir_mem_2_cry_8_c_RNITIJEZ0\
        );

    \I__3406\ : CascadeMux
    port map (
            O => \N__20228\,
            I => \N__20225\
        );

    \I__3405\ : InMux
    port map (
            O => \N__20225\,
            I => \N__20222\
        );

    \I__3404\ : LocalMux
    port map (
            O => \N__20222\,
            I => \N__20219\
        );

    \I__3403\ : Span4Mux_v
    port map (
            O => \N__20219\,
            I => \N__20216\
        );

    \I__3402\ : Odrv4
    port map (
            O => \N__20216\,
            I => \b2v_inst.dir_mem_2Z0Z_10\
        );

    \I__3401\ : InMux
    port map (
            O => \N__20213\,
            I => \N__20205\
        );

    \I__3400\ : InMux
    port map (
            O => \N__20212\,
            I => \N__20205\
        );

    \I__3399\ : InMux
    port map (
            O => \N__20211\,
            I => \N__20200\
        );

    \I__3398\ : InMux
    port map (
            O => \N__20210\,
            I => \N__20200\
        );

    \I__3397\ : LocalMux
    port map (
            O => \N__20205\,
            I => \b2v_inst.N_477\
        );

    \I__3396\ : LocalMux
    port map (
            O => \N__20200\,
            I => \b2v_inst.N_477\
        );

    \I__3395\ : InMux
    port map (
            O => \N__20195\,
            I => \N__20192\
        );

    \I__3394\ : LocalMux
    port map (
            O => \N__20192\,
            I => \N__20189\
        );

    \I__3393\ : Span4Mux_v
    port map (
            O => \N__20189\,
            I => \N__20186\
        );

    \I__3392\ : Span4Mux_v
    port map (
            O => \N__20186\,
            I => \N__20183\
        );

    \I__3391\ : Span4Mux_v
    port map (
            O => \N__20183\,
            I => \N__20180\
        );

    \I__3390\ : Sp12to4
    port map (
            O => \N__20180\,
            I => \N__20177\
        );

    \I__3389\ : Span12Mux_h
    port map (
            O => \N__20177\,
            I => \N__20174\
        );

    \I__3388\ : Odrv12
    port map (
            O => \N__20174\,
            I => swit_c_1
        );

    \I__3387\ : CascadeMux
    port map (
            O => \N__20171\,
            I => \b2v_inst.N_494_cascade_\
        );

    \I__3386\ : CascadeMux
    port map (
            O => \N__20168\,
            I => \N__20165\
        );

    \I__3385\ : InMux
    port map (
            O => \N__20165\,
            I => \N__20162\
        );

    \I__3384\ : LocalMux
    port map (
            O => \N__20162\,
            I => \N__20159\
        );

    \I__3383\ : Span4Mux_v
    port map (
            O => \N__20159\,
            I => \N__20156\
        );

    \I__3382\ : Span4Mux_h
    port map (
            O => \N__20156\,
            I => \N__20153\
        );

    \I__3381\ : Odrv4
    port map (
            O => \N__20153\,
            I => \b2v_inst.addr_ram_energia_m0_1\
        );

    \I__3380\ : CascadeMux
    port map (
            O => \N__20150\,
            I => \N__20146\
        );

    \I__3379\ : CascadeMux
    port map (
            O => \N__20149\,
            I => \N__20143\
        );

    \I__3378\ : CascadeBuf
    port map (
            O => \N__20146\,
            I => \N__20140\
        );

    \I__3377\ : CascadeBuf
    port map (
            O => \N__20143\,
            I => \N__20137\
        );

    \I__3376\ : CascadeMux
    port map (
            O => \N__20140\,
            I => \N__20134\
        );

    \I__3375\ : CascadeMux
    port map (
            O => \N__20137\,
            I => \N__20131\
        );

    \I__3374\ : CascadeBuf
    port map (
            O => \N__20134\,
            I => \N__20128\
        );

    \I__3373\ : CascadeBuf
    port map (
            O => \N__20131\,
            I => \N__20125\
        );

    \I__3372\ : CascadeMux
    port map (
            O => \N__20128\,
            I => \N__20122\
        );

    \I__3371\ : CascadeMux
    port map (
            O => \N__20125\,
            I => \N__20119\
        );

    \I__3370\ : CascadeBuf
    port map (
            O => \N__20122\,
            I => \N__20116\
        );

    \I__3369\ : CascadeBuf
    port map (
            O => \N__20119\,
            I => \N__20113\
        );

    \I__3368\ : CascadeMux
    port map (
            O => \N__20116\,
            I => \N__20110\
        );

    \I__3367\ : CascadeMux
    port map (
            O => \N__20113\,
            I => \N__20107\
        );

    \I__3366\ : CascadeBuf
    port map (
            O => \N__20110\,
            I => \N__20104\
        );

    \I__3365\ : CascadeBuf
    port map (
            O => \N__20107\,
            I => \N__20101\
        );

    \I__3364\ : CascadeMux
    port map (
            O => \N__20104\,
            I => \N__20098\
        );

    \I__3363\ : CascadeMux
    port map (
            O => \N__20101\,
            I => \N__20095\
        );

    \I__3362\ : CascadeBuf
    port map (
            O => \N__20098\,
            I => \N__20092\
        );

    \I__3361\ : CascadeBuf
    port map (
            O => \N__20095\,
            I => \N__20089\
        );

    \I__3360\ : CascadeMux
    port map (
            O => \N__20092\,
            I => \N__20086\
        );

    \I__3359\ : CascadeMux
    port map (
            O => \N__20089\,
            I => \N__20083\
        );

    \I__3358\ : CascadeBuf
    port map (
            O => \N__20086\,
            I => \N__20080\
        );

    \I__3357\ : CascadeBuf
    port map (
            O => \N__20083\,
            I => \N__20077\
        );

    \I__3356\ : CascadeMux
    port map (
            O => \N__20080\,
            I => \N__20074\
        );

    \I__3355\ : CascadeMux
    port map (
            O => \N__20077\,
            I => \N__20071\
        );

    \I__3354\ : InMux
    port map (
            O => \N__20074\,
            I => \N__20068\
        );

    \I__3353\ : InMux
    port map (
            O => \N__20071\,
            I => \N__20065\
        );

    \I__3352\ : LocalMux
    port map (
            O => \N__20068\,
            I => \N__20062\
        );

    \I__3351\ : LocalMux
    port map (
            O => \N__20065\,
            I => \N__20059\
        );

    \I__3350\ : Span4Mux_v
    port map (
            O => \N__20062\,
            I => \N__20056\
        );

    \I__3349\ : Span4Mux_v
    port map (
            O => \N__20059\,
            I => \N__20053\
        );

    \I__3348\ : Span4Mux_h
    port map (
            O => \N__20056\,
            I => \N__20048\
        );

    \I__3347\ : Span4Mux_h
    port map (
            O => \N__20053\,
            I => \N__20048\
        );

    \I__3346\ : Span4Mux_h
    port map (
            O => \N__20048\,
            I => \N__20045\
        );

    \I__3345\ : Odrv4
    port map (
            O => \N__20045\,
            I => \SYNTHESIZED_WIRE_12_10\
        );

    \I__3344\ : InMux
    port map (
            O => \N__20042\,
            I => \N__20039\
        );

    \I__3343\ : LocalMux
    port map (
            O => \N__20039\,
            I => \N__20036\
        );

    \I__3342\ : Span4Mux_h
    port map (
            O => \N__20036\,
            I => \N__20033\
        );

    \I__3341\ : Sp12to4
    port map (
            O => \N__20033\,
            I => \N__20030\
        );

    \I__3340\ : Span12Mux_v
    port map (
            O => \N__20030\,
            I => \N__20027\
        );

    \I__3339\ : Span12Mux_h
    port map (
            O => \N__20027\,
            I => \N__20024\
        );

    \I__3338\ : Odrv12
    port map (
            O => \N__20024\,
            I => swit_c_2
        );

    \I__3337\ : CascadeMux
    port map (
            O => \N__20021\,
            I => \b2v_inst.addr_ram_energia_m0_2_cascade_\
        );

    \I__3336\ : CascadeMux
    port map (
            O => \N__20018\,
            I => \N__20014\
        );

    \I__3335\ : CascadeMux
    port map (
            O => \N__20017\,
            I => \N__20011\
        );

    \I__3334\ : CascadeBuf
    port map (
            O => \N__20014\,
            I => \N__20008\
        );

    \I__3333\ : CascadeBuf
    port map (
            O => \N__20011\,
            I => \N__20005\
        );

    \I__3332\ : CascadeMux
    port map (
            O => \N__20008\,
            I => \N__20002\
        );

    \I__3331\ : CascadeMux
    port map (
            O => \N__20005\,
            I => \N__19999\
        );

    \I__3330\ : CascadeBuf
    port map (
            O => \N__20002\,
            I => \N__19996\
        );

    \I__3329\ : CascadeBuf
    port map (
            O => \N__19999\,
            I => \N__19993\
        );

    \I__3328\ : CascadeMux
    port map (
            O => \N__19996\,
            I => \N__19990\
        );

    \I__3327\ : CascadeMux
    port map (
            O => \N__19993\,
            I => \N__19987\
        );

    \I__3326\ : CascadeBuf
    port map (
            O => \N__19990\,
            I => \N__19984\
        );

    \I__3325\ : CascadeBuf
    port map (
            O => \N__19987\,
            I => \N__19981\
        );

    \I__3324\ : CascadeMux
    port map (
            O => \N__19984\,
            I => \N__19978\
        );

    \I__3323\ : CascadeMux
    port map (
            O => \N__19981\,
            I => \N__19975\
        );

    \I__3322\ : CascadeBuf
    port map (
            O => \N__19978\,
            I => \N__19972\
        );

    \I__3321\ : CascadeBuf
    port map (
            O => \N__19975\,
            I => \N__19969\
        );

    \I__3320\ : CascadeMux
    port map (
            O => \N__19972\,
            I => \N__19966\
        );

    \I__3319\ : CascadeMux
    port map (
            O => \N__19969\,
            I => \N__19963\
        );

    \I__3318\ : CascadeBuf
    port map (
            O => \N__19966\,
            I => \N__19960\
        );

    \I__3317\ : CascadeBuf
    port map (
            O => \N__19963\,
            I => \N__19957\
        );

    \I__3316\ : CascadeMux
    port map (
            O => \N__19960\,
            I => \N__19954\
        );

    \I__3315\ : CascadeMux
    port map (
            O => \N__19957\,
            I => \N__19951\
        );

    \I__3314\ : CascadeBuf
    port map (
            O => \N__19954\,
            I => \N__19948\
        );

    \I__3313\ : CascadeBuf
    port map (
            O => \N__19951\,
            I => \N__19945\
        );

    \I__3312\ : CascadeMux
    port map (
            O => \N__19948\,
            I => \N__19942\
        );

    \I__3311\ : CascadeMux
    port map (
            O => \N__19945\,
            I => \N__19939\
        );

    \I__3310\ : InMux
    port map (
            O => \N__19942\,
            I => \N__19936\
        );

    \I__3309\ : InMux
    port map (
            O => \N__19939\,
            I => \N__19933\
        );

    \I__3308\ : LocalMux
    port map (
            O => \N__19936\,
            I => \N__19928\
        );

    \I__3307\ : LocalMux
    port map (
            O => \N__19933\,
            I => \N__19928\
        );

    \I__3306\ : Span4Mux_v
    port map (
            O => \N__19928\,
            I => \N__19925\
        );

    \I__3305\ : Span4Mux_h
    port map (
            O => \N__19925\,
            I => \N__19922\
        );

    \I__3304\ : Span4Mux_h
    port map (
            O => \N__19922\,
            I => \N__19919\
        );

    \I__3303\ : Odrv4
    port map (
            O => \N__19919\,
            I => \SYNTHESIZED_WIRE_12_2\
        );

    \I__3302\ : InMux
    port map (
            O => \N__19916\,
            I => \N__19913\
        );

    \I__3301\ : LocalMux
    port map (
            O => \N__19913\,
            I => \N__19910\
        );

    \I__3300\ : Span12Mux_h
    port map (
            O => \N__19910\,
            I => \N__19907\
        );

    \I__3299\ : Odrv12
    port map (
            O => \N__19907\,
            I => swit_c_5
        );

    \I__3298\ : CascadeMux
    port map (
            O => \N__19904\,
            I => \b2v_inst.addr_ram_energia_m0_5_cascade_\
        );

    \I__3297\ : CascadeMux
    port map (
            O => \N__19901\,
            I => \N__19897\
        );

    \I__3296\ : CascadeMux
    port map (
            O => \N__19900\,
            I => \N__19894\
        );

    \I__3295\ : CascadeBuf
    port map (
            O => \N__19897\,
            I => \N__19891\
        );

    \I__3294\ : CascadeBuf
    port map (
            O => \N__19894\,
            I => \N__19888\
        );

    \I__3293\ : CascadeMux
    port map (
            O => \N__19891\,
            I => \N__19885\
        );

    \I__3292\ : CascadeMux
    port map (
            O => \N__19888\,
            I => \N__19882\
        );

    \I__3291\ : CascadeBuf
    port map (
            O => \N__19885\,
            I => \N__19879\
        );

    \I__3290\ : CascadeBuf
    port map (
            O => \N__19882\,
            I => \N__19876\
        );

    \I__3289\ : CascadeMux
    port map (
            O => \N__19879\,
            I => \N__19873\
        );

    \I__3288\ : CascadeMux
    port map (
            O => \N__19876\,
            I => \N__19870\
        );

    \I__3287\ : CascadeBuf
    port map (
            O => \N__19873\,
            I => \N__19867\
        );

    \I__3286\ : CascadeBuf
    port map (
            O => \N__19870\,
            I => \N__19864\
        );

    \I__3285\ : CascadeMux
    port map (
            O => \N__19867\,
            I => \N__19861\
        );

    \I__3284\ : CascadeMux
    port map (
            O => \N__19864\,
            I => \N__19858\
        );

    \I__3283\ : CascadeBuf
    port map (
            O => \N__19861\,
            I => \N__19855\
        );

    \I__3282\ : CascadeBuf
    port map (
            O => \N__19858\,
            I => \N__19852\
        );

    \I__3281\ : CascadeMux
    port map (
            O => \N__19855\,
            I => \N__19849\
        );

    \I__3280\ : CascadeMux
    port map (
            O => \N__19852\,
            I => \N__19846\
        );

    \I__3279\ : CascadeBuf
    port map (
            O => \N__19849\,
            I => \N__19843\
        );

    \I__3278\ : CascadeBuf
    port map (
            O => \N__19846\,
            I => \N__19840\
        );

    \I__3277\ : CascadeMux
    port map (
            O => \N__19843\,
            I => \N__19837\
        );

    \I__3276\ : CascadeMux
    port map (
            O => \N__19840\,
            I => \N__19834\
        );

    \I__3275\ : CascadeBuf
    port map (
            O => \N__19837\,
            I => \N__19831\
        );

    \I__3274\ : CascadeBuf
    port map (
            O => \N__19834\,
            I => \N__19828\
        );

    \I__3273\ : CascadeMux
    port map (
            O => \N__19831\,
            I => \N__19825\
        );

    \I__3272\ : CascadeMux
    port map (
            O => \N__19828\,
            I => \N__19822\
        );

    \I__3271\ : InMux
    port map (
            O => \N__19825\,
            I => \N__19819\
        );

    \I__3270\ : InMux
    port map (
            O => \N__19822\,
            I => \N__19816\
        );

    \I__3269\ : LocalMux
    port map (
            O => \N__19819\,
            I => \N__19811\
        );

    \I__3268\ : LocalMux
    port map (
            O => \N__19816\,
            I => \N__19811\
        );

    \I__3267\ : Span4Mux_v
    port map (
            O => \N__19811\,
            I => \N__19808\
        );

    \I__3266\ : Span4Mux_h
    port map (
            O => \N__19808\,
            I => \N__19805\
        );

    \I__3265\ : Span4Mux_h
    port map (
            O => \N__19805\,
            I => \N__19802\
        );

    \I__3264\ : Odrv4
    port map (
            O => \N__19802\,
            I => \SYNTHESIZED_WIRE_12_5\
        );

    \I__3263\ : InMux
    port map (
            O => \N__19799\,
            I => \N__19796\
        );

    \I__3262\ : LocalMux
    port map (
            O => \N__19796\,
            I => \N__19793\
        );

    \I__3261\ : Span4Mux_v
    port map (
            O => \N__19793\,
            I => \N__19790\
        );

    \I__3260\ : Sp12to4
    port map (
            O => \N__19790\,
            I => \N__19787\
        );

    \I__3259\ : Span12Mux_v
    port map (
            O => \N__19787\,
            I => \N__19784\
        );

    \I__3258\ : Span12Mux_h
    port map (
            O => \N__19784\,
            I => \N__19781\
        );

    \I__3257\ : Odrv12
    port map (
            O => \N__19781\,
            I => swit_c_10
        );

    \I__3256\ : InMux
    port map (
            O => \N__19778\,
            I => \N__19775\
        );

    \I__3255\ : LocalMux
    port map (
            O => \N__19775\,
            I => \b2v_inst.addr_ram_energia_m0_10\
        );

    \I__3254\ : InMux
    port map (
            O => \N__19772\,
            I => \N__19769\
        );

    \I__3253\ : LocalMux
    port map (
            O => \N__19769\,
            I => \N__19766\
        );

    \I__3252\ : Span4Mux_h
    port map (
            O => \N__19766\,
            I => \N__19763\
        );

    \I__3251\ : Sp12to4
    port map (
            O => \N__19763\,
            I => \N__19760\
        );

    \I__3250\ : Odrv12
    port map (
            O => \N__19760\,
            I => swit_c_3
        );

    \I__3249\ : CascadeMux
    port map (
            O => \N__19757\,
            I => \b2v_inst.N_514_cascade_\
        );

    \I__3248\ : InMux
    port map (
            O => \N__19754\,
            I => \N__19751\
        );

    \I__3247\ : LocalMux
    port map (
            O => \N__19751\,
            I => \N__19748\
        );

    \I__3246\ : Span4Mux_h
    port map (
            O => \N__19748\,
            I => \N__19745\
        );

    \I__3245\ : Span4Mux_v
    port map (
            O => \N__19745\,
            I => \N__19742\
        );

    \I__3244\ : Span4Mux_h
    port map (
            O => \N__19742\,
            I => \N__19739\
        );

    \I__3243\ : Span4Mux_h
    port map (
            O => \N__19739\,
            I => \N__19736\
        );

    \I__3242\ : Odrv4
    port map (
            O => \N__19736\,
            I => \N_116_i\
        );

    \I__3241\ : InMux
    port map (
            O => \N__19733\,
            I => \N__19730\
        );

    \I__3240\ : LocalMux
    port map (
            O => \N__19730\,
            I => \N__19725\
        );

    \I__3239\ : InMux
    port map (
            O => \N__19729\,
            I => \N__19720\
        );

    \I__3238\ : InMux
    port map (
            O => \N__19728\,
            I => \N__19720\
        );

    \I__3237\ : Odrv4
    port map (
            O => \N__19725\,
            I => \b2v_inst.stateZ0Z_16\
        );

    \I__3236\ : LocalMux
    port map (
            O => \N__19720\,
            I => \b2v_inst.stateZ0Z_16\
        );

    \I__3235\ : InMux
    port map (
            O => \N__19715\,
            I => \N__19712\
        );

    \I__3234\ : LocalMux
    port map (
            O => \N__19712\,
            I => \N__19709\
        );

    \I__3233\ : Span4Mux_h
    port map (
            O => \N__19709\,
            I => \N__19706\
        );

    \I__3232\ : Span4Mux_h
    port map (
            O => \N__19706\,
            I => \N__19703\
        );

    \I__3231\ : Odrv4
    port map (
            O => \N__19703\,
            I => \N_548_i\
        );

    \I__3230\ : CascadeMux
    port map (
            O => \N__19700\,
            I => \N__19697\
        );

    \I__3229\ : InMux
    port map (
            O => \N__19697\,
            I => \N__19694\
        );

    \I__3228\ : LocalMux
    port map (
            O => \N__19694\,
            I => \N__19688\
        );

    \I__3227\ : CascadeMux
    port map (
            O => \N__19693\,
            I => \N__19685\
        );

    \I__3226\ : CascadeMux
    port map (
            O => \N__19692\,
            I => \N__19682\
        );

    \I__3225\ : InMux
    port map (
            O => \N__19691\,
            I => \N__19679\
        );

    \I__3224\ : Span4Mux_v
    port map (
            O => \N__19688\,
            I => \N__19676\
        );

    \I__3223\ : InMux
    port map (
            O => \N__19685\,
            I => \N__19671\
        );

    \I__3222\ : InMux
    port map (
            O => \N__19682\,
            I => \N__19671\
        );

    \I__3221\ : LocalMux
    port map (
            O => \N__19679\,
            I => \b2v_inst.stateZ0Z_0\
        );

    \I__3220\ : Odrv4
    port map (
            O => \N__19676\,
            I => \b2v_inst.stateZ0Z_0\
        );

    \I__3219\ : LocalMux
    port map (
            O => \N__19671\,
            I => \b2v_inst.stateZ0Z_0\
        );

    \I__3218\ : CascadeMux
    port map (
            O => \N__19664\,
            I => \b2v_inst.N_692_cascade_\
        );

    \I__3217\ : CascadeMux
    port map (
            O => \N__19661\,
            I => \b2v_inst.addr_ram_iv_i_0_0_3_cascade_\
        );

    \I__3216\ : CascadeMux
    port map (
            O => \N__19658\,
            I => \N__19655\
        );

    \I__3215\ : CascadeBuf
    port map (
            O => \N__19655\,
            I => \N__19652\
        );

    \I__3214\ : CascadeMux
    port map (
            O => \N__19652\,
            I => \N__19648\
        );

    \I__3213\ : CascadeMux
    port map (
            O => \N__19651\,
            I => \N__19645\
        );

    \I__3212\ : CascadeBuf
    port map (
            O => \N__19648\,
            I => \N__19642\
        );

    \I__3211\ : CascadeBuf
    port map (
            O => \N__19645\,
            I => \N__19639\
        );

    \I__3210\ : CascadeMux
    port map (
            O => \N__19642\,
            I => \N__19636\
        );

    \I__3209\ : CascadeMux
    port map (
            O => \N__19639\,
            I => \N__19633\
        );

    \I__3208\ : CascadeBuf
    port map (
            O => \N__19636\,
            I => \N__19630\
        );

    \I__3207\ : CascadeBuf
    port map (
            O => \N__19633\,
            I => \N__19627\
        );

    \I__3206\ : CascadeMux
    port map (
            O => \N__19630\,
            I => \N__19624\
        );

    \I__3205\ : CascadeMux
    port map (
            O => \N__19627\,
            I => \N__19621\
        );

    \I__3204\ : CascadeBuf
    port map (
            O => \N__19624\,
            I => \N__19618\
        );

    \I__3203\ : CascadeBuf
    port map (
            O => \N__19621\,
            I => \N__19615\
        );

    \I__3202\ : CascadeMux
    port map (
            O => \N__19618\,
            I => \N__19612\
        );

    \I__3201\ : CascadeMux
    port map (
            O => \N__19615\,
            I => \N__19609\
        );

    \I__3200\ : CascadeBuf
    port map (
            O => \N__19612\,
            I => \N__19606\
        );

    \I__3199\ : CascadeBuf
    port map (
            O => \N__19609\,
            I => \N__19603\
        );

    \I__3198\ : CascadeMux
    port map (
            O => \N__19606\,
            I => \N__19600\
        );

    \I__3197\ : CascadeMux
    port map (
            O => \N__19603\,
            I => \N__19597\
        );

    \I__3196\ : InMux
    port map (
            O => \N__19600\,
            I => \N__19594\
        );

    \I__3195\ : CascadeBuf
    port map (
            O => \N__19597\,
            I => \N__19591\
        );

    \I__3194\ : LocalMux
    port map (
            O => \N__19594\,
            I => \N__19588\
        );

    \I__3193\ : CascadeMux
    port map (
            O => \N__19591\,
            I => \N__19585\
        );

    \I__3192\ : Span4Mux_v
    port map (
            O => \N__19588\,
            I => \N__19582\
        );

    \I__3191\ : InMux
    port map (
            O => \N__19585\,
            I => \N__19579\
        );

    \I__3190\ : Span4Mux_h
    port map (
            O => \N__19582\,
            I => \N__19576\
        );

    \I__3189\ : LocalMux
    port map (
            O => \N__19579\,
            I => \N__19573\
        );

    \I__3188\ : Span4Mux_h
    port map (
            O => \N__19576\,
            I => \N__19570\
        );

    \I__3187\ : Odrv12
    port map (
            O => \N__19573\,
            I => \indice_RNIIU233_3\
        );

    \I__3186\ : Odrv4
    port map (
            O => \N__19570\,
            I => \indice_RNIIU233_3\
        );

    \I__3185\ : InMux
    port map (
            O => \N__19565\,
            I => \N__19562\
        );

    \I__3184\ : LocalMux
    port map (
            O => \N__19562\,
            I => \N__19559\
        );

    \I__3183\ : Span4Mux_h
    port map (
            O => \N__19559\,
            I => \N__19556\
        );

    \I__3182\ : Span4Mux_v
    port map (
            O => \N__19556\,
            I => \N__19553\
        );

    \I__3181\ : Odrv4
    port map (
            O => \N__19553\,
            I => \b2v_inst.dir_mem_3Z0Z_3\
        );

    \I__3180\ : InMux
    port map (
            O => \N__19550\,
            I => \N__19547\
        );

    \I__3179\ : LocalMux
    port map (
            O => \N__19547\,
            I => \N__19544\
        );

    \I__3178\ : Span4Mux_v
    port map (
            O => \N__19544\,
            I => \N__19541\
        );

    \I__3177\ : Odrv4
    port map (
            O => \N__19541\,
            I => \b2v_inst.dir_mem_1Z0Z_3\
        );

    \I__3176\ : InMux
    port map (
            O => \N__19538\,
            I => \N__19535\
        );

    \I__3175\ : LocalMux
    port map (
            O => \N__19535\,
            I => \b2v_inst.addr_ram_iv_i_0_1_3\
        );

    \I__3174\ : InMux
    port map (
            O => \N__19532\,
            I => \N__19529\
        );

    \I__3173\ : LocalMux
    port map (
            O => \N__19529\,
            I => \b2v_inst.dir_memZ0Z_0\
        );

    \I__3172\ : InMux
    port map (
            O => \N__19526\,
            I => \N__19522\
        );

    \I__3171\ : InMux
    port map (
            O => \N__19525\,
            I => \N__19519\
        );

    \I__3170\ : LocalMux
    port map (
            O => \N__19522\,
            I => \N__19516\
        );

    \I__3169\ : LocalMux
    port map (
            O => \N__19519\,
            I => \N__19511\
        );

    \I__3168\ : Span4Mux_v
    port map (
            O => \N__19516\,
            I => \N__19511\
        );

    \I__3167\ : Odrv4
    port map (
            O => \N__19511\,
            I => \b2v_inst.N_618_6\
        );

    \I__3166\ : InMux
    port map (
            O => \N__19508\,
            I => \N__19505\
        );

    \I__3165\ : LocalMux
    port map (
            O => \N__19505\,
            I => \N__19502\
        );

    \I__3164\ : Odrv4
    port map (
            O => \N__19502\,
            I => \b2v_inst.dir_mem_1Z0Z_7\
        );

    \I__3163\ : InMux
    port map (
            O => \N__19499\,
            I => \N__19496\
        );

    \I__3162\ : LocalMux
    port map (
            O => \N__19496\,
            I => \N__19493\
        );

    \I__3161\ : Span4Mux_v
    port map (
            O => \N__19493\,
            I => \N__19490\
        );

    \I__3160\ : Span4Mux_h
    port map (
            O => \N__19490\,
            I => \N__19487\
        );

    \I__3159\ : Odrv4
    port map (
            O => \N__19487\,
            I => \b2v_inst.dir_mem_3Z0Z_7\
        );

    \I__3158\ : CascadeMux
    port map (
            O => \N__19484\,
            I => \b2v_inst.N_488_cascade_\
        );

    \I__3157\ : InMux
    port map (
            O => \N__19481\,
            I => \N__19478\
        );

    \I__3156\ : LocalMux
    port map (
            O => \N__19478\,
            I => \b2v_inst.addr_ram_iv_i_0_0_7\
        );

    \I__3155\ : CascadeMux
    port map (
            O => \N__19475\,
            I => \b2v_inst.addr_ram_iv_i_0_1_7_cascade_\
        );

    \I__3154\ : CascadeMux
    port map (
            O => \N__19472\,
            I => \N__19468\
        );

    \I__3153\ : CascadeMux
    port map (
            O => \N__19471\,
            I => \N__19465\
        );

    \I__3152\ : CascadeBuf
    port map (
            O => \N__19468\,
            I => \N__19462\
        );

    \I__3151\ : CascadeBuf
    port map (
            O => \N__19465\,
            I => \N__19459\
        );

    \I__3150\ : CascadeMux
    port map (
            O => \N__19462\,
            I => \N__19456\
        );

    \I__3149\ : CascadeMux
    port map (
            O => \N__19459\,
            I => \N__19453\
        );

    \I__3148\ : CascadeBuf
    port map (
            O => \N__19456\,
            I => \N__19450\
        );

    \I__3147\ : CascadeBuf
    port map (
            O => \N__19453\,
            I => \N__19447\
        );

    \I__3146\ : CascadeMux
    port map (
            O => \N__19450\,
            I => \N__19444\
        );

    \I__3145\ : CascadeMux
    port map (
            O => \N__19447\,
            I => \N__19441\
        );

    \I__3144\ : CascadeBuf
    port map (
            O => \N__19444\,
            I => \N__19438\
        );

    \I__3143\ : CascadeBuf
    port map (
            O => \N__19441\,
            I => \N__19435\
        );

    \I__3142\ : CascadeMux
    port map (
            O => \N__19438\,
            I => \N__19432\
        );

    \I__3141\ : CascadeMux
    port map (
            O => \N__19435\,
            I => \N__19429\
        );

    \I__3140\ : CascadeBuf
    port map (
            O => \N__19432\,
            I => \N__19426\
        );

    \I__3139\ : CascadeBuf
    port map (
            O => \N__19429\,
            I => \N__19423\
        );

    \I__3138\ : CascadeMux
    port map (
            O => \N__19426\,
            I => \N__19420\
        );

    \I__3137\ : CascadeMux
    port map (
            O => \N__19423\,
            I => \N__19417\
        );

    \I__3136\ : CascadeBuf
    port map (
            O => \N__19420\,
            I => \N__19414\
        );

    \I__3135\ : CascadeBuf
    port map (
            O => \N__19417\,
            I => \N__19411\
        );

    \I__3134\ : CascadeMux
    port map (
            O => \N__19414\,
            I => \N__19408\
        );

    \I__3133\ : CascadeMux
    port map (
            O => \N__19411\,
            I => \N__19405\
        );

    \I__3132\ : InMux
    port map (
            O => \N__19408\,
            I => \N__19402\
        );

    \I__3131\ : InMux
    port map (
            O => \N__19405\,
            I => \N__19399\
        );

    \I__3130\ : LocalMux
    port map (
            O => \N__19402\,
            I => \N__19394\
        );

    \I__3129\ : LocalMux
    port map (
            O => \N__19399\,
            I => \N__19394\
        );

    \I__3128\ : Span12Mux_v
    port map (
            O => \N__19394\,
            I => \N__19391\
        );

    \I__3127\ : Odrv12
    port map (
            O => \N__19391\,
            I => \indice_RNI6J333_7\
        );

    \I__3126\ : InMux
    port map (
            O => \N__19388\,
            I => \N__19385\
        );

    \I__3125\ : LocalMux
    port map (
            O => \N__19385\,
            I => \N__19382\
        );

    \I__3124\ : Span4Mux_v
    port map (
            O => \N__19382\,
            I => \N__19379\
        );

    \I__3123\ : Odrv4
    port map (
            O => \N__19379\,
            I => \b2v_inst.state_RNO_0Z0Z_29\
        );

    \I__3122\ : InMux
    port map (
            O => \N__19376\,
            I => \N__19373\
        );

    \I__3121\ : LocalMux
    port map (
            O => \N__19373\,
            I => \N__19370\
        );

    \I__3120\ : Span4Mux_v
    port map (
            O => \N__19370\,
            I => \N__19367\
        );

    \I__3119\ : Odrv4
    port map (
            O => \N__19367\,
            I => \b2v_inst.dir_mem_1Z0Z_0\
        );

    \I__3118\ : CascadeMux
    port map (
            O => \N__19364\,
            I => \N__19361\
        );

    \I__3117\ : InMux
    port map (
            O => \N__19361\,
            I => \N__19358\
        );

    \I__3116\ : LocalMux
    port map (
            O => \N__19358\,
            I => \N__19355\
        );

    \I__3115\ : Span4Mux_v
    port map (
            O => \N__19355\,
            I => \N__19352\
        );

    \I__3114\ : Span4Mux_h
    port map (
            O => \N__19352\,
            I => \N__19349\
        );

    \I__3113\ : Odrv4
    port map (
            O => \N__19349\,
            I => \b2v_inst.dir_mem_3Z0Z_0\
        );

    \I__3112\ : InMux
    port map (
            O => \N__19346\,
            I => \N__19343\
        );

    \I__3111\ : LocalMux
    port map (
            O => \N__19343\,
            I => \N__19340\
        );

    \I__3110\ : Span4Mux_v
    port map (
            O => \N__19340\,
            I => \N__19337\
        );

    \I__3109\ : Odrv4
    port map (
            O => \N__19337\,
            I => \b2v_inst.dir_mem_2Z0Z_3\
        );

    \I__3108\ : InMux
    port map (
            O => \N__19334\,
            I => \N__19331\
        );

    \I__3107\ : LocalMux
    port map (
            O => \N__19331\,
            I => \N__19328\
        );

    \I__3106\ : Span4Mux_v
    port map (
            O => \N__19328\,
            I => \N__19325\
        );

    \I__3105\ : Odrv4
    port map (
            O => \N__19325\,
            I => \b2v_inst.dir_memZ0Z_3\
        );

    \I__3104\ : InMux
    port map (
            O => \N__19322\,
            I => \N__19319\
        );

    \I__3103\ : LocalMux
    port map (
            O => \N__19319\,
            I => \N__19316\
        );

    \I__3102\ : Span4Mux_h
    port map (
            O => \N__19316\,
            I => \N__19313\
        );

    \I__3101\ : Odrv4
    port map (
            O => \N__19313\,
            I => \b2v_inst.dir_mem_3Z0Z_1\
        );

    \I__3100\ : InMux
    port map (
            O => \N__19310\,
            I => \N__19307\
        );

    \I__3099\ : LocalMux
    port map (
            O => \N__19307\,
            I => \N__19304\
        );

    \I__3098\ : Odrv4
    port map (
            O => \N__19304\,
            I => \b2v_inst.dir_memZ0Z_1\
        );

    \I__3097\ : CascadeMux
    port map (
            O => \N__19301\,
            I => \N__19298\
        );

    \I__3096\ : InMux
    port map (
            O => \N__19298\,
            I => \N__19295\
        );

    \I__3095\ : LocalMux
    port map (
            O => \N__19295\,
            I => \N__19292\
        );

    \I__3094\ : Span4Mux_v
    port map (
            O => \N__19292\,
            I => \N__19289\
        );

    \I__3093\ : Odrv4
    port map (
            O => \N__19289\,
            I => \b2v_inst.dir_mem_2Z0Z_1\
        );

    \I__3092\ : InMux
    port map (
            O => \N__19286\,
            I => \N__19283\
        );

    \I__3091\ : LocalMux
    port map (
            O => \N__19283\,
            I => \N__19279\
        );

    \I__3090\ : InMux
    port map (
            O => \N__19282\,
            I => \N__19276\
        );

    \I__3089\ : Span4Mux_h
    port map (
            O => \N__19279\,
            I => \N__19270\
        );

    \I__3088\ : LocalMux
    port map (
            O => \N__19276\,
            I => \N__19270\
        );

    \I__3087\ : CascadeMux
    port map (
            O => \N__19275\,
            I => \N__19267\
        );

    \I__3086\ : Span4Mux_h
    port map (
            O => \N__19270\,
            I => \N__19264\
        );

    \I__3085\ : InMux
    port map (
            O => \N__19267\,
            I => \N__19261\
        );

    \I__3084\ : Odrv4
    port map (
            O => \N__19264\,
            I => \b2v_inst.un8_dir_mem_1_cry_0_c_RNI4SNCZ0\
        );

    \I__3083\ : LocalMux
    port map (
            O => \N__19261\,
            I => \b2v_inst.un8_dir_mem_1_cry_0_c_RNI4SNCZ0\
        );

    \I__3082\ : InMux
    port map (
            O => \N__19256\,
            I => \N__19253\
        );

    \I__3081\ : LocalMux
    port map (
            O => \N__19253\,
            I => \b2v_inst.dir_mem_1Z0Z_1\
        );

    \I__3080\ : InMux
    port map (
            O => \N__19250\,
            I => \N__19236\
        );

    \I__3079\ : InMux
    port map (
            O => \N__19249\,
            I => \N__19236\
        );

    \I__3078\ : InMux
    port map (
            O => \N__19248\,
            I => \N__19229\
        );

    \I__3077\ : InMux
    port map (
            O => \N__19247\,
            I => \N__19229\
        );

    \I__3076\ : InMux
    port map (
            O => \N__19246\,
            I => \N__19229\
        );

    \I__3075\ : InMux
    port map (
            O => \N__19245\,
            I => \N__19218\
        );

    \I__3074\ : InMux
    port map (
            O => \N__19244\,
            I => \N__19218\
        );

    \I__3073\ : InMux
    port map (
            O => \N__19243\,
            I => \N__19218\
        );

    \I__3072\ : InMux
    port map (
            O => \N__19242\,
            I => \N__19218\
        );

    \I__3071\ : InMux
    port map (
            O => \N__19241\,
            I => \N__19218\
        );

    \I__3070\ : LocalMux
    port map (
            O => \N__19236\,
            I => \b2v_inst.dir_mem_115lt11\
        );

    \I__3069\ : LocalMux
    port map (
            O => \N__19229\,
            I => \b2v_inst.dir_mem_115lt11\
        );

    \I__3068\ : LocalMux
    port map (
            O => \N__19218\,
            I => \b2v_inst.dir_mem_115lt11\
        );

    \I__3067\ : InMux
    port map (
            O => \N__19211\,
            I => \N__19207\
        );

    \I__3066\ : InMux
    port map (
            O => \N__19210\,
            I => \N__19204\
        );

    \I__3065\ : LocalMux
    port map (
            O => \N__19207\,
            I => \N__19201\
        );

    \I__3064\ : LocalMux
    port map (
            O => \N__19204\,
            I => \N__19195\
        );

    \I__3063\ : Span4Mux_v
    port map (
            O => \N__19201\,
            I => \N__19195\
        );

    \I__3062\ : CascadeMux
    port map (
            O => \N__19200\,
            I => \N__19192\
        );

    \I__3061\ : Span4Mux_h
    port map (
            O => \N__19195\,
            I => \N__19189\
        );

    \I__3060\ : InMux
    port map (
            O => \N__19192\,
            I => \N__19186\
        );

    \I__3059\ : Odrv4
    port map (
            O => \N__19189\,
            I => \b2v_inst.indice_RNILHHBZ0Z_2\
        );

    \I__3058\ : LocalMux
    port map (
            O => \N__19186\,
            I => \b2v_inst.indice_RNILHHBZ0Z_2\
        );

    \I__3057\ : CascadeMux
    port map (
            O => \N__19181\,
            I => \N__19175\
        );

    \I__3056\ : CascadeMux
    port map (
            O => \N__19180\,
            I => \N__19172\
        );

    \I__3055\ : CascadeMux
    port map (
            O => \N__19179\,
            I => \N__19169\
        );

    \I__3054\ : InMux
    port map (
            O => \N__19178\,
            I => \N__19159\
        );

    \I__3053\ : InMux
    port map (
            O => \N__19175\,
            I => \N__19159\
        );

    \I__3052\ : InMux
    port map (
            O => \N__19172\,
            I => \N__19156\
        );

    \I__3051\ : InMux
    port map (
            O => \N__19169\,
            I => \N__19151\
        );

    \I__3050\ : InMux
    port map (
            O => \N__19168\,
            I => \N__19151\
        );

    \I__3049\ : InMux
    port map (
            O => \N__19167\,
            I => \N__19142\
        );

    \I__3048\ : InMux
    port map (
            O => \N__19166\,
            I => \N__19142\
        );

    \I__3047\ : InMux
    port map (
            O => \N__19165\,
            I => \N__19142\
        );

    \I__3046\ : InMux
    port map (
            O => \N__19164\,
            I => \N__19142\
        );

    \I__3045\ : LocalMux
    port map (
            O => \N__19159\,
            I => \N__19139\
        );

    \I__3044\ : LocalMux
    port map (
            O => \N__19156\,
            I => \b2v_inst.dir_mem_115lto11_0\
        );

    \I__3043\ : LocalMux
    port map (
            O => \N__19151\,
            I => \b2v_inst.dir_mem_115lto11_0\
        );

    \I__3042\ : LocalMux
    port map (
            O => \N__19142\,
            I => \b2v_inst.dir_mem_115lto11_0\
        );

    \I__3041\ : Odrv12
    port map (
            O => \N__19139\,
            I => \b2v_inst.dir_mem_115lto11_0\
        );

    \I__3040\ : InMux
    port map (
            O => \N__19130\,
            I => \N__19127\
        );

    \I__3039\ : LocalMux
    port map (
            O => \N__19127\,
            I => \N__19124\
        );

    \I__3038\ : Span12Mux_h
    port map (
            O => \N__19124\,
            I => \N__19120\
        );

    \I__3037\ : InMux
    port map (
            O => \N__19123\,
            I => \N__19117\
        );

    \I__3036\ : Odrv12
    port map (
            O => \N__19120\,
            I => \b2v_inst.un8_dir_mem_1_cry_1_c_RNI6VOCZ0\
        );

    \I__3035\ : LocalMux
    port map (
            O => \N__19117\,
            I => \b2v_inst.un8_dir_mem_1_cry_1_c_RNI6VOCZ0\
        );

    \I__3034\ : CEMux
    port map (
            O => \N__19112\,
            I => \N__19108\
        );

    \I__3033\ : CEMux
    port map (
            O => \N__19111\,
            I => \N__19105\
        );

    \I__3032\ : LocalMux
    port map (
            O => \N__19108\,
            I => \N__19101\
        );

    \I__3031\ : LocalMux
    port map (
            O => \N__19105\,
            I => \N__19098\
        );

    \I__3030\ : CEMux
    port map (
            O => \N__19104\,
            I => \N__19095\
        );

    \I__3029\ : Span4Mux_v
    port map (
            O => \N__19101\,
            I => \N__19092\
        );

    \I__3028\ : Span4Mux_h
    port map (
            O => \N__19098\,
            I => \N__19089\
        );

    \I__3027\ : LocalMux
    port map (
            O => \N__19095\,
            I => \N__19086\
        );

    \I__3026\ : Odrv4
    port map (
            O => \N__19092\,
            I => \b2v_inst.N_363_i\
        );

    \I__3025\ : Odrv4
    port map (
            O => \N__19089\,
            I => \b2v_inst.N_363_i\
        );

    \I__3024\ : Odrv4
    port map (
            O => \N__19086\,
            I => \b2v_inst.N_363_i\
        );

    \I__3023\ : InMux
    port map (
            O => \N__19079\,
            I => \N__19076\
        );

    \I__3022\ : LocalMux
    port map (
            O => \N__19076\,
            I => \N__19073\
        );

    \I__3021\ : Odrv4
    port map (
            O => \N__19073\,
            I => \b2v_inst.dir_mem_2Z0Z_6\
        );

    \I__3020\ : CascadeMux
    port map (
            O => \N__19070\,
            I => \b2v_inst.N_489_cascade_\
        );

    \I__3019\ : InMux
    port map (
            O => \N__19067\,
            I => \N__19064\
        );

    \I__3018\ : LocalMux
    port map (
            O => \N__19064\,
            I => \N__19061\
        );

    \I__3017\ : Span4Mux_h
    port map (
            O => \N__19061\,
            I => \N__19056\
        );

    \I__3016\ : InMux
    port map (
            O => \N__19060\,
            I => \N__19053\
        );

    \I__3015\ : InMux
    port map (
            O => \N__19059\,
            I => \N__19050\
        );

    \I__3014\ : Odrv4
    port map (
            O => \N__19056\,
            I => \b2v_inst.un8_dir_mem_2_cry_1_c_RNI88LLZ0\
        );

    \I__3013\ : LocalMux
    port map (
            O => \N__19053\,
            I => \b2v_inst.un8_dir_mem_2_cry_1_c_RNI88LLZ0\
        );

    \I__3012\ : LocalMux
    port map (
            O => \N__19050\,
            I => \b2v_inst.un8_dir_mem_2_cry_1_c_RNI88LLZ0\
        );

    \I__3011\ : InMux
    port map (
            O => \N__19043\,
            I => \N__19040\
        );

    \I__3010\ : LocalMux
    port map (
            O => \N__19040\,
            I => \N__19037\
        );

    \I__3009\ : Span4Mux_h
    port map (
            O => \N__19037\,
            I => \N__19032\
        );

    \I__3008\ : InMux
    port map (
            O => \N__19036\,
            I => \N__19029\
        );

    \I__3007\ : InMux
    port map (
            O => \N__19035\,
            I => \N__19026\
        );

    \I__3006\ : Odrv4
    port map (
            O => \N__19032\,
            I => \b2v_inst.un8_dir_mem_2_cry_2_c_RNIABMLZ0\
        );

    \I__3005\ : LocalMux
    port map (
            O => \N__19029\,
            I => \b2v_inst.un8_dir_mem_2_cry_2_c_RNIABMLZ0\
        );

    \I__3004\ : LocalMux
    port map (
            O => \N__19026\,
            I => \b2v_inst.un8_dir_mem_2_cry_2_c_RNIABMLZ0\
        );

    \I__3003\ : CascadeMux
    port map (
            O => \N__19019\,
            I => \N__19016\
        );

    \I__3002\ : InMux
    port map (
            O => \N__19016\,
            I => \N__19013\
        );

    \I__3001\ : LocalMux
    port map (
            O => \N__19013\,
            I => \N__19010\
        );

    \I__3000\ : Span4Mux_v
    port map (
            O => \N__19010\,
            I => \N__19007\
        );

    \I__2999\ : Odrv4
    port map (
            O => \N__19007\,
            I => \b2v_inst.dir_mem_2Z0Z_4\
        );

    \I__2998\ : InMux
    port map (
            O => \N__19004\,
            I => \N__19001\
        );

    \I__2997\ : LocalMux
    port map (
            O => \N__19001\,
            I => \N__18998\
        );

    \I__2996\ : Span4Mux_h
    port map (
            O => \N__18998\,
            I => \N__18994\
        );

    \I__2995\ : InMux
    port map (
            O => \N__18997\,
            I => \N__18991\
        );

    \I__2994\ : Odrv4
    port map (
            O => \N__18994\,
            I => \b2v_inst.un8_dir_mem_2_cry_3_c_RNICENLZ0\
        );

    \I__2993\ : LocalMux
    port map (
            O => \N__18991\,
            I => \b2v_inst.un8_dir_mem_2_cry_3_c_RNICENLZ0\
        );

    \I__2992\ : InMux
    port map (
            O => \N__18986\,
            I => \N__18983\
        );

    \I__2991\ : LocalMux
    port map (
            O => \N__18983\,
            I => \N__18980\
        );

    \I__2990\ : Span4Mux_v
    port map (
            O => \N__18980\,
            I => \N__18976\
        );

    \I__2989\ : InMux
    port map (
            O => \N__18979\,
            I => \N__18973\
        );

    \I__2988\ : Odrv4
    port map (
            O => \N__18976\,
            I => \b2v_inst.un8_dir_mem_2_cry_4_c_RNIEHOLZ0\
        );

    \I__2987\ : LocalMux
    port map (
            O => \N__18973\,
            I => \b2v_inst.un8_dir_mem_2_cry_4_c_RNIEHOLZ0\
        );

    \I__2986\ : InMux
    port map (
            O => \N__18968\,
            I => \N__18961\
        );

    \I__2985\ : InMux
    port map (
            O => \N__18967\,
            I => \N__18961\
        );

    \I__2984\ : InMux
    port map (
            O => \N__18966\,
            I => \N__18958\
        );

    \I__2983\ : LocalMux
    port map (
            O => \N__18961\,
            I => \N__18953\
        );

    \I__2982\ : LocalMux
    port map (
            O => \N__18958\,
            I => \N__18953\
        );

    \I__2981\ : Odrv12
    port map (
            O => \N__18953\,
            I => \b2v_inst.un8_dir_mem_1_cry_10_THRU_CO\
        );

    \I__2980\ : InMux
    port map (
            O => \N__18950\,
            I => \N__18943\
        );

    \I__2979\ : InMux
    port map (
            O => \N__18949\,
            I => \N__18943\
        );

    \I__2978\ : InMux
    port map (
            O => \N__18948\,
            I => \N__18940\
        );

    \I__2977\ : LocalMux
    port map (
            O => \N__18943\,
            I => \N__18935\
        );

    \I__2976\ : LocalMux
    port map (
            O => \N__18940\,
            I => \N__18935\
        );

    \I__2975\ : Odrv12
    port map (
            O => \N__18935\,
            I => \b2v_inst.un8_dir_mem_1_cry_9_c_RNITCOLZ0\
        );

    \I__2974\ : InMux
    port map (
            O => \N__18932\,
            I => \N__18929\
        );

    \I__2973\ : LocalMux
    port map (
            O => \N__18929\,
            I => \b2v_inst.dir_mem_1Z0Z_8\
        );

    \I__2972\ : CascadeMux
    port map (
            O => \N__18926\,
            I => \N__18923\
        );

    \I__2971\ : InMux
    port map (
            O => \N__18923\,
            I => \N__18920\
        );

    \I__2970\ : LocalMux
    port map (
            O => \N__18920\,
            I => \N__18917\
        );

    \I__2969\ : Odrv4
    port map (
            O => \N__18917\,
            I => \b2v_inst.dir_mem_3Z0Z_8\
        );

    \I__2968\ : InMux
    port map (
            O => \N__18914\,
            I => \N__18911\
        );

    \I__2967\ : LocalMux
    port map (
            O => \N__18911\,
            I => \N__18908\
        );

    \I__2966\ : Span4Mux_h
    port map (
            O => \N__18908\,
            I => \N__18905\
        );

    \I__2965\ : Sp12to4
    port map (
            O => \N__18905\,
            I => \N__18902\
        );

    \I__2964\ : Span12Mux_v
    port map (
            O => \N__18902\,
            I => \N__18899\
        );

    \I__2963\ : Span12Mux_h
    port map (
            O => \N__18899\,
            I => \N__18896\
        );

    \I__2962\ : Odrv12
    port map (
            O => \N__18896\,
            I => swit_c_7
        );

    \I__2961\ : CascadeMux
    port map (
            O => \N__18893\,
            I => \N__18890\
        );

    \I__2960\ : InMux
    port map (
            O => \N__18890\,
            I => \N__18887\
        );

    \I__2959\ : LocalMux
    port map (
            O => \N__18887\,
            I => \N__18884\
        );

    \I__2958\ : Span4Mux_h
    port map (
            O => \N__18884\,
            I => \N__18881\
        );

    \I__2957\ : Span4Mux_h
    port map (
            O => \N__18881\,
            I => \N__18878\
        );

    \I__2956\ : Odrv4
    port map (
            O => \N__18878\,
            I => \b2v_inst.addr_ram_energia_m0_7\
        );

    \I__2955\ : IoInMux
    port map (
            O => \N__18875\,
            I => \N__18871\
        );

    \I__2954\ : InMux
    port map (
            O => \N__18874\,
            I => \N__18868\
        );

    \I__2953\ : LocalMux
    port map (
            O => \N__18871\,
            I => \N__18865\
        );

    \I__2952\ : LocalMux
    port map (
            O => \N__18868\,
            I => \N__18862\
        );

    \I__2951\ : Span4Mux_s3_h
    port map (
            O => \N__18865\,
            I => \N__18859\
        );

    \I__2950\ : Span4Mux_v
    port map (
            O => \N__18862\,
            I => \N__18856\
        );

    \I__2949\ : Span4Mux_h
    port map (
            O => \N__18859\,
            I => \N__18853\
        );

    \I__2948\ : Span4Mux_h
    port map (
            O => \N__18856\,
            I => \N__18850\
        );

    \I__2947\ : Odrv4
    port map (
            O => \N__18853\,
            I => leds_c_12
        );

    \I__2946\ : Odrv4
    port map (
            O => \N__18850\,
            I => leds_c_12
        );

    \I__2945\ : InMux
    port map (
            O => \N__18845\,
            I => \N__18842\
        );

    \I__2944\ : LocalMux
    port map (
            O => \N__18842\,
            I => \N__18838\
        );

    \I__2943\ : InMux
    port map (
            O => \N__18841\,
            I => \N__18835\
        );

    \I__2942\ : Span4Mux_v
    port map (
            O => \N__18838\,
            I => \N__18831\
        );

    \I__2941\ : LocalMux
    port map (
            O => \N__18835\,
            I => \N__18828\
        );

    \I__2940\ : InMux
    port map (
            O => \N__18834\,
            I => \N__18825\
        );

    \I__2939\ : Span4Mux_h
    port map (
            O => \N__18831\,
            I => \N__18820\
        );

    \I__2938\ : Span4Mux_v
    port map (
            O => \N__18828\,
            I => \N__18820\
        );

    \I__2937\ : LocalMux
    port map (
            O => \N__18825\,
            I => \N__18817\
        );

    \I__2936\ : Odrv4
    port map (
            O => \N__18820\,
            I => \b2v_inst.un1_indice_cry_4_c_RNI46NGZ0\
        );

    \I__2935\ : Odrv4
    port map (
            O => \N__18817\,
            I => \b2v_inst.un1_indice_cry_4_c_RNI46NGZ0\
        );

    \I__2934\ : InMux
    port map (
            O => \N__18812\,
            I => \N__18809\
        );

    \I__2933\ : LocalMux
    port map (
            O => \N__18809\,
            I => \N__18805\
        );

    \I__2932\ : InMux
    port map (
            O => \N__18808\,
            I => \N__18802\
        );

    \I__2931\ : Span4Mux_v
    port map (
            O => \N__18805\,
            I => \N__18797\
        );

    \I__2930\ : LocalMux
    port map (
            O => \N__18802\,
            I => \N__18797\
        );

    \I__2929\ : Span4Mux_h
    port map (
            O => \N__18797\,
            I => \N__18793\
        );

    \I__2928\ : InMux
    port map (
            O => \N__18796\,
            I => \N__18790\
        );

    \I__2927\ : Odrv4
    port map (
            O => \N__18793\,
            I => \b2v_inst.un1_indice_cry_8_c_RNICIRGZ0\
        );

    \I__2926\ : LocalMux
    port map (
            O => \N__18790\,
            I => \b2v_inst.un1_indice_cry_8_c_RNICIRGZ0\
        );

    \I__2925\ : InMux
    port map (
            O => \N__18785\,
            I => \N__18781\
        );

    \I__2924\ : InMux
    port map (
            O => \N__18784\,
            I => \N__18777\
        );

    \I__2923\ : LocalMux
    port map (
            O => \N__18781\,
            I => \N__18774\
        );

    \I__2922\ : CascadeMux
    port map (
            O => \N__18780\,
            I => \N__18771\
        );

    \I__2921\ : LocalMux
    port map (
            O => \N__18777\,
            I => \N__18768\
        );

    \I__2920\ : Span4Mux_h
    port map (
            O => \N__18774\,
            I => \N__18765\
        );

    \I__2919\ : InMux
    port map (
            O => \N__18771\,
            I => \N__18762\
        );

    \I__2918\ : Span4Mux_h
    port map (
            O => \N__18768\,
            I => \N__18759\
        );

    \I__2917\ : Span4Mux_h
    port map (
            O => \N__18765\,
            I => \N__18754\
        );

    \I__2916\ : LocalMux
    port map (
            O => \N__18762\,
            I => \N__18754\
        );

    \I__2915\ : Odrv4
    port map (
            O => \N__18759\,
            I => \b2v_inst.dir_mem_316lto7\
        );

    \I__2914\ : Odrv4
    port map (
            O => \N__18754\,
            I => \b2v_inst.dir_mem_316lto7\
        );

    \I__2913\ : InMux
    port map (
            O => \N__18749\,
            I => \N__18746\
        );

    \I__2912\ : LocalMux
    port map (
            O => \N__18746\,
            I => \N__18743\
        );

    \I__2911\ : Span4Mux_h
    port map (
            O => \N__18743\,
            I => \N__18740\
        );

    \I__2910\ : Sp12to4
    port map (
            O => \N__18740\,
            I => \N__18737\
        );

    \I__2909\ : Span12Mux_v
    port map (
            O => \N__18737\,
            I => \N__18734\
        );

    \I__2908\ : Span12Mux_h
    port map (
            O => \N__18734\,
            I => \N__18731\
        );

    \I__2907\ : Odrv12
    port map (
            O => \N__18731\,
            I => swit_c_6
        );

    \I__2906\ : CascadeMux
    port map (
            O => \N__18728\,
            I => \b2v_inst.addr_ram_energia_m0_6_cascade_\
        );

    \I__2905\ : CascadeMux
    port map (
            O => \N__18725\,
            I => \N__18721\
        );

    \I__2904\ : CascadeMux
    port map (
            O => \N__18724\,
            I => \N__18718\
        );

    \I__2903\ : CascadeBuf
    port map (
            O => \N__18721\,
            I => \N__18715\
        );

    \I__2902\ : CascadeBuf
    port map (
            O => \N__18718\,
            I => \N__18712\
        );

    \I__2901\ : CascadeMux
    port map (
            O => \N__18715\,
            I => \N__18709\
        );

    \I__2900\ : CascadeMux
    port map (
            O => \N__18712\,
            I => \N__18706\
        );

    \I__2899\ : CascadeBuf
    port map (
            O => \N__18709\,
            I => \N__18703\
        );

    \I__2898\ : CascadeBuf
    port map (
            O => \N__18706\,
            I => \N__18700\
        );

    \I__2897\ : CascadeMux
    port map (
            O => \N__18703\,
            I => \N__18697\
        );

    \I__2896\ : CascadeMux
    port map (
            O => \N__18700\,
            I => \N__18694\
        );

    \I__2895\ : CascadeBuf
    port map (
            O => \N__18697\,
            I => \N__18691\
        );

    \I__2894\ : CascadeBuf
    port map (
            O => \N__18694\,
            I => \N__18688\
        );

    \I__2893\ : CascadeMux
    port map (
            O => \N__18691\,
            I => \N__18685\
        );

    \I__2892\ : CascadeMux
    port map (
            O => \N__18688\,
            I => \N__18682\
        );

    \I__2891\ : CascadeBuf
    port map (
            O => \N__18685\,
            I => \N__18679\
        );

    \I__2890\ : CascadeBuf
    port map (
            O => \N__18682\,
            I => \N__18676\
        );

    \I__2889\ : CascadeMux
    port map (
            O => \N__18679\,
            I => \N__18673\
        );

    \I__2888\ : CascadeMux
    port map (
            O => \N__18676\,
            I => \N__18670\
        );

    \I__2887\ : CascadeBuf
    port map (
            O => \N__18673\,
            I => \N__18667\
        );

    \I__2886\ : CascadeBuf
    port map (
            O => \N__18670\,
            I => \N__18664\
        );

    \I__2885\ : CascadeMux
    port map (
            O => \N__18667\,
            I => \N__18661\
        );

    \I__2884\ : CascadeMux
    port map (
            O => \N__18664\,
            I => \N__18658\
        );

    \I__2883\ : CascadeBuf
    port map (
            O => \N__18661\,
            I => \N__18655\
        );

    \I__2882\ : CascadeBuf
    port map (
            O => \N__18658\,
            I => \N__18652\
        );

    \I__2881\ : CascadeMux
    port map (
            O => \N__18655\,
            I => \N__18649\
        );

    \I__2880\ : CascadeMux
    port map (
            O => \N__18652\,
            I => \N__18646\
        );

    \I__2879\ : InMux
    port map (
            O => \N__18649\,
            I => \N__18643\
        );

    \I__2878\ : InMux
    port map (
            O => \N__18646\,
            I => \N__18640\
        );

    \I__2877\ : LocalMux
    port map (
            O => \N__18643\,
            I => \N__18635\
        );

    \I__2876\ : LocalMux
    port map (
            O => \N__18640\,
            I => \N__18635\
        );

    \I__2875\ : Span12Mux_s11_v
    port map (
            O => \N__18635\,
            I => \N__18632\
        );

    \I__2874\ : Odrv12
    port map (
            O => \N__18632\,
            I => \SYNTHESIZED_WIRE_12_6\
        );

    \I__2873\ : InMux
    port map (
            O => \N__18629\,
            I => \N__18626\
        );

    \I__2872\ : LocalMux
    port map (
            O => \N__18626\,
            I => \N__18623\
        );

    \I__2871\ : Odrv4
    port map (
            O => \N__18623\,
            I => \b2v_inst.state_ns_0_i_a2_0_0_23\
        );

    \I__2870\ : CascadeMux
    port map (
            O => \N__18620\,
            I => \b2v_inst.state_ns_i_0_a2_11_o2_4_0_6_1_3_cascade_\
        );

    \I__2869\ : InMux
    port map (
            O => \N__18617\,
            I => \N__18614\
        );

    \I__2868\ : LocalMux
    port map (
            O => \N__18614\,
            I => \b2v_inst.state_ns_i_0_a2_11_o2_4_0_1_3\
        );

    \I__2867\ : InMux
    port map (
            O => \N__18611\,
            I => \N__18608\
        );

    \I__2866\ : LocalMux
    port map (
            O => \N__18608\,
            I => \N__18605\
        );

    \I__2865\ : Odrv12
    port map (
            O => \N__18605\,
            I => \b2v_inst.N_11\
        );

    \I__2864\ : CascadeMux
    port map (
            O => \N__18602\,
            I => \b2v_inst.N_4_i_i_1_cascade_\
        );

    \I__2863\ : InMux
    port map (
            O => \N__18599\,
            I => \N__18596\
        );

    \I__2862\ : LocalMux
    port map (
            O => \N__18596\,
            I => \b2v_inst.g3_i_1\
        );

    \I__2861\ : InMux
    port map (
            O => \N__18593\,
            I => \N__18590\
        );

    \I__2860\ : LocalMux
    port map (
            O => \N__18590\,
            I => \N__18587\
        );

    \I__2859\ : Span4Mux_v
    port map (
            O => \N__18587\,
            I => \N__18584\
        );

    \I__2858\ : Sp12to4
    port map (
            O => \N__18584\,
            I => \N__18581\
        );

    \I__2857\ : Span12Mux_h
    port map (
            O => \N__18581\,
            I => \N__18578\
        );

    \I__2856\ : Span12Mux_h
    port map (
            O => \N__18578\,
            I => \N__18575\
        );

    \I__2855\ : Span12Mux_v
    port map (
            O => \N__18575\,
            I => \N__18572\
        );

    \I__2854\ : Odrv12
    port map (
            O => \N__18572\,
            I => swit_c_8
        );

    \I__2853\ : InMux
    port map (
            O => \N__18569\,
            I => \N__18566\
        );

    \I__2852\ : LocalMux
    port map (
            O => \N__18566\,
            I => \N__18563\
        );

    \I__2851\ : Span12Mux_v
    port map (
            O => \N__18563\,
            I => \N__18560\
        );

    \I__2850\ : Odrv12
    port map (
            O => \N__18560\,
            I => \b2v_inst.addr_ram_energia_m0_8\
        );

    \I__2849\ : InMux
    port map (
            O => \N__18557\,
            I => \N__18554\
        );

    \I__2848\ : LocalMux
    port map (
            O => \N__18554\,
            I => \b2v_inst.state_ns_i_0_a2_11_o2_4_0_5_3\
        );

    \I__2847\ : InMux
    port map (
            O => \N__18551\,
            I => \N__18548\
        );

    \I__2846\ : LocalMux
    port map (
            O => \N__18548\,
            I => \b2v_inst.state_RNO_2Z0Z_29\
        );

    \I__2845\ : CascadeMux
    port map (
            O => \N__18545\,
            I => \b2v_inst.state_ns_i_0_a2_11_o2_4_0_7_3_cascade_\
        );

    \I__2844\ : InMux
    port map (
            O => \N__18542\,
            I => \N__18539\
        );

    \I__2843\ : LocalMux
    port map (
            O => \N__18539\,
            I => \N__18536\
        );

    \I__2842\ : Odrv4
    port map (
            O => \N__18536\,
            I => \b2v_inst.state_RNO_1Z0Z_29\
        );

    \I__2841\ : InMux
    port map (
            O => \N__18533\,
            I => \N__18530\
        );

    \I__2840\ : LocalMux
    port map (
            O => \N__18530\,
            I => \b2v_inst.dir_energia_RNO_0Z0Z_0\
        );

    \I__2839\ : CascadeMux
    port map (
            O => \N__18527\,
            I => \N__18524\
        );

    \I__2838\ : InMux
    port map (
            O => \N__18524\,
            I => \N__18521\
        );

    \I__2837\ : LocalMux
    port map (
            O => \N__18521\,
            I => \N__18518\
        );

    \I__2836\ : Span4Mux_h
    port map (
            O => \N__18518\,
            I => \N__18515\
        );

    \I__2835\ : Odrv4
    port map (
            O => \N__18515\,
            I => \b2v_inst.dir_mem_3Z0Z_5\
        );

    \I__2834\ : CascadeMux
    port map (
            O => \N__18512\,
            I => \N__18509\
        );

    \I__2833\ : InMux
    port map (
            O => \N__18509\,
            I => \N__18506\
        );

    \I__2832\ : LocalMux
    port map (
            O => \N__18506\,
            I => \N__18503\
        );

    \I__2831\ : Span4Mux_v
    port map (
            O => \N__18503\,
            I => \N__18500\
        );

    \I__2830\ : Span4Mux_h
    port map (
            O => \N__18500\,
            I => \N__18497\
        );

    \I__2829\ : Span4Mux_h
    port map (
            O => \N__18497\,
            I => \N__18494\
        );

    \I__2828\ : Span4Mux_h
    port map (
            O => \N__18494\,
            I => \N__18491\
        );

    \I__2827\ : Odrv4
    port map (
            O => \N__18491\,
            I => \SYNTHESIZED_WIRE_1_5\
        );

    \I__2826\ : InMux
    port map (
            O => \N__18488\,
            I => \N__18485\
        );

    \I__2825\ : LocalMux
    port map (
            O => \N__18485\,
            I => \N__18482\
        );

    \I__2824\ : Span4Mux_h
    port map (
            O => \N__18482\,
            I => \N__18479\
        );

    \I__2823\ : Odrv4
    port map (
            O => \N__18479\,
            I => \b2v_inst.dir_memZ0Z_4\
        );

    \I__2822\ : CascadeMux
    port map (
            O => \N__18476\,
            I => \b2v_inst.addr_ram_iv_i_0_4_cascade_\
        );

    \I__2821\ : CascadeMux
    port map (
            O => \N__18473\,
            I => \N__18470\
        );

    \I__2820\ : CascadeBuf
    port map (
            O => \N__18470\,
            I => \N__18466\
        );

    \I__2819\ : CascadeMux
    port map (
            O => \N__18469\,
            I => \N__18463\
        );

    \I__2818\ : CascadeMux
    port map (
            O => \N__18466\,
            I => \N__18460\
        );

    \I__2817\ : CascadeBuf
    port map (
            O => \N__18463\,
            I => \N__18457\
        );

    \I__2816\ : CascadeBuf
    port map (
            O => \N__18460\,
            I => \N__18454\
        );

    \I__2815\ : CascadeMux
    port map (
            O => \N__18457\,
            I => \N__18451\
        );

    \I__2814\ : CascadeMux
    port map (
            O => \N__18454\,
            I => \N__18448\
        );

    \I__2813\ : CascadeBuf
    port map (
            O => \N__18451\,
            I => \N__18445\
        );

    \I__2812\ : CascadeBuf
    port map (
            O => \N__18448\,
            I => \N__18442\
        );

    \I__2811\ : CascadeMux
    port map (
            O => \N__18445\,
            I => \N__18439\
        );

    \I__2810\ : CascadeMux
    port map (
            O => \N__18442\,
            I => \N__18436\
        );

    \I__2809\ : CascadeBuf
    port map (
            O => \N__18439\,
            I => \N__18433\
        );

    \I__2808\ : CascadeBuf
    port map (
            O => \N__18436\,
            I => \N__18430\
        );

    \I__2807\ : CascadeMux
    port map (
            O => \N__18433\,
            I => \N__18427\
        );

    \I__2806\ : CascadeMux
    port map (
            O => \N__18430\,
            I => \N__18424\
        );

    \I__2805\ : CascadeBuf
    port map (
            O => \N__18427\,
            I => \N__18421\
        );

    \I__2804\ : CascadeBuf
    port map (
            O => \N__18424\,
            I => \N__18418\
        );

    \I__2803\ : CascadeMux
    port map (
            O => \N__18421\,
            I => \N__18415\
        );

    \I__2802\ : CascadeMux
    port map (
            O => \N__18418\,
            I => \N__18412\
        );

    \I__2801\ : CascadeBuf
    port map (
            O => \N__18415\,
            I => \N__18409\
        );

    \I__2800\ : InMux
    port map (
            O => \N__18412\,
            I => \N__18406\
        );

    \I__2799\ : CascadeMux
    port map (
            O => \N__18409\,
            I => \N__18403\
        );

    \I__2798\ : LocalMux
    port map (
            O => \N__18406\,
            I => \N__18400\
        );

    \I__2797\ : InMux
    port map (
            O => \N__18403\,
            I => \N__18397\
        );

    \I__2796\ : Span4Mux_h
    port map (
            O => \N__18400\,
            I => \N__18394\
        );

    \I__2795\ : LocalMux
    port map (
            O => \N__18397\,
            I => \N__18391\
        );

    \I__2794\ : Span4Mux_h
    port map (
            O => \N__18394\,
            I => \N__18388\
        );

    \I__2793\ : Span12Mux_s11_h
    port map (
            O => \N__18391\,
            I => \N__18385\
        );

    \I__2792\ : Span4Mux_h
    port map (
            O => \N__18388\,
            I => \N__18382\
        );

    \I__2791\ : Odrv12
    port map (
            O => \N__18385\,
            I => \indice_RNIN3333_4\
        );

    \I__2790\ : Odrv4
    port map (
            O => \N__18382\,
            I => \indice_RNIN3333_4\
        );

    \I__2789\ : InMux
    port map (
            O => \N__18377\,
            I => \N__18374\
        );

    \I__2788\ : LocalMux
    port map (
            O => \N__18374\,
            I => \N__18371\
        );

    \I__2787\ : Odrv12
    port map (
            O => \N__18371\,
            I => \b2v_inst.dir_mem_1Z0Z_4\
        );

    \I__2786\ : InMux
    port map (
            O => \N__18368\,
            I => \N__18365\
        );

    \I__2785\ : LocalMux
    port map (
            O => \N__18365\,
            I => \b2v_inst.addr_ram_iv_i_1_4\
        );

    \I__2784\ : InMux
    port map (
            O => \N__18362\,
            I => \N__18358\
        );

    \I__2783\ : InMux
    port map (
            O => \N__18361\,
            I => \N__18355\
        );

    \I__2782\ : LocalMux
    port map (
            O => \N__18358\,
            I => \N__18352\
        );

    \I__2781\ : LocalMux
    port map (
            O => \N__18355\,
            I => \N__18348\
        );

    \I__2780\ : Span4Mux_v
    port map (
            O => \N__18352\,
            I => \N__18345\
        );

    \I__2779\ : InMux
    port map (
            O => \N__18351\,
            I => \N__18342\
        );

    \I__2778\ : Span4Mux_h
    port map (
            O => \N__18348\,
            I => \N__18335\
        );

    \I__2777\ : Span4Mux_h
    port map (
            O => \N__18345\,
            I => \N__18335\
        );

    \I__2776\ : LocalMux
    port map (
            O => \N__18342\,
            I => \N__18335\
        );

    \I__2775\ : Odrv4
    port map (
            O => \N__18335\,
            I => \b2v_inst.un1_indice_cry_3_c_RNI23MGZ0\
        );

    \I__2774\ : CascadeMux
    port map (
            O => \N__18332\,
            I => \N__18329\
        );

    \I__2773\ : InMux
    port map (
            O => \N__18329\,
            I => \N__18326\
        );

    \I__2772\ : LocalMux
    port map (
            O => \N__18326\,
            I => \N__18319\
        );

    \I__2771\ : CascadeMux
    port map (
            O => \N__18325\,
            I => \N__18315\
        );

    \I__2770\ : CascadeMux
    port map (
            O => \N__18324\,
            I => \N__18310\
        );

    \I__2769\ : CascadeMux
    port map (
            O => \N__18323\,
            I => \N__18307\
        );

    \I__2768\ : CascadeMux
    port map (
            O => \N__18322\,
            I => \N__18303\
        );

    \I__2767\ : Span4Mux_h
    port map (
            O => \N__18319\,
            I => \N__18300\
        );

    \I__2766\ : InMux
    port map (
            O => \N__18318\,
            I => \N__18295\
        );

    \I__2765\ : InMux
    port map (
            O => \N__18315\,
            I => \N__18295\
        );

    \I__2764\ : InMux
    port map (
            O => \N__18314\,
            I => \N__18288\
        );

    \I__2763\ : InMux
    port map (
            O => \N__18313\,
            I => \N__18288\
        );

    \I__2762\ : InMux
    port map (
            O => \N__18310\,
            I => \N__18288\
        );

    \I__2761\ : InMux
    port map (
            O => \N__18307\,
            I => \N__18285\
        );

    \I__2760\ : InMux
    port map (
            O => \N__18306\,
            I => \N__18280\
        );

    \I__2759\ : InMux
    port map (
            O => \N__18303\,
            I => \N__18280\
        );

    \I__2758\ : Odrv4
    port map (
            O => \N__18300\,
            I => \b2v_inst.dir_mem_316lto11_0\
        );

    \I__2757\ : LocalMux
    port map (
            O => \N__18295\,
            I => \b2v_inst.dir_mem_316lto11_0\
        );

    \I__2756\ : LocalMux
    port map (
            O => \N__18288\,
            I => \b2v_inst.dir_mem_316lto11_0\
        );

    \I__2755\ : LocalMux
    port map (
            O => \N__18285\,
            I => \b2v_inst.dir_mem_316lto11_0\
        );

    \I__2754\ : LocalMux
    port map (
            O => \N__18280\,
            I => \b2v_inst.dir_mem_316lto11_0\
        );

    \I__2753\ : InMux
    port map (
            O => \N__18269\,
            I => \N__18266\
        );

    \I__2752\ : LocalMux
    port map (
            O => \N__18266\,
            I => \N__18263\
        );

    \I__2751\ : Span4Mux_v
    port map (
            O => \N__18263\,
            I => \N__18250\
        );

    \I__2750\ : InMux
    port map (
            O => \N__18262\,
            I => \N__18247\
        );

    \I__2749\ : InMux
    port map (
            O => \N__18261\,
            I => \N__18242\
        );

    \I__2748\ : InMux
    port map (
            O => \N__18260\,
            I => \N__18242\
        );

    \I__2747\ : InMux
    port map (
            O => \N__18259\,
            I => \N__18227\
        );

    \I__2746\ : InMux
    port map (
            O => \N__18258\,
            I => \N__18227\
        );

    \I__2745\ : InMux
    port map (
            O => \N__18257\,
            I => \N__18227\
        );

    \I__2744\ : InMux
    port map (
            O => \N__18256\,
            I => \N__18227\
        );

    \I__2743\ : InMux
    port map (
            O => \N__18255\,
            I => \N__18227\
        );

    \I__2742\ : InMux
    port map (
            O => \N__18254\,
            I => \N__18227\
        );

    \I__2741\ : InMux
    port map (
            O => \N__18253\,
            I => \N__18227\
        );

    \I__2740\ : Odrv4
    port map (
            O => \N__18250\,
            I => \b2v_inst.dir_mem_316lt11\
        );

    \I__2739\ : LocalMux
    port map (
            O => \N__18247\,
            I => \b2v_inst.dir_mem_316lt11\
        );

    \I__2738\ : LocalMux
    port map (
            O => \N__18242\,
            I => \b2v_inst.dir_mem_316lt11\
        );

    \I__2737\ : LocalMux
    port map (
            O => \N__18227\,
            I => \b2v_inst.dir_mem_316lt11\
        );

    \I__2736\ : CascadeMux
    port map (
            O => \N__18218\,
            I => \N__18215\
        );

    \I__2735\ : InMux
    port map (
            O => \N__18215\,
            I => \N__18212\
        );

    \I__2734\ : LocalMux
    port map (
            O => \N__18212\,
            I => \b2v_inst.dir_mem_3Z0Z_4\
        );

    \I__2733\ : CEMux
    port map (
            O => \N__18209\,
            I => \N__18205\
        );

    \I__2732\ : CEMux
    port map (
            O => \N__18208\,
            I => \N__18200\
        );

    \I__2731\ : LocalMux
    port map (
            O => \N__18205\,
            I => \N__18197\
        );

    \I__2730\ : CEMux
    port map (
            O => \N__18204\,
            I => \N__18194\
        );

    \I__2729\ : CEMux
    port map (
            O => \N__18203\,
            I => \N__18191\
        );

    \I__2728\ : LocalMux
    port map (
            O => \N__18200\,
            I => \N__18188\
        );

    \I__2727\ : Span4Mux_v
    port map (
            O => \N__18197\,
            I => \N__18183\
        );

    \I__2726\ : LocalMux
    port map (
            O => \N__18194\,
            I => \N__18183\
        );

    \I__2725\ : LocalMux
    port map (
            O => \N__18191\,
            I => \N__18180\
        );

    \I__2724\ : Span4Mux_h
    port map (
            O => \N__18188\,
            I => \N__18177\
        );

    \I__2723\ : Sp12to4
    port map (
            O => \N__18183\,
            I => \N__18174\
        );

    \I__2722\ : Odrv4
    port map (
            O => \N__18180\,
            I => \b2v_inst.N_362_i\
        );

    \I__2721\ : Odrv4
    port map (
            O => \N__18177\,
            I => \b2v_inst.N_362_i\
        );

    \I__2720\ : Odrv12
    port map (
            O => \N__18174\,
            I => \b2v_inst.N_362_i\
        );

    \I__2719\ : InMux
    port map (
            O => \N__18167\,
            I => \N__18161\
        );

    \I__2718\ : InMux
    port map (
            O => \N__18166\,
            I => \N__18161\
        );

    \I__2717\ : LocalMux
    port map (
            O => \N__18161\,
            I => \N__18158\
        );

    \I__2716\ : Odrv12
    port map (
            O => \N__18158\,
            I => \b2v_inst.un8_dir_mem_1_cry_7_c_RNIIHVCZ0\
        );

    \I__2715\ : CascadeMux
    port map (
            O => \N__18155\,
            I => \N__18152\
        );

    \I__2714\ : InMux
    port map (
            O => \N__18152\,
            I => \N__18149\
        );

    \I__2713\ : LocalMux
    port map (
            O => \N__18149\,
            I => \N__18146\
        );

    \I__2712\ : Span4Mux_h
    port map (
            O => \N__18146\,
            I => \N__18143\
        );

    \I__2711\ : Odrv4
    port map (
            O => \N__18143\,
            I => \b2v_inst.dir_mem_1_RNO_0Z0Z_8\
        );

    \I__2710\ : InMux
    port map (
            O => \N__18140\,
            I => \N__18134\
        );

    \I__2709\ : InMux
    port map (
            O => \N__18139\,
            I => \N__18134\
        );

    \I__2708\ : LocalMux
    port map (
            O => \N__18134\,
            I => \N__18131\
        );

    \I__2707\ : Odrv4
    port map (
            O => \N__18131\,
            I => \b2v_inst.un8_dir_mem_1_cry_8_c_RNIKK0DZ0\
        );

    \I__2706\ : CascadeMux
    port map (
            O => \N__18128\,
            I => \N__18125\
        );

    \I__2705\ : InMux
    port map (
            O => \N__18125\,
            I => \N__18122\
        );

    \I__2704\ : LocalMux
    port map (
            O => \N__18122\,
            I => \N__18119\
        );

    \I__2703\ : Span4Mux_h
    port map (
            O => \N__18119\,
            I => \N__18116\
        );

    \I__2702\ : Odrv4
    port map (
            O => \N__18116\,
            I => \b2v_inst.dir_mem_1_RNO_0Z0Z_9\
        );

    \I__2701\ : InMux
    port map (
            O => \N__18113\,
            I => \N__18109\
        );

    \I__2700\ : InMux
    port map (
            O => \N__18112\,
            I => \N__18106\
        );

    \I__2699\ : LocalMux
    port map (
            O => \N__18109\,
            I => \N__18103\
        );

    \I__2698\ : LocalMux
    port map (
            O => \N__18106\,
            I => \N__18100\
        );

    \I__2697\ : Span4Mux_v
    port map (
            O => \N__18103\,
            I => \N__18097\
        );

    \I__2696\ : Span4Mux_v
    port map (
            O => \N__18100\,
            I => \N__18094\
        );

    \I__2695\ : Odrv4
    port map (
            O => \N__18097\,
            I => \b2v_inst.un8_dir_mem_1_cry_4_c_RNIC8SCZ0\
        );

    \I__2694\ : Odrv4
    port map (
            O => \N__18094\,
            I => \b2v_inst.un8_dir_mem_1_cry_4_c_RNIC8SCZ0\
        );

    \I__2693\ : CascadeMux
    port map (
            O => \N__18089\,
            I => \N__18086\
        );

    \I__2692\ : InMux
    port map (
            O => \N__18086\,
            I => \N__18083\
        );

    \I__2691\ : LocalMux
    port map (
            O => \N__18083\,
            I => \N__18080\
        );

    \I__2690\ : Span4Mux_h
    port map (
            O => \N__18080\,
            I => \N__18077\
        );

    \I__2689\ : Odrv4
    port map (
            O => \N__18077\,
            I => \b2v_inst.dir_mem_1_RNO_0Z0Z_5\
        );

    \I__2688\ : InMux
    port map (
            O => \N__18074\,
            I => \N__18071\
        );

    \I__2687\ : LocalMux
    port map (
            O => \N__18071\,
            I => \N__18068\
        );

    \I__2686\ : Odrv4
    port map (
            O => \N__18068\,
            I => \b2v_inst.dir_mem_1Z0Z_6\
        );

    \I__2685\ : CascadeMux
    port map (
            O => \N__18065\,
            I => \N__18062\
        );

    \I__2684\ : InMux
    port map (
            O => \N__18062\,
            I => \N__18059\
        );

    \I__2683\ : LocalMux
    port map (
            O => \N__18059\,
            I => \N__18056\
        );

    \I__2682\ : Span4Mux_v
    port map (
            O => \N__18056\,
            I => \N__18053\
        );

    \I__2681\ : Odrv4
    port map (
            O => \N__18053\,
            I => \b2v_inst.dir_mem_3Z0Z_6\
        );

    \I__2680\ : InMux
    port map (
            O => \N__18050\,
            I => \N__18047\
        );

    \I__2679\ : LocalMux
    port map (
            O => \N__18047\,
            I => \N__18044\
        );

    \I__2678\ : Odrv4
    port map (
            O => \N__18044\,
            I => \b2v_inst.dir_memZ0Z_7\
        );

    \I__2677\ : CascadeMux
    port map (
            O => \N__18041\,
            I => \b2v_inst.N_450_i_1_cascade_\
        );

    \I__2676\ : InMux
    port map (
            O => \N__18038\,
            I => \N__18035\
        );

    \I__2675\ : LocalMux
    port map (
            O => \N__18035\,
            I => \N__18032\
        );

    \I__2674\ : Span4Mux_h
    port map (
            O => \N__18032\,
            I => \N__18029\
        );

    \I__2673\ : Odrv4
    port map (
            O => \N__18029\,
            I => \b2v_inst.dir_memZ0Z_10\
        );

    \I__2672\ : InMux
    port map (
            O => \N__18026\,
            I => \N__18023\
        );

    \I__2671\ : LocalMux
    port map (
            O => \N__18023\,
            I => \N__18020\
        );

    \I__2670\ : Odrv4
    port map (
            O => \N__18020\,
            I => \b2v_inst.dir_mem_1Z0Z_5\
        );

    \I__2669\ : InMux
    port map (
            O => \N__18017\,
            I => \N__18014\
        );

    \I__2668\ : LocalMux
    port map (
            O => \N__18014\,
            I => \N__18010\
        );

    \I__2667\ : InMux
    port map (
            O => \N__18013\,
            I => \N__18007\
        );

    \I__2666\ : Odrv4
    port map (
            O => \N__18010\,
            I => \b2v_inst.un8_dir_mem_1_cry_2_c_RNI82QCZ0\
        );

    \I__2665\ : LocalMux
    port map (
            O => \N__18007\,
            I => \b2v_inst.un8_dir_mem_1_cry_2_c_RNI82QCZ0\
        );

    \I__2664\ : InMux
    port map (
            O => \N__18002\,
            I => \N__17999\
        );

    \I__2663\ : LocalMux
    port map (
            O => \N__17999\,
            I => \N__17995\
        );

    \I__2662\ : InMux
    port map (
            O => \N__17998\,
            I => \N__17992\
        );

    \I__2661\ : Odrv4
    port map (
            O => \N__17995\,
            I => \b2v_inst.un8_dir_mem_1_cry_3_c_RNIA5RCZ0\
        );

    \I__2660\ : LocalMux
    port map (
            O => \N__17992\,
            I => \b2v_inst.un8_dir_mem_1_cry_3_c_RNIA5RCZ0\
        );

    \I__2659\ : InMux
    port map (
            O => \N__17987\,
            I => \N__17983\
        );

    \I__2658\ : InMux
    port map (
            O => \N__17986\,
            I => \N__17980\
        );

    \I__2657\ : LocalMux
    port map (
            O => \N__17983\,
            I => \N__17977\
        );

    \I__2656\ : LocalMux
    port map (
            O => \N__17980\,
            I => \N__17974\
        );

    \I__2655\ : Span4Mux_h
    port map (
            O => \N__17977\,
            I => \N__17971\
        );

    \I__2654\ : Odrv12
    port map (
            O => \N__17974\,
            I => \b2v_inst.un8_dir_mem_1_cry_5_c_RNIEBTCZ0\
        );

    \I__2653\ : Odrv4
    port map (
            O => \N__17971\,
            I => \b2v_inst.un8_dir_mem_1_cry_5_c_RNIEBTCZ0\
        );

    \I__2652\ : CascadeMux
    port map (
            O => \N__17966\,
            I => \N__17963\
        );

    \I__2651\ : InMux
    port map (
            O => \N__17963\,
            I => \N__17960\
        );

    \I__2650\ : LocalMux
    port map (
            O => \N__17960\,
            I => \N__17957\
        );

    \I__2649\ : Sp12to4
    port map (
            O => \N__17957\,
            I => \N__17954\
        );

    \I__2648\ : Span12Mux_s10_v
    port map (
            O => \N__17954\,
            I => \N__17951\
        );

    \I__2647\ : Odrv12
    port map (
            O => \N__17951\,
            I => \b2v_inst.dir_mem_1_RNO_0Z0Z_6\
        );

    \I__2646\ : InMux
    port map (
            O => \N__17948\,
            I => \N__17945\
        );

    \I__2645\ : LocalMux
    port map (
            O => \N__17945\,
            I => \b2v_inst.dir_mem_215lt7\
        );

    \I__2644\ : InMux
    port map (
            O => \N__17942\,
            I => \N__17939\
        );

    \I__2643\ : LocalMux
    port map (
            O => \N__17939\,
            I => \b2v_inst.dir_mem_115lt7\
        );

    \I__2642\ : InMux
    port map (
            O => \N__17936\,
            I => \N__17933\
        );

    \I__2641\ : LocalMux
    port map (
            O => \N__17933\,
            I => \N__17930\
        );

    \I__2640\ : Span4Mux_h
    port map (
            O => \N__17930\,
            I => \N__17927\
        );

    \I__2639\ : Odrv4
    port map (
            O => \N__17927\,
            I => \b2v_inst.dir_mem_1_RNO_0Z0Z_10\
        );

    \I__2638\ : CascadeMux
    port map (
            O => \N__17924\,
            I => \b2v_inst.dir_mem_115lt11_cascade_\
        );

    \I__2637\ : CascadeMux
    port map (
            O => \N__17921\,
            I => \N__17917\
        );

    \I__2636\ : InMux
    port map (
            O => \N__17920\,
            I => \N__17914\
        );

    \I__2635\ : InMux
    port map (
            O => \N__17917\,
            I => \N__17911\
        );

    \I__2634\ : LocalMux
    port map (
            O => \N__17914\,
            I => \N__17906\
        );

    \I__2633\ : LocalMux
    port map (
            O => \N__17911\,
            I => \N__17906\
        );

    \I__2632\ : Span4Mux_h
    port map (
            O => \N__17906\,
            I => \N__17903\
        );

    \I__2631\ : Odrv4
    port map (
            O => \N__17903\,
            I => \b2v_inst.dir_mem_115lto7\
        );

    \I__2630\ : CascadeMux
    port map (
            O => \N__17900\,
            I => \N__17897\
        );

    \I__2629\ : InMux
    port map (
            O => \N__17897\,
            I => \N__17894\
        );

    \I__2628\ : LocalMux
    port map (
            O => \N__17894\,
            I => \N__17891\
        );

    \I__2627\ : Span4Mux_h
    port map (
            O => \N__17891\,
            I => \N__17888\
        );

    \I__2626\ : Odrv4
    port map (
            O => \N__17888\,
            I => \b2v_inst.dir_mem_1_RNO_0Z0Z_7\
        );

    \I__2625\ : CascadeMux
    port map (
            O => \N__17885\,
            I => \b2v_inst.N_512_cascade_\
        );

    \I__2624\ : InMux
    port map (
            O => \N__17882\,
            I => \N__17879\
        );

    \I__2623\ : LocalMux
    port map (
            O => \N__17879\,
            I => \N__17876\
        );

    \I__2622\ : Odrv4
    port map (
            O => \N__17876\,
            I => \b2v_inst.N_430_tz\
        );

    \I__2621\ : CascadeMux
    port map (
            O => \N__17873\,
            I => \b2v_inst.g0_4_4_cascade_\
        );

    \I__2620\ : InMux
    port map (
            O => \N__17870\,
            I => \N__17867\
        );

    \I__2619\ : LocalMux
    port map (
            O => \N__17867\,
            I => \N__17864\
        );

    \I__2618\ : Odrv12
    port map (
            O => \N__17864\,
            I => \b2v_inst.g3_0_0\
        );

    \I__2617\ : CascadeMux
    port map (
            O => \N__17861\,
            I => \N__17858\
        );

    \I__2616\ : InMux
    port map (
            O => \N__17858\,
            I => \N__17854\
        );

    \I__2615\ : InMux
    port map (
            O => \N__17857\,
            I => \N__17851\
        );

    \I__2614\ : LocalMux
    port map (
            O => \N__17854\,
            I => \N__17848\
        );

    \I__2613\ : LocalMux
    port map (
            O => \N__17851\,
            I => \N__17843\
        );

    \I__2612\ : Span4Mux_v
    port map (
            O => \N__17848\,
            I => \N__17843\
        );

    \I__2611\ : Odrv4
    port map (
            O => \N__17843\,
            I => \b2v_inst.un4_pix_count_intlto18Z0Z_0\
        );

    \I__2610\ : CascadeMux
    port map (
            O => \N__17840\,
            I => \b2v_inst.g0_0_cascade_\
        );

    \I__2609\ : InMux
    port map (
            O => \N__17837\,
            I => \N__17834\
        );

    \I__2608\ : LocalMux
    port map (
            O => \N__17834\,
            I => \b2v_inst.g3_0\
        );

    \I__2607\ : InMux
    port map (
            O => \N__17831\,
            I => \N__17828\
        );

    \I__2606\ : LocalMux
    port map (
            O => \N__17828\,
            I => \b2v_inst.g0_4_5\
        );

    \I__2605\ : IoInMux
    port map (
            O => \N__17825\,
            I => \N__17822\
        );

    \I__2604\ : LocalMux
    port map (
            O => \N__17822\,
            I => \N__17818\
        );

    \I__2603\ : InMux
    port map (
            O => \N__17821\,
            I => \N__17815\
        );

    \I__2602\ : Span4Mux_s3_h
    port map (
            O => \N__17818\,
            I => \N__17812\
        );

    \I__2601\ : LocalMux
    port map (
            O => \N__17815\,
            I => \N__17809\
        );

    \I__2600\ : Span4Mux_h
    port map (
            O => \N__17812\,
            I => \N__17806\
        );

    \I__2599\ : Span4Mux_h
    port map (
            O => \N__17809\,
            I => \N__17803\
        );

    \I__2598\ : Span4Mux_v
    port map (
            O => \N__17806\,
            I => \N__17798\
        );

    \I__2597\ : Span4Mux_h
    port map (
            O => \N__17803\,
            I => \N__17798\
        );

    \I__2596\ : Odrv4
    port map (
            O => \N__17798\,
            I => leds_c_10
        );

    \I__2595\ : IoInMux
    port map (
            O => \N__17795\,
            I => \N__17792\
        );

    \I__2594\ : LocalMux
    port map (
            O => \N__17792\,
            I => \N__17789\
        );

    \I__2593\ : IoSpan4Mux
    port map (
            O => \N__17789\,
            I => \N__17786\
        );

    \I__2592\ : Span4Mux_s2_v
    port map (
            O => \N__17786\,
            I => \N__17783\
        );

    \I__2591\ : Span4Mux_h
    port map (
            O => \N__17783\,
            I => \N__17779\
        );

    \I__2590\ : InMux
    port map (
            O => \N__17782\,
            I => \N__17776\
        );

    \I__2589\ : Span4Mux_v
    port map (
            O => \N__17779\,
            I => \N__17773\
        );

    \I__2588\ : LocalMux
    port map (
            O => \N__17776\,
            I => \N__17770\
        );

    \I__2587\ : Odrv4
    port map (
            O => \N__17773\,
            I => leds_c_11
        );

    \I__2586\ : Odrv12
    port map (
            O => \N__17770\,
            I => leds_c_11
        );

    \I__2585\ : InMux
    port map (
            O => \N__17765\,
            I => \N__17761\
        );

    \I__2584\ : IoInMux
    port map (
            O => \N__17764\,
            I => \N__17758\
        );

    \I__2583\ : LocalMux
    port map (
            O => \N__17761\,
            I => \N__17755\
        );

    \I__2582\ : LocalMux
    port map (
            O => \N__17758\,
            I => \N__17752\
        );

    \I__2581\ : Span4Mux_h
    port map (
            O => \N__17755\,
            I => \N__17749\
        );

    \I__2580\ : Span12Mux_s7_h
    port map (
            O => \N__17752\,
            I => \N__17746\
        );

    \I__2579\ : Span4Mux_v
    port map (
            O => \N__17749\,
            I => \N__17743\
        );

    \I__2578\ : Odrv12
    port map (
            O => \N__17746\,
            I => leds_c_7
        );

    \I__2577\ : Odrv4
    port map (
            O => \N__17743\,
            I => leds_c_7
        );

    \I__2576\ : InMux
    port map (
            O => \N__17738\,
            I => \N__17735\
        );

    \I__2575\ : LocalMux
    port map (
            O => \N__17735\,
            I => \b2v_inst.G_40_i_3\
        );

    \I__2574\ : InMux
    port map (
            O => \N__17732\,
            I => \N__17724\
        );

    \I__2573\ : InMux
    port map (
            O => \N__17731\,
            I => \N__17715\
        );

    \I__2572\ : InMux
    port map (
            O => \N__17730\,
            I => \N__17715\
        );

    \I__2571\ : InMux
    port map (
            O => \N__17729\,
            I => \N__17715\
        );

    \I__2570\ : InMux
    port map (
            O => \N__17728\,
            I => \N__17710\
        );

    \I__2569\ : CascadeMux
    port map (
            O => \N__17727\,
            I => \N__17706\
        );

    \I__2568\ : LocalMux
    port map (
            O => \N__17724\,
            I => \N__17702\
        );

    \I__2567\ : CascadeMux
    port map (
            O => \N__17723\,
            I => \N__17699\
        );

    \I__2566\ : InMux
    port map (
            O => \N__17722\,
            I => \N__17696\
        );

    \I__2565\ : LocalMux
    port map (
            O => \N__17715\,
            I => \N__17692\
        );

    \I__2564\ : InMux
    port map (
            O => \N__17714\,
            I => \N__17689\
        );

    \I__2563\ : InMux
    port map (
            O => \N__17713\,
            I => \N__17686\
        );

    \I__2562\ : LocalMux
    port map (
            O => \N__17710\,
            I => \N__17682\
        );

    \I__2561\ : InMux
    port map (
            O => \N__17709\,
            I => \N__17677\
        );

    \I__2560\ : InMux
    port map (
            O => \N__17706\,
            I => \N__17677\
        );

    \I__2559\ : InMux
    port map (
            O => \N__17705\,
            I => \N__17674\
        );

    \I__2558\ : Span4Mux_v
    port map (
            O => \N__17702\,
            I => \N__17671\
        );

    \I__2557\ : InMux
    port map (
            O => \N__17699\,
            I => \N__17668\
        );

    \I__2556\ : LocalMux
    port map (
            O => \N__17696\,
            I => \N__17665\
        );

    \I__2555\ : InMux
    port map (
            O => \N__17695\,
            I => \N__17662\
        );

    \I__2554\ : Span4Mux_h
    port map (
            O => \N__17692\,
            I => \N__17659\
        );

    \I__2553\ : LocalMux
    port map (
            O => \N__17689\,
            I => \N__17656\
        );

    \I__2552\ : LocalMux
    port map (
            O => \N__17686\,
            I => \N__17653\
        );

    \I__2551\ : InMux
    port map (
            O => \N__17685\,
            I => \N__17650\
        );

    \I__2550\ : Span4Mux_h
    port map (
            O => \N__17682\,
            I => \N__17645\
        );

    \I__2549\ : LocalMux
    port map (
            O => \N__17677\,
            I => \N__17645\
        );

    \I__2548\ : LocalMux
    port map (
            O => \N__17674\,
            I => \N__17636\
        );

    \I__2547\ : Span4Mux_h
    port map (
            O => \N__17671\,
            I => \N__17636\
        );

    \I__2546\ : LocalMux
    port map (
            O => \N__17668\,
            I => \N__17636\
        );

    \I__2545\ : Span4Mux_v
    port map (
            O => \N__17665\,
            I => \N__17636\
        );

    \I__2544\ : LocalMux
    port map (
            O => \N__17662\,
            I => \SYNTHESIZED_WIRE_4_19\
        );

    \I__2543\ : Odrv4
    port map (
            O => \N__17659\,
            I => \SYNTHESIZED_WIRE_4_19\
        );

    \I__2542\ : Odrv4
    port map (
            O => \N__17656\,
            I => \SYNTHESIZED_WIRE_4_19\
        );

    \I__2541\ : Odrv4
    port map (
            O => \N__17653\,
            I => \SYNTHESIZED_WIRE_4_19\
        );

    \I__2540\ : LocalMux
    port map (
            O => \N__17650\,
            I => \SYNTHESIZED_WIRE_4_19\
        );

    \I__2539\ : Odrv4
    port map (
            O => \N__17645\,
            I => \SYNTHESIZED_WIRE_4_19\
        );

    \I__2538\ : Odrv4
    port map (
            O => \N__17636\,
            I => \SYNTHESIZED_WIRE_4_19\
        );

    \I__2537\ : InMux
    port map (
            O => \N__17621\,
            I => \N__17617\
        );

    \I__2536\ : InMux
    port map (
            O => \N__17620\,
            I => \N__17614\
        );

    \I__2535\ : LocalMux
    port map (
            O => \N__17617\,
            I => \N__17605\
        );

    \I__2534\ : LocalMux
    port map (
            O => \N__17614\,
            I => \N__17605\
        );

    \I__2533\ : InMux
    port map (
            O => \N__17613\,
            I => \N__17602\
        );

    \I__2532\ : InMux
    port map (
            O => \N__17612\,
            I => \N__17599\
        );

    \I__2531\ : InMux
    port map (
            O => \N__17611\,
            I => \N__17595\
        );

    \I__2530\ : InMux
    port map (
            O => \N__17610\,
            I => \N__17589\
        );

    \I__2529\ : Span4Mux_v
    port map (
            O => \N__17605\,
            I => \N__17584\
        );

    \I__2528\ : LocalMux
    port map (
            O => \N__17602\,
            I => \N__17584\
        );

    \I__2527\ : LocalMux
    port map (
            O => \N__17599\,
            I => \N__17581\
        );

    \I__2526\ : InMux
    port map (
            O => \N__17598\,
            I => \N__17578\
        );

    \I__2525\ : LocalMux
    port map (
            O => \N__17595\,
            I => \N__17575\
        );

    \I__2524\ : InMux
    port map (
            O => \N__17594\,
            I => \N__17572\
        );

    \I__2523\ : InMux
    port map (
            O => \N__17593\,
            I => \N__17569\
        );

    \I__2522\ : InMux
    port map (
            O => \N__17592\,
            I => \N__17566\
        );

    \I__2521\ : LocalMux
    port map (
            O => \N__17589\,
            I => \N__17562\
        );

    \I__2520\ : Span4Mux_h
    port map (
            O => \N__17584\,
            I => \N__17559\
        );

    \I__2519\ : Span4Mux_h
    port map (
            O => \N__17581\,
            I => \N__17552\
        );

    \I__2518\ : LocalMux
    port map (
            O => \N__17578\,
            I => \N__17552\
        );

    \I__2517\ : Span4Mux_v
    port map (
            O => \N__17575\,
            I => \N__17552\
        );

    \I__2516\ : LocalMux
    port map (
            O => \N__17572\,
            I => \N__17549\
        );

    \I__2515\ : LocalMux
    port map (
            O => \N__17569\,
            I => \N__17544\
        );

    \I__2514\ : LocalMux
    port map (
            O => \N__17566\,
            I => \N__17544\
        );

    \I__2513\ : InMux
    port map (
            O => \N__17565\,
            I => \N__17541\
        );

    \I__2512\ : Span4Mux_h
    port map (
            O => \N__17562\,
            I => \N__17538\
        );

    \I__2511\ : Odrv4
    port map (
            O => \N__17559\,
            I => \SYNTHESIZED_WIRE_4_16\
        );

    \I__2510\ : Odrv4
    port map (
            O => \N__17552\,
            I => \SYNTHESIZED_WIRE_4_16\
        );

    \I__2509\ : Odrv4
    port map (
            O => \N__17549\,
            I => \SYNTHESIZED_WIRE_4_16\
        );

    \I__2508\ : Odrv4
    port map (
            O => \N__17544\,
            I => \SYNTHESIZED_WIRE_4_16\
        );

    \I__2507\ : LocalMux
    port map (
            O => \N__17541\,
            I => \SYNTHESIZED_WIRE_4_16\
        );

    \I__2506\ : Odrv4
    port map (
            O => \N__17538\,
            I => \SYNTHESIZED_WIRE_4_16\
        );

    \I__2505\ : InMux
    port map (
            O => \N__17525\,
            I => \N__17521\
        );

    \I__2504\ : InMux
    port map (
            O => \N__17524\,
            I => \N__17518\
        );

    \I__2503\ : LocalMux
    port map (
            O => \N__17521\,
            I => \b2v_inst.N_5\
        );

    \I__2502\ : LocalMux
    port map (
            O => \N__17518\,
            I => \b2v_inst.N_5\
        );

    \I__2501\ : CascadeMux
    port map (
            O => \N__17513\,
            I => \b2v_inst.N_430_i_1_cascade_\
        );

    \I__2500\ : InMux
    port map (
            O => \N__17510\,
            I => \N__17506\
        );

    \I__2499\ : InMux
    port map (
            O => \N__17509\,
            I => \N__17503\
        );

    \I__2498\ : LocalMux
    port map (
            O => \N__17506\,
            I => \N__17497\
        );

    \I__2497\ : LocalMux
    port map (
            O => \N__17503\,
            I => \N__17494\
        );

    \I__2496\ : InMux
    port map (
            O => \N__17502\,
            I => \N__17491\
        );

    \I__2495\ : InMux
    port map (
            O => \N__17501\,
            I => \N__17485\
        );

    \I__2494\ : InMux
    port map (
            O => \N__17500\,
            I => \N__17485\
        );

    \I__2493\ : Span4Mux_v
    port map (
            O => \N__17497\,
            I => \N__17476\
        );

    \I__2492\ : Span4Mux_v
    port map (
            O => \N__17494\,
            I => \N__17476\
        );

    \I__2491\ : LocalMux
    port map (
            O => \N__17491\,
            I => \N__17476\
        );

    \I__2490\ : InMux
    port map (
            O => \N__17490\,
            I => \N__17473\
        );

    \I__2489\ : LocalMux
    port map (
            O => \N__17485\,
            I => \N__17470\
        );

    \I__2488\ : InMux
    port map (
            O => \N__17484\,
            I => \N__17467\
        );

    \I__2487\ : InMux
    port map (
            O => \N__17483\,
            I => \N__17464\
        );

    \I__2486\ : Span4Mux_h
    port map (
            O => \N__17476\,
            I => \N__17461\
        );

    \I__2485\ : LocalMux
    port map (
            O => \N__17473\,
            I => \N__17456\
        );

    \I__2484\ : Span4Mux_v
    port map (
            O => \N__17470\,
            I => \N__17456\
        );

    \I__2483\ : LocalMux
    port map (
            O => \N__17467\,
            I => \SYNTHESIZED_WIRE_4_18\
        );

    \I__2482\ : LocalMux
    port map (
            O => \N__17464\,
            I => \SYNTHESIZED_WIRE_4_18\
        );

    \I__2481\ : Odrv4
    port map (
            O => \N__17461\,
            I => \SYNTHESIZED_WIRE_4_18\
        );

    \I__2480\ : Odrv4
    port map (
            O => \N__17456\,
            I => \SYNTHESIZED_WIRE_4_18\
        );

    \I__2479\ : InMux
    port map (
            O => \N__17447\,
            I => \N__17441\
        );

    \I__2478\ : InMux
    port map (
            O => \N__17446\,
            I => \N__17438\
        );

    \I__2477\ : InMux
    port map (
            O => \N__17445\,
            I => \N__17433\
        );

    \I__2476\ : InMux
    port map (
            O => \N__17444\,
            I => \N__17428\
        );

    \I__2475\ : LocalMux
    port map (
            O => \N__17441\,
            I => \N__17423\
        );

    \I__2474\ : LocalMux
    port map (
            O => \N__17438\,
            I => \N__17423\
        );

    \I__2473\ : InMux
    port map (
            O => \N__17437\,
            I => \N__17420\
        );

    \I__2472\ : InMux
    port map (
            O => \N__17436\,
            I => \N__17417\
        );

    \I__2471\ : LocalMux
    port map (
            O => \N__17433\,
            I => \N__17414\
        );

    \I__2470\ : InMux
    port map (
            O => \N__17432\,
            I => \N__17411\
        );

    \I__2469\ : InMux
    port map (
            O => \N__17431\,
            I => \N__17408\
        );

    \I__2468\ : LocalMux
    port map (
            O => \N__17428\,
            I => \N__17405\
        );

    \I__2467\ : Span4Mux_v
    port map (
            O => \N__17423\,
            I => \N__17402\
        );

    \I__2466\ : LocalMux
    port map (
            O => \N__17420\,
            I => \N__17397\
        );

    \I__2465\ : LocalMux
    port map (
            O => \N__17417\,
            I => \N__17397\
        );

    \I__2464\ : Span4Mux_h
    port map (
            O => \N__17414\,
            I => \N__17394\
        );

    \I__2463\ : LocalMux
    port map (
            O => \N__17411\,
            I => \SYNTHESIZED_WIRE_4_17\
        );

    \I__2462\ : LocalMux
    port map (
            O => \N__17408\,
            I => \SYNTHESIZED_WIRE_4_17\
        );

    \I__2461\ : Odrv4
    port map (
            O => \N__17405\,
            I => \SYNTHESIZED_WIRE_4_17\
        );

    \I__2460\ : Odrv4
    port map (
            O => \N__17402\,
            I => \SYNTHESIZED_WIRE_4_17\
        );

    \I__2459\ : Odrv4
    port map (
            O => \N__17397\,
            I => \SYNTHESIZED_WIRE_4_17\
        );

    \I__2458\ : Odrv4
    port map (
            O => \N__17394\,
            I => \SYNTHESIZED_WIRE_4_17\
        );

    \I__2457\ : CascadeMux
    port map (
            O => \N__17381\,
            I => \N__17377\
        );

    \I__2456\ : CascadeMux
    port map (
            O => \N__17380\,
            I => \N__17373\
        );

    \I__2455\ : InMux
    port map (
            O => \N__17377\,
            I => \N__17370\
        );

    \I__2454\ : InMux
    port map (
            O => \N__17376\,
            I => \N__17365\
        );

    \I__2453\ : InMux
    port map (
            O => \N__17373\,
            I => \N__17365\
        );

    \I__2452\ : LocalMux
    port map (
            O => \N__17370\,
            I => \b2v_inst.g1Z0Z_0\
        );

    \I__2451\ : LocalMux
    port map (
            O => \N__17365\,
            I => \b2v_inst.g1Z0Z_0\
        );

    \I__2450\ : InMux
    port map (
            O => \N__17360\,
            I => \N__17357\
        );

    \I__2449\ : LocalMux
    port map (
            O => \N__17357\,
            I => \b2v_inst.pix_count_anterior5\
        );

    \I__2448\ : CascadeMux
    port map (
            O => \N__17354\,
            I => \b2v_inst.state_ns_0_i_o2_6_23_cascade_\
        );

    \I__2447\ : InMux
    port map (
            O => \N__17351\,
            I => \N__17348\
        );

    \I__2446\ : LocalMux
    port map (
            O => \N__17348\,
            I => \b2v_inst.state_ns_0_i_o2_7_23\
        );

    \I__2445\ : CascadeMux
    port map (
            O => \N__17345\,
            I => \b2v_inst.g0_6_cascade_\
        );

    \I__2444\ : InMux
    port map (
            O => \N__17342\,
            I => \N__17339\
        );

    \I__2443\ : LocalMux
    port map (
            O => \N__17339\,
            I => \b2v_inst.o2\
        );

    \I__2442\ : CascadeMux
    port map (
            O => \N__17336\,
            I => \b2v_inst.G_40_i_6_cascade_\
        );

    \I__2441\ : InMux
    port map (
            O => \N__17333\,
            I => \N__17330\
        );

    \I__2440\ : LocalMux
    port map (
            O => \N__17330\,
            I => \b2v_inst.state_ns_i_0_a2_11_a2_0_3_3\
        );

    \I__2439\ : InMux
    port map (
            O => \N__17327\,
            I => \N__17324\
        );

    \I__2438\ : LocalMux
    port map (
            O => \N__17324\,
            I => \b2v_inst.N_618_5\
        );

    \I__2437\ : InMux
    port map (
            O => \N__17321\,
            I => \N__17318\
        );

    \I__2436\ : LocalMux
    port map (
            O => \N__17318\,
            I => \N__17315\
        );

    \I__2435\ : Span4Mux_h
    port map (
            O => \N__17315\,
            I => \N__17311\
        );

    \I__2434\ : InMux
    port map (
            O => \N__17314\,
            I => \N__17308\
        );

    \I__2433\ : Odrv4
    port map (
            O => \N__17311\,
            I => \b2v_inst1.N_49\
        );

    \I__2432\ : LocalMux
    port map (
            O => \N__17308\,
            I => \b2v_inst1.N_49\
        );

    \I__2431\ : InMux
    port map (
            O => \N__17303\,
            I => \N__17294\
        );

    \I__2430\ : InMux
    port map (
            O => \N__17302\,
            I => \N__17294\
        );

    \I__2429\ : InMux
    port map (
            O => \N__17301\,
            I => \N__17291\
        );

    \I__2428\ : InMux
    port map (
            O => \N__17300\,
            I => \N__17286\
        );

    \I__2427\ : InMux
    port map (
            O => \N__17299\,
            I => \N__17282\
        );

    \I__2426\ : LocalMux
    port map (
            O => \N__17294\,
            I => \N__17279\
        );

    \I__2425\ : LocalMux
    port map (
            O => \N__17291\,
            I => \N__17276\
        );

    \I__2424\ : InMux
    port map (
            O => \N__17290\,
            I => \N__17273\
        );

    \I__2423\ : InMux
    port map (
            O => \N__17289\,
            I => \N__17270\
        );

    \I__2422\ : LocalMux
    port map (
            O => \N__17286\,
            I => \N__17267\
        );

    \I__2421\ : InMux
    port map (
            O => \N__17285\,
            I => \N__17264\
        );

    \I__2420\ : LocalMux
    port map (
            O => \N__17282\,
            I => \N__17261\
        );

    \I__2419\ : Span4Mux_v
    port map (
            O => \N__17279\,
            I => \N__17254\
        );

    \I__2418\ : Span4Mux_v
    port map (
            O => \N__17276\,
            I => \N__17254\
        );

    \I__2417\ : LocalMux
    port map (
            O => \N__17273\,
            I => \N__17254\
        );

    \I__2416\ : LocalMux
    port map (
            O => \N__17270\,
            I => \N__17247\
        );

    \I__2415\ : Span4Mux_h
    port map (
            O => \N__17267\,
            I => \N__17247\
        );

    \I__2414\ : LocalMux
    port map (
            O => \N__17264\,
            I => \N__17247\
        );

    \I__2413\ : Span4Mux_v
    port map (
            O => \N__17261\,
            I => \N__17242\
        );

    \I__2412\ : Span4Mux_h
    port map (
            O => \N__17254\,
            I => \N__17242\
        );

    \I__2411\ : Span4Mux_v
    port map (
            O => \N__17247\,
            I => \N__17239\
        );

    \I__2410\ : Odrv4
    port map (
            O => \N__17242\,
            I => \b2v_inst1.r_RX_Byte_1_sqmuxa\
        );

    \I__2409\ : Odrv4
    port map (
            O => \N__17239\,
            I => \b2v_inst1.r_RX_Byte_1_sqmuxa\
        );

    \I__2408\ : InMux
    port map (
            O => \N__17234\,
            I => \N__17231\
        );

    \I__2407\ : LocalMux
    port map (
            O => \N__17231\,
            I => \b2v_inst.N_618_3\
        );

    \I__2406\ : InMux
    port map (
            O => \N__17228\,
            I => \N__17225\
        );

    \I__2405\ : LocalMux
    port map (
            O => \N__17225\,
            I => \b2v_inst.state_ns_i_0_a2_11_o2_4_0_3_3\
        );

    \I__2404\ : CascadeMux
    port map (
            O => \N__17222\,
            I => \N__17218\
        );

    \I__2403\ : InMux
    port map (
            O => \N__17221\,
            I => \N__17214\
        );

    \I__2402\ : InMux
    port map (
            O => \N__17218\,
            I => \N__17209\
        );

    \I__2401\ : InMux
    port map (
            O => \N__17217\,
            I => \N__17209\
        );

    \I__2400\ : LocalMux
    port map (
            O => \N__17214\,
            I => \N__17206\
        );

    \I__2399\ : LocalMux
    port map (
            O => \N__17209\,
            I => \b2v_inst.un4_pix_count_intlto19_0_0\
        );

    \I__2398\ : Odrv12
    port map (
            O => \N__17206\,
            I => \b2v_inst.un4_pix_count_intlto19_0_0\
        );

    \I__2397\ : CascadeMux
    port map (
            O => \N__17201\,
            I => \N__17198\
        );

    \I__2396\ : InMux
    port map (
            O => \N__17198\,
            I => \N__17195\
        );

    \I__2395\ : LocalMux
    port map (
            O => \N__17195\,
            I => \b2v_inst.G_40_i_2\
        );

    \I__2394\ : IoInMux
    port map (
            O => \N__17192\,
            I => \N__17189\
        );

    \I__2393\ : LocalMux
    port map (
            O => \N__17189\,
            I => \N__17186\
        );

    \I__2392\ : IoSpan4Mux
    port map (
            O => \N__17186\,
            I => \N__17182\
        );

    \I__2391\ : InMux
    port map (
            O => \N__17185\,
            I => \N__17179\
        );

    \I__2390\ : Span4Mux_s3_v
    port map (
            O => \N__17182\,
            I => \N__17176\
        );

    \I__2389\ : LocalMux
    port map (
            O => \N__17179\,
            I => \N__17173\
        );

    \I__2388\ : Span4Mux_v
    port map (
            O => \N__17176\,
            I => \N__17170\
        );

    \I__2387\ : Span4Mux_v
    port map (
            O => \N__17173\,
            I => \N__17167\
        );

    \I__2386\ : Span4Mux_v
    port map (
            O => \N__17170\,
            I => \N__17164\
        );

    \I__2385\ : Span4Mux_h
    port map (
            O => \N__17167\,
            I => \N__17161\
        );

    \I__2384\ : Odrv4
    port map (
            O => \N__17164\,
            I => leds_c_4
        );

    \I__2383\ : Odrv4
    port map (
            O => \N__17161\,
            I => leds_c_4
        );

    \I__2382\ : IoInMux
    port map (
            O => \N__17156\,
            I => \N__17153\
        );

    \I__2381\ : LocalMux
    port map (
            O => \N__17153\,
            I => \N__17150\
        );

    \I__2380\ : Span4Mux_s3_v
    port map (
            O => \N__17150\,
            I => \N__17146\
        );

    \I__2379\ : InMux
    port map (
            O => \N__17149\,
            I => \N__17143\
        );

    \I__2378\ : Sp12to4
    port map (
            O => \N__17146\,
            I => \N__17140\
        );

    \I__2377\ : LocalMux
    port map (
            O => \N__17143\,
            I => \N__17137\
        );

    \I__2376\ : Span12Mux_s11_h
    port map (
            O => \N__17140\,
            I => \N__17134\
        );

    \I__2375\ : Span4Mux_h
    port map (
            O => \N__17137\,
            I => \N__17131\
        );

    \I__2374\ : Span12Mux_v
    port map (
            O => \N__17134\,
            I => \N__17128\
        );

    \I__2373\ : Span4Mux_v
    port map (
            O => \N__17131\,
            I => \N__17125\
        );

    \I__2372\ : Odrv12
    port map (
            O => \N__17128\,
            I => leds_c_5
        );

    \I__2371\ : Odrv4
    port map (
            O => \N__17125\,
            I => leds_c_5
        );

    \I__2370\ : InMux
    port map (
            O => \N__17120\,
            I => \N__17117\
        );

    \I__2369\ : LocalMux
    port map (
            O => \N__17117\,
            I => \b2v_inst.dir_mem_115lt6_0\
        );

    \I__2368\ : CascadeMux
    port map (
            O => \N__17114\,
            I => \b2v_inst.g0_1_0_cascade_\
        );

    \I__2367\ : InMux
    port map (
            O => \N__17111\,
            I => \N__17108\
        );

    \I__2366\ : LocalMux
    port map (
            O => \N__17108\,
            I => \N__17105\
        );

    \I__2365\ : Span4Mux_h
    port map (
            O => \N__17105\,
            I => \N__17101\
        );

    \I__2364\ : InMux
    port map (
            O => \N__17104\,
            I => \N__17098\
        );

    \I__2363\ : Span4Mux_h
    port map (
            O => \N__17101\,
            I => \N__17095\
        );

    \I__2362\ : LocalMux
    port map (
            O => \N__17098\,
            I => \N__17092\
        );

    \I__2361\ : Odrv4
    port map (
            O => \N__17095\,
            I => \b2v_inst.un7_pix_count_int_0_N_2_THRU_CO\
        );

    \I__2360\ : Odrv12
    port map (
            O => \N__17092\,
            I => \b2v_inst.un7_pix_count_int_0_N_2_THRU_CO\
        );

    \I__2359\ : InMux
    port map (
            O => \N__17087\,
            I => \b2v_inst.un8_dir_mem_2_cry_4\
        );

    \I__2358\ : InMux
    port map (
            O => \N__17084\,
            I => \b2v_inst.un8_dir_mem_2_cry_5\
        );

    \I__2357\ : InMux
    port map (
            O => \N__17081\,
            I => \b2v_inst.un8_dir_mem_2_cry_6\
        );

    \I__2356\ : InMux
    port map (
            O => \N__17078\,
            I => \b2v_inst.un8_dir_mem_2_cry_7\
        );

    \I__2355\ : InMux
    port map (
            O => \N__17075\,
            I => \bfn_9_6_0_\
        );

    \I__2354\ : InMux
    port map (
            O => \N__17072\,
            I => \b2v_inst.un8_dir_mem_2_cry_9\
        );

    \I__2353\ : InMux
    port map (
            O => \N__17069\,
            I => \N__17066\
        );

    \I__2352\ : LocalMux
    port map (
            O => \N__17066\,
            I => \b2v_inst.dir_mem_215lt6_0\
        );

    \I__2351\ : CascadeMux
    port map (
            O => \N__17063\,
            I => \b2v_inst1.N_36_cascade_\
        );

    \I__2350\ : CascadeMux
    port map (
            O => \N__17060\,
            I => \N__17057\
        );

    \I__2349\ : InMux
    port map (
            O => \N__17057\,
            I => \N__17049\
        );

    \I__2348\ : InMux
    port map (
            O => \N__17056\,
            I => \N__17049\
        );

    \I__2347\ : CascadeMux
    port map (
            O => \N__17055\,
            I => \N__17043\
        );

    \I__2346\ : InMux
    port map (
            O => \N__17054\,
            I => \N__17038\
        );

    \I__2345\ : LocalMux
    port map (
            O => \N__17049\,
            I => \N__17035\
        );

    \I__2344\ : InMux
    port map (
            O => \N__17048\,
            I => \N__17028\
        );

    \I__2343\ : InMux
    port map (
            O => \N__17047\,
            I => \N__17028\
        );

    \I__2342\ : InMux
    port map (
            O => \N__17046\,
            I => \N__17028\
        );

    \I__2341\ : InMux
    port map (
            O => \N__17043\,
            I => \N__17021\
        );

    \I__2340\ : InMux
    port map (
            O => \N__17042\,
            I => \N__17021\
        );

    \I__2339\ : InMux
    port map (
            O => \N__17041\,
            I => \N__17021\
        );

    \I__2338\ : LocalMux
    port map (
            O => \N__17038\,
            I => \b2v_inst1.r_Bit_IndexZ0Z_1\
        );

    \I__2337\ : Odrv12
    port map (
            O => \N__17035\,
            I => \b2v_inst1.r_Bit_IndexZ0Z_1\
        );

    \I__2336\ : LocalMux
    port map (
            O => \N__17028\,
            I => \b2v_inst1.r_Bit_IndexZ0Z_1\
        );

    \I__2335\ : LocalMux
    port map (
            O => \N__17021\,
            I => \b2v_inst1.r_Bit_IndexZ0Z_1\
        );

    \I__2334\ : InMux
    port map (
            O => \N__17012\,
            I => \N__17006\
        );

    \I__2333\ : InMux
    port map (
            O => \N__17011\,
            I => \N__17001\
        );

    \I__2332\ : InMux
    port map (
            O => \N__17010\,
            I => \N__17001\
        );

    \I__2331\ : InMux
    port map (
            O => \N__17009\,
            I => \N__16992\
        );

    \I__2330\ : LocalMux
    port map (
            O => \N__17006\,
            I => \N__16987\
        );

    \I__2329\ : LocalMux
    port map (
            O => \N__17001\,
            I => \N__16987\
        );

    \I__2328\ : InMux
    port map (
            O => \N__17000\,
            I => \N__16982\
        );

    \I__2327\ : InMux
    port map (
            O => \N__16999\,
            I => \N__16982\
        );

    \I__2326\ : InMux
    port map (
            O => \N__16998\,
            I => \N__16973\
        );

    \I__2325\ : InMux
    port map (
            O => \N__16997\,
            I => \N__16973\
        );

    \I__2324\ : InMux
    port map (
            O => \N__16996\,
            I => \N__16973\
        );

    \I__2323\ : InMux
    port map (
            O => \N__16995\,
            I => \N__16973\
        );

    \I__2322\ : LocalMux
    port map (
            O => \N__16992\,
            I => \b2v_inst1.r_Bit_IndexZ0Z_0\
        );

    \I__2321\ : Odrv4
    port map (
            O => \N__16987\,
            I => \b2v_inst1.r_Bit_IndexZ0Z_0\
        );

    \I__2320\ : LocalMux
    port map (
            O => \N__16982\,
            I => \b2v_inst1.r_Bit_IndexZ0Z_0\
        );

    \I__2319\ : LocalMux
    port map (
            O => \N__16973\,
            I => \b2v_inst1.r_Bit_IndexZ0Z_0\
        );

    \I__2318\ : InMux
    port map (
            O => \N__16964\,
            I => \N__16961\
        );

    \I__2317\ : LocalMux
    port map (
            O => \N__16961\,
            I => \b2v_inst1.N_50\
        );

    \I__2316\ : CascadeMux
    port map (
            O => \N__16958\,
            I => \N__16955\
        );

    \I__2315\ : InMux
    port map (
            O => \N__16955\,
            I => \N__16952\
        );

    \I__2314\ : LocalMux
    port map (
            O => \N__16952\,
            I => \b2v_inst1.r_RX_Bytece_0_5\
        );

    \I__2313\ : InMux
    port map (
            O => \N__16949\,
            I => \N__16946\
        );

    \I__2312\ : LocalMux
    port map (
            O => \N__16946\,
            I => \N__16943\
        );

    \I__2311\ : Odrv12
    port map (
            O => \N__16943\,
            I => \N_460_i\
        );

    \I__2310\ : InMux
    port map (
            O => \N__16940\,
            I => \N__16937\
        );

    \I__2309\ : LocalMux
    port map (
            O => \N__16937\,
            I => \N__16934\
        );

    \I__2308\ : Span4Mux_v
    port map (
            O => \N__16934\,
            I => \N__16931\
        );

    \I__2307\ : Odrv4
    port map (
            O => \N__16931\,
            I => \N_459_i\
        );

    \I__2306\ : InMux
    port map (
            O => \N__16928\,
            I => \b2v_inst.un8_dir_mem_2_cry_1\
        );

    \I__2305\ : InMux
    port map (
            O => \N__16925\,
            I => \b2v_inst.un8_dir_mem_2_cry_2\
        );

    \I__2304\ : InMux
    port map (
            O => \N__16922\,
            I => \b2v_inst.un8_dir_mem_2_cry_3\
        );

    \I__2303\ : InMux
    port map (
            O => \N__16919\,
            I => \N__16916\
        );

    \I__2302\ : LocalMux
    port map (
            O => \N__16916\,
            I => \b2v_inst1.r_RX_Bytece_0_6\
        );

    \I__2301\ : CascadeMux
    port map (
            O => \N__16913\,
            I => \N__16910\
        );

    \I__2300\ : InMux
    port map (
            O => \N__16910\,
            I => \N__16907\
        );

    \I__2299\ : LocalMux
    port map (
            O => \N__16907\,
            I => \N__16898\
        );

    \I__2298\ : InMux
    port map (
            O => \N__16906\,
            I => \N__16893\
        );

    \I__2297\ : InMux
    port map (
            O => \N__16905\,
            I => \N__16893\
        );

    \I__2296\ : InMux
    port map (
            O => \N__16904\,
            I => \N__16890\
        );

    \I__2295\ : InMux
    port map (
            O => \N__16903\,
            I => \N__16887\
        );

    \I__2294\ : InMux
    port map (
            O => \N__16902\,
            I => \N__16882\
        );

    \I__2293\ : InMux
    port map (
            O => \N__16901\,
            I => \N__16882\
        );

    \I__2292\ : Span4Mux_h
    port map (
            O => \N__16898\,
            I => \N__16879\
        );

    \I__2291\ : LocalMux
    port map (
            O => \N__16893\,
            I => \N__16876\
        );

    \I__2290\ : LocalMux
    port map (
            O => \N__16890\,
            I => \b2v_inst1.r_Clk_CountZ0Z_2\
        );

    \I__2289\ : LocalMux
    port map (
            O => \N__16887\,
            I => \b2v_inst1.r_Clk_CountZ0Z_2\
        );

    \I__2288\ : LocalMux
    port map (
            O => \N__16882\,
            I => \b2v_inst1.r_Clk_CountZ0Z_2\
        );

    \I__2287\ : Odrv4
    port map (
            O => \N__16879\,
            I => \b2v_inst1.r_Clk_CountZ0Z_2\
        );

    \I__2286\ : Odrv4
    port map (
            O => \N__16876\,
            I => \b2v_inst1.r_Clk_CountZ0Z_2\
        );

    \I__2285\ : CascadeMux
    port map (
            O => \N__16865\,
            I => \b2v_inst1.m16_0_o2_cascade_\
        );

    \I__2284\ : InMux
    port map (
            O => \N__16862\,
            I => \N__16859\
        );

    \I__2283\ : LocalMux
    port map (
            O => \N__16859\,
            I => \N__16856\
        );

    \I__2282\ : Odrv4
    port map (
            O => \N__16856\,
            I => \b2v_inst.g0_1_0_0\
        );

    \I__2281\ : InMux
    port map (
            O => \N__16853\,
            I => \N__16849\
        );

    \I__2280\ : CascadeMux
    port map (
            O => \N__16852\,
            I => \N__16844\
        );

    \I__2279\ : LocalMux
    port map (
            O => \N__16849\,
            I => \N__16839\
        );

    \I__2278\ : InMux
    port map (
            O => \N__16848\,
            I => \N__16836\
        );

    \I__2277\ : InMux
    port map (
            O => \N__16847\,
            I => \N__16833\
        );

    \I__2276\ : InMux
    port map (
            O => \N__16844\,
            I => \N__16828\
        );

    \I__2275\ : InMux
    port map (
            O => \N__16843\,
            I => \N__16828\
        );

    \I__2274\ : InMux
    port map (
            O => \N__16842\,
            I => \N__16825\
        );

    \I__2273\ : Span4Mux_v
    port map (
            O => \N__16839\,
            I => \N__16816\
        );

    \I__2272\ : LocalMux
    port map (
            O => \N__16836\,
            I => \N__16816\
        );

    \I__2271\ : LocalMux
    port map (
            O => \N__16833\,
            I => \N__16813\
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__16828\,
            I => \N__16810\
        );

    \I__2269\ : LocalMux
    port map (
            O => \N__16825\,
            I => \N__16807\
        );

    \I__2268\ : InMux
    port map (
            O => \N__16824\,
            I => \N__16800\
        );

    \I__2267\ : InMux
    port map (
            O => \N__16823\,
            I => \N__16800\
        );

    \I__2266\ : InMux
    port map (
            O => \N__16822\,
            I => \N__16800\
        );

    \I__2265\ : InMux
    port map (
            O => \N__16821\,
            I => \N__16797\
        );

    \I__2264\ : Span4Mux_h
    port map (
            O => \N__16816\,
            I => \N__16794\
        );

    \I__2263\ : Span4Mux_v
    port map (
            O => \N__16813\,
            I => \N__16789\
        );

    \I__2262\ : Span4Mux_v
    port map (
            O => \N__16810\,
            I => \N__16789\
        );

    \I__2261\ : Span4Mux_h
    port map (
            O => \N__16807\,
            I => \N__16784\
        );

    \I__2260\ : LocalMux
    port map (
            O => \N__16800\,
            I => \N__16784\
        );

    \I__2259\ : LocalMux
    port map (
            O => \N__16797\,
            I => \SYNTHESIZED_WIRE_4_7\
        );

    \I__2258\ : Odrv4
    port map (
            O => \N__16794\,
            I => \SYNTHESIZED_WIRE_4_7\
        );

    \I__2257\ : Odrv4
    port map (
            O => \N__16789\,
            I => \SYNTHESIZED_WIRE_4_7\
        );

    \I__2256\ : Odrv4
    port map (
            O => \N__16784\,
            I => \SYNTHESIZED_WIRE_4_7\
        );

    \I__2255\ : CascadeMux
    port map (
            O => \N__16775\,
            I => \N__16772\
        );

    \I__2254\ : InMux
    port map (
            O => \N__16772\,
            I => \N__16769\
        );

    \I__2253\ : LocalMux
    port map (
            O => \N__16769\,
            I => \N__16766\
        );

    \I__2252\ : Span4Mux_v
    port map (
            O => \N__16766\,
            I => \N__16763\
        );

    \I__2251\ : Span4Mux_h
    port map (
            O => \N__16763\,
            I => \N__16760\
        );

    \I__2250\ : Odrv4
    port map (
            O => \N__16760\,
            I => \b2v_inst.un4_pix_count_intlto6_d_1_2\
        );

    \I__2249\ : InMux
    port map (
            O => \N__16757\,
            I => \N__16753\
        );

    \I__2248\ : InMux
    port map (
            O => \N__16756\,
            I => \N__16749\
        );

    \I__2247\ : LocalMux
    port map (
            O => \N__16753\,
            I => \N__16741\
        );

    \I__2246\ : InMux
    port map (
            O => \N__16752\,
            I => \N__16738\
        );

    \I__2245\ : LocalMux
    port map (
            O => \N__16749\,
            I => \N__16735\
        );

    \I__2244\ : InMux
    port map (
            O => \N__16748\,
            I => \N__16728\
        );

    \I__2243\ : InMux
    port map (
            O => \N__16747\,
            I => \N__16728\
        );

    \I__2242\ : InMux
    port map (
            O => \N__16746\,
            I => \N__16728\
        );

    \I__2241\ : InMux
    port map (
            O => \N__16745\,
            I => \N__16724\
        );

    \I__2240\ : InMux
    port map (
            O => \N__16744\,
            I => \N__16721\
        );

    \I__2239\ : Span4Mux_v
    port map (
            O => \N__16741\,
            I => \N__16716\
        );

    \I__2238\ : LocalMux
    port map (
            O => \N__16738\,
            I => \N__16716\
        );

    \I__2237\ : Span4Mux_v
    port map (
            O => \N__16735\,
            I => \N__16711\
        );

    \I__2236\ : LocalMux
    port map (
            O => \N__16728\,
            I => \N__16711\
        );

    \I__2235\ : InMux
    port map (
            O => \N__16727\,
            I => \N__16708\
        );

    \I__2234\ : LocalMux
    port map (
            O => \N__16724\,
            I => \N__16703\
        );

    \I__2233\ : LocalMux
    port map (
            O => \N__16721\,
            I => \N__16703\
        );

    \I__2232\ : Span4Mux_v
    port map (
            O => \N__16716\,
            I => \N__16700\
        );

    \I__2231\ : Span4Mux_h
    port map (
            O => \N__16711\,
            I => \N__16697\
        );

    \I__2230\ : LocalMux
    port map (
            O => \N__16708\,
            I => \SYNTHESIZED_WIRE_4_4\
        );

    \I__2229\ : Odrv4
    port map (
            O => \N__16703\,
            I => \SYNTHESIZED_WIRE_4_4\
        );

    \I__2228\ : Odrv4
    port map (
            O => \N__16700\,
            I => \SYNTHESIZED_WIRE_4_4\
        );

    \I__2227\ : Odrv4
    port map (
            O => \N__16697\,
            I => \SYNTHESIZED_WIRE_4_4\
        );

    \I__2226\ : InMux
    port map (
            O => \N__16688\,
            I => \N__16685\
        );

    \I__2225\ : LocalMux
    port map (
            O => \N__16685\,
            I => \b2v_inst.g1_0_0\
        );

    \I__2224\ : InMux
    port map (
            O => \N__16682\,
            I => \N__16679\
        );

    \I__2223\ : LocalMux
    port map (
            O => \N__16679\,
            I => \b2v_inst.g1_0_0Z0Z_2\
        );

    \I__2222\ : CascadeMux
    port map (
            O => \N__16676\,
            I => \N__16673\
        );

    \I__2221\ : InMux
    port map (
            O => \N__16673\,
            I => \N__16670\
        );

    \I__2220\ : LocalMux
    port map (
            O => \N__16670\,
            I => \b2v_inst.g1_0_a4Z0Z_0\
        );

    \I__2219\ : InMux
    port map (
            O => \N__16667\,
            I => \N__16664\
        );

    \I__2218\ : LocalMux
    port map (
            O => \N__16664\,
            I => \N__16661\
        );

    \I__2217\ : Sp12to4
    port map (
            O => \N__16661\,
            I => \N__16658\
        );

    \I__2216\ : Span12Mux_v
    port map (
            O => \N__16658\,
            I => \N__16655\
        );

    \I__2215\ : Span12Mux_h
    port map (
            O => \N__16655\,
            I => \N__16652\
        );

    \I__2214\ : Odrv12
    port map (
            O => \N__16652\,
            I => swit_c_9
        );

    \I__2213\ : InMux
    port map (
            O => \N__16649\,
            I => \N__16646\
        );

    \I__2212\ : LocalMux
    port map (
            O => \N__16646\,
            I => \b2v_inst.addr_ram_energia_m0_9\
        );

    \I__2211\ : CascadeMux
    port map (
            O => \N__16643\,
            I => \b2v_inst1.N_38_cascade_\
        );

    \I__2210\ : InMux
    port map (
            O => \N__16640\,
            I => \N__16633\
        );

    \I__2209\ : InMux
    port map (
            O => \N__16639\,
            I => \N__16633\
        );

    \I__2208\ : InMux
    port map (
            O => \N__16638\,
            I => \N__16624\
        );

    \I__2207\ : LocalMux
    port map (
            O => \N__16633\,
            I => \N__16621\
        );

    \I__2206\ : InMux
    port map (
            O => \N__16632\,
            I => \N__16618\
        );

    \I__2205\ : InMux
    port map (
            O => \N__16631\,
            I => \N__16615\
        );

    \I__2204\ : InMux
    port map (
            O => \N__16630\,
            I => \N__16612\
        );

    \I__2203\ : InMux
    port map (
            O => \N__16629\,
            I => \N__16609\
        );

    \I__2202\ : InMux
    port map (
            O => \N__16628\,
            I => \N__16606\
        );

    \I__2201\ : InMux
    port map (
            O => \N__16627\,
            I => \N__16603\
        );

    \I__2200\ : LocalMux
    port map (
            O => \N__16624\,
            I => \N__16596\
        );

    \I__2199\ : Span4Mux_v
    port map (
            O => \N__16621\,
            I => \N__16596\
        );

    \I__2198\ : LocalMux
    port map (
            O => \N__16618\,
            I => \N__16596\
        );

    \I__2197\ : LocalMux
    port map (
            O => \N__16615\,
            I => \b2v_inst1.r_Bit_IndexZ0Z_2\
        );

    \I__2196\ : LocalMux
    port map (
            O => \N__16612\,
            I => \b2v_inst1.r_Bit_IndexZ0Z_2\
        );

    \I__2195\ : LocalMux
    port map (
            O => \N__16609\,
            I => \b2v_inst1.r_Bit_IndexZ0Z_2\
        );

    \I__2194\ : LocalMux
    port map (
            O => \N__16606\,
            I => \b2v_inst1.r_Bit_IndexZ0Z_2\
        );

    \I__2193\ : LocalMux
    port map (
            O => \N__16603\,
            I => \b2v_inst1.r_Bit_IndexZ0Z_2\
        );

    \I__2192\ : Odrv4
    port map (
            O => \N__16596\,
            I => \b2v_inst1.r_Bit_IndexZ0Z_2\
        );

    \I__2191\ : InMux
    port map (
            O => \N__16583\,
            I => \N__16580\
        );

    \I__2190\ : LocalMux
    port map (
            O => \N__16580\,
            I => \b2v_inst1.N_44\
        );

    \I__2189\ : CascadeMux
    port map (
            O => \N__16577\,
            I => \b2v_inst1.N_96_cascade_\
        );

    \I__2188\ : InMux
    port map (
            O => \N__16574\,
            I => \N__16571\
        );

    \I__2187\ : LocalMux
    port map (
            O => \N__16571\,
            I => \b2v_inst.g0_0_i_a4Z0Z_0\
        );

    \I__2186\ : InMux
    port map (
            O => \N__16568\,
            I => \N__16565\
        );

    \I__2185\ : LocalMux
    port map (
            O => \N__16565\,
            I => \N__16562\
        );

    \I__2184\ : Odrv4
    port map (
            O => \N__16562\,
            I => \b2v_inst.g0_0_iZ0Z_2\
        );

    \I__2183\ : CascadeMux
    port map (
            O => \N__16559\,
            I => \N__16556\
        );

    \I__2182\ : InMux
    port map (
            O => \N__16556\,
            I => \N__16553\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__16553\,
            I => \N__16550\
        );

    \I__2180\ : Span12Mux_h
    port map (
            O => \N__16550\,
            I => \N__16547\
        );

    \I__2179\ : Odrv12
    port map (
            O => \N__16547\,
            I => \b2v_inst.g2Z0Z_1\
        );

    \I__2178\ : CascadeMux
    port map (
            O => \N__16544\,
            I => \b2v_inst1.N_58_i_cascade_\
        );

    \I__2177\ : InMux
    port map (
            O => \N__16541\,
            I => \N__16537\
        );

    \I__2176\ : InMux
    port map (
            O => \N__16540\,
            I => \N__16533\
        );

    \I__2175\ : LocalMux
    port map (
            O => \N__16537\,
            I => \N__16530\
        );

    \I__2174\ : InMux
    port map (
            O => \N__16536\,
            I => \N__16527\
        );

    \I__2173\ : LocalMux
    port map (
            O => \N__16533\,
            I => \N__16524\
        );

    \I__2172\ : Odrv12
    port map (
            O => \N__16530\,
            I => \b2v_inst1.un22_r_clk_count_ac0_3\
        );

    \I__2171\ : LocalMux
    port map (
            O => \N__16527\,
            I => \b2v_inst1.un22_r_clk_count_ac0_3\
        );

    \I__2170\ : Odrv4
    port map (
            O => \N__16524\,
            I => \b2v_inst1.un22_r_clk_count_ac0_3\
        );

    \I__2169\ : InMux
    port map (
            O => \N__16517\,
            I => \b2v_inst.un3_dir_mem_cry_5\
        );

    \I__2168\ : InMux
    port map (
            O => \N__16514\,
            I => \b2v_inst.un3_dir_mem_cry_6\
        );

    \I__2167\ : InMux
    port map (
            O => \N__16511\,
            I => \bfn_8_10_0_\
        );

    \I__2166\ : InMux
    port map (
            O => \N__16508\,
            I => \b2v_inst.un3_dir_mem_cry_8\
        );

    \I__2165\ : InMux
    port map (
            O => \N__16505\,
            I => \b2v_inst.un3_dir_mem_cry_9\
        );

    \I__2164\ : InMux
    port map (
            O => \N__16502\,
            I => \N__16495\
        );

    \I__2163\ : InMux
    port map (
            O => \N__16501\,
            I => \N__16491\
        );

    \I__2162\ : InMux
    port map (
            O => \N__16500\,
            I => \N__16488\
        );

    \I__2161\ : InMux
    port map (
            O => \N__16499\,
            I => \N__16485\
        );

    \I__2160\ : InMux
    port map (
            O => \N__16498\,
            I => \N__16482\
        );

    \I__2159\ : LocalMux
    port map (
            O => \N__16495\,
            I => \N__16479\
        );

    \I__2158\ : InMux
    port map (
            O => \N__16494\,
            I => \N__16476\
        );

    \I__2157\ : LocalMux
    port map (
            O => \N__16491\,
            I => \N__16470\
        );

    \I__2156\ : LocalMux
    port map (
            O => \N__16488\,
            I => \N__16465\
        );

    \I__2155\ : LocalMux
    port map (
            O => \N__16485\,
            I => \N__16465\
        );

    \I__2154\ : LocalMux
    port map (
            O => \N__16482\,
            I => \N__16458\
        );

    \I__2153\ : Span4Mux_h
    port map (
            O => \N__16479\,
            I => \N__16458\
        );

    \I__2152\ : LocalMux
    port map (
            O => \N__16476\,
            I => \N__16458\
        );

    \I__2151\ : InMux
    port map (
            O => \N__16475\,
            I => \N__16453\
        );

    \I__2150\ : InMux
    port map (
            O => \N__16474\,
            I => \N__16453\
        );

    \I__2149\ : InMux
    port map (
            O => \N__16473\,
            I => \N__16450\
        );

    \I__2148\ : Span4Mux_v
    port map (
            O => \N__16470\,
            I => \N__16447\
        );

    \I__2147\ : Span4Mux_v
    port map (
            O => \N__16465\,
            I => \N__16442\
        );

    \I__2146\ : Span4Mux_v
    port map (
            O => \N__16458\,
            I => \N__16442\
        );

    \I__2145\ : LocalMux
    port map (
            O => \N__16453\,
            I => \N__16439\
        );

    \I__2144\ : LocalMux
    port map (
            O => \N__16450\,
            I => \SYNTHESIZED_WIRE_4_13\
        );

    \I__2143\ : Odrv4
    port map (
            O => \N__16447\,
            I => \SYNTHESIZED_WIRE_4_13\
        );

    \I__2142\ : Odrv4
    port map (
            O => \N__16442\,
            I => \SYNTHESIZED_WIRE_4_13\
        );

    \I__2141\ : Odrv4
    port map (
            O => \N__16439\,
            I => \SYNTHESIZED_WIRE_4_13\
        );

    \I__2140\ : InMux
    port map (
            O => \N__16430\,
            I => \N__16426\
        );

    \I__2139\ : InMux
    port map (
            O => \N__16429\,
            I => \N__16420\
        );

    \I__2138\ : LocalMux
    port map (
            O => \N__16426\,
            I => \N__16417\
        );

    \I__2137\ : InMux
    port map (
            O => \N__16425\,
            I => \N__16414\
        );

    \I__2136\ : InMux
    port map (
            O => \N__16424\,
            I => \N__16411\
        );

    \I__2135\ : InMux
    port map (
            O => \N__16423\,
            I => \N__16404\
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__16420\,
            I => \N__16399\
        );

    \I__2133\ : Span4Mux_h
    port map (
            O => \N__16417\,
            I => \N__16399\
        );

    \I__2132\ : LocalMux
    port map (
            O => \N__16414\,
            I => \N__16394\
        );

    \I__2131\ : LocalMux
    port map (
            O => \N__16411\,
            I => \N__16394\
        );

    \I__2130\ : InMux
    port map (
            O => \N__16410\,
            I => \N__16387\
        );

    \I__2129\ : InMux
    port map (
            O => \N__16409\,
            I => \N__16387\
        );

    \I__2128\ : InMux
    port map (
            O => \N__16408\,
            I => \N__16387\
        );

    \I__2127\ : InMux
    port map (
            O => \N__16407\,
            I => \N__16384\
        );

    \I__2126\ : LocalMux
    port map (
            O => \N__16404\,
            I => \N__16379\
        );

    \I__2125\ : Span4Mux_v
    port map (
            O => \N__16399\,
            I => \N__16379\
        );

    \I__2124\ : Span4Mux_h
    port map (
            O => \N__16394\,
            I => \N__16376\
        );

    \I__2123\ : LocalMux
    port map (
            O => \N__16387\,
            I => \N__16373\
        );

    \I__2122\ : LocalMux
    port map (
            O => \N__16384\,
            I => \SYNTHESIZED_WIRE_4_15\
        );

    \I__2121\ : Odrv4
    port map (
            O => \N__16379\,
            I => \SYNTHESIZED_WIRE_4_15\
        );

    \I__2120\ : Odrv4
    port map (
            O => \N__16376\,
            I => \SYNTHESIZED_WIRE_4_15\
        );

    \I__2119\ : Odrv4
    port map (
            O => \N__16373\,
            I => \SYNTHESIZED_WIRE_4_15\
        );

    \I__2118\ : CascadeMux
    port map (
            O => \N__16364\,
            I => \N__16359\
        );

    \I__2117\ : InMux
    port map (
            O => \N__16363\,
            I => \N__16355\
        );

    \I__2116\ : InMux
    port map (
            O => \N__16362\,
            I => \N__16351\
        );

    \I__2115\ : InMux
    port map (
            O => \N__16359\,
            I => \N__16347\
        );

    \I__2114\ : InMux
    port map (
            O => \N__16358\,
            I => \N__16344\
        );

    \I__2113\ : LocalMux
    port map (
            O => \N__16355\,
            I => \N__16341\
        );

    \I__2112\ : InMux
    port map (
            O => \N__16354\,
            I => \N__16335\
        );

    \I__2111\ : LocalMux
    port map (
            O => \N__16351\,
            I => \N__16332\
        );

    \I__2110\ : InMux
    port map (
            O => \N__16350\,
            I => \N__16329\
        );

    \I__2109\ : LocalMux
    port map (
            O => \N__16347\,
            I => \N__16326\
        );

    \I__2108\ : LocalMux
    port map (
            O => \N__16344\,
            I => \N__16323\
        );

    \I__2107\ : Span4Mux_h
    port map (
            O => \N__16341\,
            I => \N__16320\
        );

    \I__2106\ : InMux
    port map (
            O => \N__16340\,
            I => \N__16313\
        );

    \I__2105\ : InMux
    port map (
            O => \N__16339\,
            I => \N__16313\
        );

    \I__2104\ : InMux
    port map (
            O => \N__16338\,
            I => \N__16313\
        );

    \I__2103\ : LocalMux
    port map (
            O => \N__16335\,
            I => \N__16306\
        );

    \I__2102\ : Span4Mux_v
    port map (
            O => \N__16332\,
            I => \N__16306\
        );

    \I__2101\ : LocalMux
    port map (
            O => \N__16329\,
            I => \N__16306\
        );

    \I__2100\ : Span4Mux_h
    port map (
            O => \N__16326\,
            I => \N__16301\
        );

    \I__2099\ : Span4Mux_h
    port map (
            O => \N__16323\,
            I => \N__16301\
        );

    \I__2098\ : Span4Mux_v
    port map (
            O => \N__16320\,
            I => \N__16296\
        );

    \I__2097\ : LocalMux
    port map (
            O => \N__16313\,
            I => \N__16296\
        );

    \I__2096\ : Odrv4
    port map (
            O => \N__16306\,
            I => \SYNTHESIZED_WIRE_4_14\
        );

    \I__2095\ : Odrv4
    port map (
            O => \N__16301\,
            I => \SYNTHESIZED_WIRE_4_14\
        );

    \I__2094\ : Odrv4
    port map (
            O => \N__16296\,
            I => \SYNTHESIZED_WIRE_4_14\
        );

    \I__2093\ : InMux
    port map (
            O => \N__16289\,
            I => \N__16286\
        );

    \I__2092\ : LocalMux
    port map (
            O => \N__16286\,
            I => \b2v_inst.state_RNO_25Z0Z_29\
        );

    \I__2091\ : InMux
    port map (
            O => \N__16283\,
            I => \N__16280\
        );

    \I__2090\ : LocalMux
    port map (
            O => \N__16280\,
            I => \N__16277\
        );

    \I__2089\ : Odrv4
    port map (
            O => \N__16277\,
            I => \b2v_inst.g2_1_0\
        );

    \I__2088\ : CascadeMux
    port map (
            O => \N__16274\,
            I => \b2v_inst.m29_2_cascade_\
        );

    \I__2087\ : InMux
    port map (
            O => \N__16271\,
            I => \N__16268\
        );

    \I__2086\ : LocalMux
    port map (
            O => \N__16268\,
            I => \N__16263\
        );

    \I__2085\ : InMux
    port map (
            O => \N__16267\,
            I => \N__16260\
        );

    \I__2084\ : InMux
    port map (
            O => \N__16266\,
            I => \N__16257\
        );

    \I__2083\ : Odrv12
    port map (
            O => \N__16263\,
            I => \b2v_inst.un4_pix_count_intlto10_1_d_0\
        );

    \I__2082\ : LocalMux
    port map (
            O => \N__16260\,
            I => \b2v_inst.un4_pix_count_intlto10_1_d_0\
        );

    \I__2081\ : LocalMux
    port map (
            O => \N__16257\,
            I => \b2v_inst.un4_pix_count_intlto10_1_d_0\
        );

    \I__2080\ : CascadeMux
    port map (
            O => \N__16250\,
            I => \N__16247\
        );

    \I__2079\ : InMux
    port map (
            O => \N__16247\,
            I => \N__16242\
        );

    \I__2078\ : InMux
    port map (
            O => \N__16246\,
            I => \N__16239\
        );

    \I__2077\ : InMux
    port map (
            O => \N__16245\,
            I => \N__16236\
        );

    \I__2076\ : LocalMux
    port map (
            O => \N__16242\,
            I => \N__16233\
        );

    \I__2075\ : LocalMux
    port map (
            O => \N__16239\,
            I => \N__16230\
        );

    \I__2074\ : LocalMux
    port map (
            O => \N__16236\,
            I => \N__16225\
        );

    \I__2073\ : Span4Mux_v
    port map (
            O => \N__16233\,
            I => \N__16225\
        );

    \I__2072\ : Odrv12
    port map (
            O => \N__16230\,
            I => \b2v_inst.indice_RNIJFHBZ0Z_0\
        );

    \I__2071\ : Odrv4
    port map (
            O => \N__16225\,
            I => \b2v_inst.indice_RNIJFHBZ0Z_0\
        );

    \I__2070\ : InMux
    port map (
            O => \N__16220\,
            I => \N__16217\
        );

    \I__2069\ : LocalMux
    port map (
            O => \N__16217\,
            I => \N__16212\
        );

    \I__2068\ : InMux
    port map (
            O => \N__16216\,
            I => \N__16209\
        );

    \I__2067\ : InMux
    port map (
            O => \N__16215\,
            I => \N__16206\
        );

    \I__2066\ : Span4Mux_h
    port map (
            O => \N__16212\,
            I => \N__16203\
        );

    \I__2065\ : LocalMux
    port map (
            O => \N__16209\,
            I => \N__16200\
        );

    \I__2064\ : LocalMux
    port map (
            O => \N__16206\,
            I => \b2v_inst.un1_indice_cry_5_c_RNI69OGZ0\
        );

    \I__2063\ : Odrv4
    port map (
            O => \N__16203\,
            I => \b2v_inst.un1_indice_cry_5_c_RNI69OGZ0\
        );

    \I__2062\ : Odrv4
    port map (
            O => \N__16200\,
            I => \b2v_inst.un1_indice_cry_5_c_RNI69OGZ0\
        );

    \I__2061\ : CascadeMux
    port map (
            O => \N__16193\,
            I => \N__16190\
        );

    \I__2060\ : InMux
    port map (
            O => \N__16190\,
            I => \N__16187\
        );

    \I__2059\ : LocalMux
    port map (
            O => \N__16187\,
            I => \N__16184\
        );

    \I__2058\ : Span4Mux_v
    port map (
            O => \N__16184\,
            I => \N__16181\
        );

    \I__2057\ : Span4Mux_h
    port map (
            O => \N__16181\,
            I => \N__16178\
        );

    \I__2056\ : Odrv4
    port map (
            O => \N__16178\,
            I => \b2v_inst.dir_mem_3_RNO_0Z0Z_6\
        );

    \I__2055\ : InMux
    port map (
            O => \N__16175\,
            I => \b2v_inst.un3_dir_mem_cry_1\
        );

    \I__2054\ : InMux
    port map (
            O => \N__16172\,
            I => \b2v_inst.un3_dir_mem_cry_2\
        );

    \I__2053\ : InMux
    port map (
            O => \N__16169\,
            I => \b2v_inst.un3_dir_mem_cry_3\
        );

    \I__2052\ : InMux
    port map (
            O => \N__16166\,
            I => \b2v_inst.un3_dir_mem_cry_4\
        );

    \I__2051\ : InMux
    port map (
            O => \N__16163\,
            I => \b2v_inst.un2_dir_mem_1_cry_8\
        );

    \I__2050\ : CascadeMux
    port map (
            O => \N__16160\,
            I => \N__16156\
        );

    \I__2049\ : InMux
    port map (
            O => \N__16159\,
            I => \N__16151\
        );

    \I__2048\ : InMux
    port map (
            O => \N__16156\,
            I => \N__16151\
        );

    \I__2047\ : LocalMux
    port map (
            O => \N__16151\,
            I => \N__16147\
        );

    \I__2046\ : InMux
    port map (
            O => \N__16150\,
            I => \N__16144\
        );

    \I__2045\ : Odrv4
    port map (
            O => \N__16147\,
            I => \b2v_inst.un1_indice_cry_10_THRU_CO\
        );

    \I__2044\ : LocalMux
    port map (
            O => \N__16144\,
            I => \b2v_inst.un1_indice_cry_10_THRU_CO\
        );

    \I__2043\ : CascadeMux
    port map (
            O => \N__16139\,
            I => \N__16136\
        );

    \I__2042\ : InMux
    port map (
            O => \N__16136\,
            I => \N__16133\
        );

    \I__2041\ : LocalMux
    port map (
            O => \N__16133\,
            I => \N__16130\
        );

    \I__2040\ : Span4Mux_h
    port map (
            O => \N__16130\,
            I => \N__16127\
        );

    \I__2039\ : Span4Mux_h
    port map (
            O => \N__16127\,
            I => \N__16124\
        );

    \I__2038\ : Odrv4
    port map (
            O => \N__16124\,
            I => \b2v_inst.dir_mem_3_RNO_0Z0Z_10\
        );

    \I__2037\ : CascadeMux
    port map (
            O => \N__16121\,
            I => \N__16118\
        );

    \I__2036\ : InMux
    port map (
            O => \N__16118\,
            I => \N__16115\
        );

    \I__2035\ : LocalMux
    port map (
            O => \N__16115\,
            I => \N__16112\
        );

    \I__2034\ : Span4Mux_v
    port map (
            O => \N__16112\,
            I => \N__16109\
        );

    \I__2033\ : Odrv4
    port map (
            O => \N__16109\,
            I => \b2v_inst.dir_mem_3_RNO_0Z0Z_7\
        );

    \I__2032\ : CascadeMux
    port map (
            O => \N__16106\,
            I => \N__16103\
        );

    \I__2031\ : InMux
    port map (
            O => \N__16103\,
            I => \N__16100\
        );

    \I__2030\ : LocalMux
    port map (
            O => \N__16100\,
            I => \N__16097\
        );

    \I__2029\ : Span4Mux_v
    port map (
            O => \N__16097\,
            I => \N__16094\
        );

    \I__2028\ : Odrv4
    port map (
            O => \N__16094\,
            I => \b2v_inst.dir_mem_3_RNO_0Z0Z_8\
        );

    \I__2027\ : CascadeMux
    port map (
            O => \N__16091\,
            I => \N__16088\
        );

    \I__2026\ : InMux
    port map (
            O => \N__16088\,
            I => \N__16085\
        );

    \I__2025\ : LocalMux
    port map (
            O => \N__16085\,
            I => \N__16082\
        );

    \I__2024\ : Span4Mux_h
    port map (
            O => \N__16082\,
            I => \N__16079\
        );

    \I__2023\ : Odrv4
    port map (
            O => \N__16079\,
            I => \b2v_inst.dir_mem_3_RNO_0Z0Z_9\
        );

    \I__2022\ : InMux
    port map (
            O => \N__16076\,
            I => \N__16073\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__16073\,
            I => \N__16068\
        );

    \I__2020\ : InMux
    port map (
            O => \N__16072\,
            I => \N__16065\
        );

    \I__2019\ : InMux
    port map (
            O => \N__16071\,
            I => \N__16062\
        );

    \I__2018\ : Span4Mux_h
    port map (
            O => \N__16068\,
            I => \N__16059\
        );

    \I__2017\ : LocalMux
    port map (
            O => \N__16065\,
            I => \N__16056\
        );

    \I__2016\ : LocalMux
    port map (
            O => \N__16062\,
            I => \b2v_inst.un1_indice_cry_2_c_RNI00LGZ0\
        );

    \I__2015\ : Odrv4
    port map (
            O => \N__16059\,
            I => \b2v_inst.un1_indice_cry_2_c_RNI00LGZ0\
        );

    \I__2014\ : Odrv4
    port map (
            O => \N__16056\,
            I => \b2v_inst.un1_indice_cry_2_c_RNI00LGZ0\
        );

    \I__2013\ : InMux
    port map (
            O => \N__16049\,
            I => \b2v_inst.un2_dir_mem_1_cry_3\
        );

    \I__2012\ : InMux
    port map (
            O => \N__16046\,
            I => \b2v_inst.un2_dir_mem_1_cry_4\
        );

    \I__2011\ : InMux
    port map (
            O => \N__16043\,
            I => \b2v_inst.un2_dir_mem_1_cry_5\
        );

    \I__2010\ : InMux
    port map (
            O => \N__16040\,
            I => \b2v_inst.un2_dir_mem_1_cry_6\
        );

    \I__2009\ : InMux
    port map (
            O => \N__16037\,
            I => \bfn_8_6_0_\
        );

    \I__2008\ : CascadeMux
    port map (
            O => \N__16034\,
            I => \N__16031\
        );

    \I__2007\ : InMux
    port map (
            O => \N__16031\,
            I => \N__16028\
        );

    \I__2006\ : LocalMux
    port map (
            O => \N__16028\,
            I => \b2v_inst.N_8\
        );

    \I__2005\ : InMux
    port map (
            O => \N__16025\,
            I => \N__16022\
        );

    \I__2004\ : LocalMux
    port map (
            O => \N__16022\,
            I => \b2v_inst1.N_42\
        );

    \I__2003\ : InMux
    port map (
            O => \N__16019\,
            I => \N__16016\
        );

    \I__2002\ : LocalMux
    port map (
            O => \N__16016\,
            I => \N__16012\
        );

    \I__2001\ : InMux
    port map (
            O => \N__16015\,
            I => \N__16009\
        );

    \I__2000\ : Odrv4
    port map (
            O => \N__16012\,
            I => \b2v_inst1.r_SM_Main_d_4\
        );

    \I__1999\ : LocalMux
    port map (
            O => \N__16009\,
            I => \b2v_inst1.r_SM_Main_d_4\
        );

    \I__1998\ : InMux
    port map (
            O => \N__16004\,
            I => \N__15999\
        );

    \I__1997\ : InMux
    port map (
            O => \N__16003\,
            I => \N__15994\
        );

    \I__1996\ : InMux
    port map (
            O => \N__16002\,
            I => \N__15994\
        );

    \I__1995\ : LocalMux
    port map (
            O => \N__15999\,
            I => \N__15989\
        );

    \I__1994\ : LocalMux
    port map (
            O => \N__15994\,
            I => \N__15989\
        );

    \I__1993\ : Odrv4
    port map (
            O => \N__15989\,
            I => \b2v_inst1.N_47\
        );

    \I__1992\ : CascadeMux
    port map (
            O => \N__15986\,
            I => \b2v_inst1.r_SM_Main_d_4_cascade_\
        );

    \I__1991\ : InMux
    port map (
            O => \N__15983\,
            I => \N__15980\
        );

    \I__1990\ : LocalMux
    port map (
            O => \N__15980\,
            I => \b2v_inst1.N_51\
        );

    \I__1989\ : CascadeMux
    port map (
            O => \N__15977\,
            I => \N__15973\
        );

    \I__1988\ : CascadeMux
    port map (
            O => \N__15976\,
            I => \N__15970\
        );

    \I__1987\ : CascadeBuf
    port map (
            O => \N__15973\,
            I => \N__15967\
        );

    \I__1986\ : CascadeBuf
    port map (
            O => \N__15970\,
            I => \N__15964\
        );

    \I__1985\ : CascadeMux
    port map (
            O => \N__15967\,
            I => \N__15961\
        );

    \I__1984\ : CascadeMux
    port map (
            O => \N__15964\,
            I => \N__15958\
        );

    \I__1983\ : CascadeBuf
    port map (
            O => \N__15961\,
            I => \N__15955\
        );

    \I__1982\ : CascadeBuf
    port map (
            O => \N__15958\,
            I => \N__15952\
        );

    \I__1981\ : CascadeMux
    port map (
            O => \N__15955\,
            I => \N__15949\
        );

    \I__1980\ : CascadeMux
    port map (
            O => \N__15952\,
            I => \N__15946\
        );

    \I__1979\ : CascadeBuf
    port map (
            O => \N__15949\,
            I => \N__15943\
        );

    \I__1978\ : CascadeBuf
    port map (
            O => \N__15946\,
            I => \N__15940\
        );

    \I__1977\ : CascadeMux
    port map (
            O => \N__15943\,
            I => \N__15937\
        );

    \I__1976\ : CascadeMux
    port map (
            O => \N__15940\,
            I => \N__15934\
        );

    \I__1975\ : CascadeBuf
    port map (
            O => \N__15937\,
            I => \N__15931\
        );

    \I__1974\ : CascadeBuf
    port map (
            O => \N__15934\,
            I => \N__15928\
        );

    \I__1973\ : CascadeMux
    port map (
            O => \N__15931\,
            I => \N__15925\
        );

    \I__1972\ : CascadeMux
    port map (
            O => \N__15928\,
            I => \N__15922\
        );

    \I__1971\ : CascadeBuf
    port map (
            O => \N__15925\,
            I => \N__15919\
        );

    \I__1970\ : CascadeBuf
    port map (
            O => \N__15922\,
            I => \N__15916\
        );

    \I__1969\ : CascadeMux
    port map (
            O => \N__15919\,
            I => \N__15913\
        );

    \I__1968\ : CascadeMux
    port map (
            O => \N__15916\,
            I => \N__15910\
        );

    \I__1967\ : CascadeBuf
    port map (
            O => \N__15913\,
            I => \N__15907\
        );

    \I__1966\ : CascadeBuf
    port map (
            O => \N__15910\,
            I => \N__15904\
        );

    \I__1965\ : CascadeMux
    port map (
            O => \N__15907\,
            I => \N__15901\
        );

    \I__1964\ : CascadeMux
    port map (
            O => \N__15904\,
            I => \N__15898\
        );

    \I__1963\ : InMux
    port map (
            O => \N__15901\,
            I => \N__15895\
        );

    \I__1962\ : InMux
    port map (
            O => \N__15898\,
            I => \N__15892\
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__15895\,
            I => \N__15887\
        );

    \I__1960\ : LocalMux
    port map (
            O => \N__15892\,
            I => \N__15887\
        );

    \I__1959\ : Span4Mux_v
    port map (
            O => \N__15887\,
            I => \N__15884\
        );

    \I__1958\ : Span4Mux_h
    port map (
            O => \N__15884\,
            I => \N__15881\
        );

    \I__1957\ : Odrv4
    port map (
            O => \N__15881\,
            I => \SYNTHESIZED_WIRE_12_9\
        );

    \I__1956\ : InMux
    port map (
            O => \N__15878\,
            I => \N__15872\
        );

    \I__1955\ : InMux
    port map (
            O => \N__15877\,
            I => \N__15869\
        );

    \I__1954\ : InMux
    port map (
            O => \N__15876\,
            I => \N__15866\
        );

    \I__1953\ : InMux
    port map (
            O => \N__15875\,
            I => \N__15863\
        );

    \I__1952\ : LocalMux
    port map (
            O => \N__15872\,
            I => \N__15860\
        );

    \I__1951\ : LocalMux
    port map (
            O => \N__15869\,
            I => \N__15854\
        );

    \I__1950\ : LocalMux
    port map (
            O => \N__15866\,
            I => \N__15854\
        );

    \I__1949\ : LocalMux
    port map (
            O => \N__15863\,
            I => \N__15849\
        );

    \I__1948\ : Span4Mux_v
    port map (
            O => \N__15860\,
            I => \N__15849\
        );

    \I__1947\ : CascadeMux
    port map (
            O => \N__15859\,
            I => \N__15845\
        );

    \I__1946\ : Span4Mux_h
    port map (
            O => \N__15854\,
            I => \N__15842\
        );

    \I__1945\ : Sp12to4
    port map (
            O => \N__15849\,
            I => \N__15839\
        );

    \I__1944\ : InMux
    port map (
            O => \N__15848\,
            I => \N__15834\
        );

    \I__1943\ : InMux
    port map (
            O => \N__15845\,
            I => \N__15834\
        );

    \I__1942\ : Odrv4
    port map (
            O => \N__15842\,
            I => \SYNTHESIZED_WIRE_4_6\
        );

    \I__1941\ : Odrv12
    port map (
            O => \N__15839\,
            I => \SYNTHESIZED_WIRE_4_6\
        );

    \I__1940\ : LocalMux
    port map (
            O => \N__15834\,
            I => \SYNTHESIZED_WIRE_4_6\
        );

    \I__1939\ : InMux
    port map (
            O => \N__15827\,
            I => \N__15821\
        );

    \I__1938\ : InMux
    port map (
            O => \N__15826\,
            I => \N__15818\
        );

    \I__1937\ : InMux
    port map (
            O => \N__15825\,
            I => \N__15813\
        );

    \I__1936\ : InMux
    port map (
            O => \N__15824\,
            I => \N__15813\
        );

    \I__1935\ : LocalMux
    port map (
            O => \N__15821\,
            I => \N__15808\
        );

    \I__1934\ : LocalMux
    port map (
            O => \N__15818\,
            I => \N__15808\
        );

    \I__1933\ : LocalMux
    port map (
            O => \N__15813\,
            I => \N__15802\
        );

    \I__1932\ : Span4Mux_h
    port map (
            O => \N__15808\,
            I => \N__15802\
        );

    \I__1931\ : CascadeMux
    port map (
            O => \N__15807\,
            I => \N__15798\
        );

    \I__1930\ : Span4Mux_h
    port map (
            O => \N__15802\,
            I => \N__15795\
        );

    \I__1929\ : InMux
    port map (
            O => \N__15801\,
            I => \N__15792\
        );

    \I__1928\ : InMux
    port map (
            O => \N__15798\,
            I => \N__15789\
        );

    \I__1927\ : Odrv4
    port map (
            O => \N__15795\,
            I => \SYNTHESIZED_WIRE_4_5\
        );

    \I__1926\ : LocalMux
    port map (
            O => \N__15792\,
            I => \SYNTHESIZED_WIRE_4_5\
        );

    \I__1925\ : LocalMux
    port map (
            O => \N__15789\,
            I => \SYNTHESIZED_WIRE_4_5\
        );

    \I__1924\ : CascadeMux
    port map (
            O => \N__15782\,
            I => \b2v_inst.un4_pix_count_intlto6_d_1_0_cascade_\
        );

    \I__1923\ : CascadeMux
    port map (
            O => \N__15779\,
            I => \N__15775\
        );

    \I__1922\ : CascadeMux
    port map (
            O => \N__15778\,
            I => \N__15770\
        );

    \I__1921\ : InMux
    port map (
            O => \N__15775\,
            I => \N__15767\
        );

    \I__1920\ : CascadeMux
    port map (
            O => \N__15774\,
            I => \N__15764\
        );

    \I__1919\ : InMux
    port map (
            O => \N__15773\,
            I => \N__15761\
        );

    \I__1918\ : InMux
    port map (
            O => \N__15770\,
            I => \N__15758\
        );

    \I__1917\ : LocalMux
    port map (
            O => \N__15767\,
            I => \N__15755\
        );

    \I__1916\ : InMux
    port map (
            O => \N__15764\,
            I => \N__15752\
        );

    \I__1915\ : LocalMux
    port map (
            O => \N__15761\,
            I => \N__15749\
        );

    \I__1914\ : LocalMux
    port map (
            O => \N__15758\,
            I => \N__15744\
        );

    \I__1913\ : Span4Mux_v
    port map (
            O => \N__15755\,
            I => \N__15744\
        );

    \I__1912\ : LocalMux
    port map (
            O => \N__15752\,
            I => \N__15741\
        );

    \I__1911\ : Odrv4
    port map (
            O => \N__15749\,
            I => \SYNTHESIZED_WIRE_4_10_rep1\
        );

    \I__1910\ : Odrv4
    port map (
            O => \N__15744\,
            I => \SYNTHESIZED_WIRE_4_10_rep1\
        );

    \I__1909\ : Odrv4
    port map (
            O => \N__15741\,
            I => \SYNTHESIZED_WIRE_4_10_rep1\
        );

    \I__1908\ : CascadeMux
    port map (
            O => \N__15734\,
            I => \N__15731\
        );

    \I__1907\ : InMux
    port map (
            O => \N__15731\,
            I => \N__15726\
        );

    \I__1906\ : InMux
    port map (
            O => \N__15730\,
            I => \N__15722\
        );

    \I__1905\ : InMux
    port map (
            O => \N__15729\,
            I => \N__15719\
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__15726\,
            I => \N__15716\
        );

    \I__1903\ : InMux
    port map (
            O => \N__15725\,
            I => \N__15713\
        );

    \I__1902\ : LocalMux
    port map (
            O => \N__15722\,
            I => \N__15710\
        );

    \I__1901\ : LocalMux
    port map (
            O => \N__15719\,
            I => \N__15707\
        );

    \I__1900\ : Span4Mux_h
    port map (
            O => \N__15716\,
            I => \N__15704\
        );

    \I__1899\ : LocalMux
    port map (
            O => \N__15713\,
            I => \N__15699\
        );

    \I__1898\ : Span4Mux_h
    port map (
            O => \N__15710\,
            I => \N__15699\
        );

    \I__1897\ : Span4Mux_h
    port map (
            O => \N__15707\,
            I => \N__15696\
        );

    \I__1896\ : Span4Mux_h
    port map (
            O => \N__15704\,
            I => \N__15693\
        );

    \I__1895\ : Span4Mux_h
    port map (
            O => \N__15699\,
            I => \N__15690\
        );

    \I__1894\ : Odrv4
    port map (
            O => \N__15696\,
            I => b2v_inst4_pix_count_int_fast_11
        );

    \I__1893\ : Odrv4
    port map (
            O => \N__15693\,
            I => b2v_inst4_pix_count_int_fast_11
        );

    \I__1892\ : Odrv4
    port map (
            O => \N__15690\,
            I => b2v_inst4_pix_count_int_fast_11
        );

    \I__1891\ : InMux
    port map (
            O => \N__15683\,
            I => \N__15678\
        );

    \I__1890\ : CascadeMux
    port map (
            O => \N__15682\,
            I => \N__15675\
        );

    \I__1889\ : InMux
    port map (
            O => \N__15681\,
            I => \N__15671\
        );

    \I__1888\ : LocalMux
    port map (
            O => \N__15678\,
            I => \N__15668\
        );

    \I__1887\ : InMux
    port map (
            O => \N__15675\,
            I => \N__15665\
        );

    \I__1886\ : InMux
    port map (
            O => \N__15674\,
            I => \N__15662\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__15671\,
            I => \N__15659\
        );

    \I__1884\ : Span4Mux_v
    port map (
            O => \N__15668\,
            I => \N__15654\
        );

    \I__1883\ : LocalMux
    port map (
            O => \N__15665\,
            I => \N__15654\
        );

    \I__1882\ : LocalMux
    port map (
            O => \N__15662\,
            I => \N__15649\
        );

    \I__1881\ : Span4Mux_h
    port map (
            O => \N__15659\,
            I => \N__15649\
        );

    \I__1880\ : Span4Mux_h
    port map (
            O => \N__15654\,
            I => \N__15646\
        );

    \I__1879\ : Odrv4
    port map (
            O => \N__15649\,
            I => b2v_inst4_pix_count_int_fast_12
        );

    \I__1878\ : Odrv4
    port map (
            O => \N__15646\,
            I => b2v_inst4_pix_count_int_fast_12
        );

    \I__1877\ : InMux
    port map (
            O => \N__15641\,
            I => \N__15638\
        );

    \I__1876\ : LocalMux
    port map (
            O => \N__15638\,
            I => \N__15635\
        );

    \I__1875\ : Span4Mux_h
    port map (
            O => \N__15635\,
            I => \N__15631\
        );

    \I__1874\ : CascadeMux
    port map (
            O => \N__15634\,
            I => \N__15628\
        );

    \I__1873\ : Span4Mux_h
    port map (
            O => \N__15631\,
            I => \N__15625\
        );

    \I__1872\ : InMux
    port map (
            O => \N__15628\,
            I => \N__15622\
        );

    \I__1871\ : Odrv4
    port map (
            O => \N__15625\,
            I => b2v_inst_un4_pix_count_intlto12_0
        );

    \I__1870\ : LocalMux
    port map (
            O => \N__15622\,
            I => b2v_inst_un4_pix_count_intlto12_0
        );

    \I__1869\ : InMux
    port map (
            O => \N__15617\,
            I => \N__15613\
        );

    \I__1868\ : InMux
    port map (
            O => \N__15616\,
            I => \N__15610\
        );

    \I__1867\ : LocalMux
    port map (
            O => \N__15613\,
            I => \N__15606\
        );

    \I__1866\ : LocalMux
    port map (
            O => \N__15610\,
            I => \N__15603\
        );

    \I__1865\ : InMux
    port map (
            O => \N__15609\,
            I => \N__15600\
        );

    \I__1864\ : Span4Mux_v
    port map (
            O => \N__15606\,
            I => \N__15593\
        );

    \I__1863\ : Span4Mux_h
    port map (
            O => \N__15603\,
            I => \N__15588\
        );

    \I__1862\ : LocalMux
    port map (
            O => \N__15600\,
            I => \N__15588\
        );

    \I__1861\ : InMux
    port map (
            O => \N__15599\,
            I => \N__15585\
        );

    \I__1860\ : InMux
    port map (
            O => \N__15598\,
            I => \N__15582\
        );

    \I__1859\ : InMux
    port map (
            O => \N__15597\,
            I => \N__15577\
        );

    \I__1858\ : InMux
    port map (
            O => \N__15596\,
            I => \N__15577\
        );

    \I__1857\ : Odrv4
    port map (
            O => \N__15593\,
            I => \SYNTHESIZED_WIRE_4_10\
        );

    \I__1856\ : Odrv4
    port map (
            O => \N__15588\,
            I => \SYNTHESIZED_WIRE_4_10\
        );

    \I__1855\ : LocalMux
    port map (
            O => \N__15585\,
            I => \SYNTHESIZED_WIRE_4_10\
        );

    \I__1854\ : LocalMux
    port map (
            O => \N__15582\,
            I => \SYNTHESIZED_WIRE_4_10\
        );

    \I__1853\ : LocalMux
    port map (
            O => \N__15577\,
            I => \SYNTHESIZED_WIRE_4_10\
        );

    \I__1852\ : InMux
    port map (
            O => \N__15566\,
            I => \N__15561\
        );

    \I__1851\ : CascadeMux
    port map (
            O => \N__15565\,
            I => \N__15558\
        );

    \I__1850\ : InMux
    port map (
            O => \N__15564\,
            I => \N__15555\
        );

    \I__1849\ : LocalMux
    port map (
            O => \N__15561\,
            I => \N__15552\
        );

    \I__1848\ : InMux
    port map (
            O => \N__15558\,
            I => \N__15549\
        );

    \I__1847\ : LocalMux
    port map (
            O => \N__15555\,
            I => \N__15543\
        );

    \I__1846\ : Span4Mux_v
    port map (
            O => \N__15552\,
            I => \N__15538\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__15549\,
            I => \N__15538\
        );

    \I__1844\ : InMux
    port map (
            O => \N__15548\,
            I => \N__15533\
        );

    \I__1843\ : InMux
    port map (
            O => \N__15547\,
            I => \N__15533\
        );

    \I__1842\ : CascadeMux
    port map (
            O => \N__15546\,
            I => \N__15530\
        );

    \I__1841\ : Span4Mux_v
    port map (
            O => \N__15543\,
            I => \N__15526\
        );

    \I__1840\ : Span4Mux_h
    port map (
            O => \N__15538\,
            I => \N__15521\
        );

    \I__1839\ : LocalMux
    port map (
            O => \N__15533\,
            I => \N__15521\
        );

    \I__1838\ : InMux
    port map (
            O => \N__15530\,
            I => \N__15518\
        );

    \I__1837\ : InMux
    port map (
            O => \N__15529\,
            I => \N__15515\
        );

    \I__1836\ : Odrv4
    port map (
            O => \N__15526\,
            I => \SYNTHESIZED_WIRE_4_9\
        );

    \I__1835\ : Odrv4
    port map (
            O => \N__15521\,
            I => \SYNTHESIZED_WIRE_4_9\
        );

    \I__1834\ : LocalMux
    port map (
            O => \N__15518\,
            I => \SYNTHESIZED_WIRE_4_9\
        );

    \I__1833\ : LocalMux
    port map (
            O => \N__15515\,
            I => \SYNTHESIZED_WIRE_4_9\
        );

    \I__1832\ : CascadeMux
    port map (
            O => \N__15506\,
            I => \b2v_inst_un4_pix_count_intlto12_0_cascade_\
        );

    \I__1831\ : InMux
    port map (
            O => \N__15503\,
            I => \N__15496\
        );

    \I__1830\ : InMux
    port map (
            O => \N__15502\,
            I => \N__15492\
        );

    \I__1829\ : InMux
    port map (
            O => \N__15501\,
            I => \N__15487\
        );

    \I__1828\ : InMux
    port map (
            O => \N__15500\,
            I => \N__15487\
        );

    \I__1827\ : InMux
    port map (
            O => \N__15499\,
            I => \N__15484\
        );

    \I__1826\ : LocalMux
    port map (
            O => \N__15496\,
            I => \N__15481\
        );

    \I__1825\ : InMux
    port map (
            O => \N__15495\,
            I => \N__15478\
        );

    \I__1824\ : LocalMux
    port map (
            O => \N__15492\,
            I => \N__15474\
        );

    \I__1823\ : LocalMux
    port map (
            O => \N__15487\,
            I => \N__15471\
        );

    \I__1822\ : LocalMux
    port map (
            O => \N__15484\,
            I => \N__15468\
        );

    \I__1821\ : Span4Mux_v
    port map (
            O => \N__15481\,
            I => \N__15463\
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__15478\,
            I => \N__15463\
        );

    \I__1819\ : InMux
    port map (
            O => \N__15477\,
            I => \N__15460\
        );

    \I__1818\ : Span4Mux_v
    port map (
            O => \N__15474\,
            I => \N__15455\
        );

    \I__1817\ : Span4Mux_v
    port map (
            O => \N__15471\,
            I => \N__15455\
        );

    \I__1816\ : Span4Mux_h
    port map (
            O => \N__15468\,
            I => \N__15450\
        );

    \I__1815\ : Span4Mux_h
    port map (
            O => \N__15463\,
            I => \N__15450\
        );

    \I__1814\ : LocalMux
    port map (
            O => \N__15460\,
            I => \SYNTHESIZED_WIRE_4_8\
        );

    \I__1813\ : Odrv4
    port map (
            O => \N__15455\,
            I => \SYNTHESIZED_WIRE_4_8\
        );

    \I__1812\ : Odrv4
    port map (
            O => \N__15450\,
            I => \SYNTHESIZED_WIRE_4_8\
        );

    \I__1811\ : InMux
    port map (
            O => \N__15443\,
            I => \N__15440\
        );

    \I__1810\ : LocalMux
    port map (
            O => \N__15440\,
            I => \N__15437\
        );

    \I__1809\ : Odrv12
    port map (
            O => \N__15437\,
            I => \N_457_i\
        );

    \I__1808\ : InMux
    port map (
            O => \N__15434\,
            I => \N__15431\
        );

    \I__1807\ : LocalMux
    port map (
            O => \N__15431\,
            I => \b2v_inst1.N_48\
        );

    \I__1806\ : CascadeMux
    port map (
            O => \N__15428\,
            I => \b2v_inst1.N_44_cascade_\
        );

    \I__1805\ : InMux
    port map (
            O => \N__15425\,
            I => \N__15422\
        );

    \I__1804\ : LocalMux
    port map (
            O => \N__15422\,
            I => \b2v_inst.un4_pix_count_intlto10_1_0Z0Z_0\
        );

    \I__1803\ : CascadeMux
    port map (
            O => \N__15419\,
            I => \b2v_inst.un4_pix_count_intlt8_cascade_\
        );

    \I__1802\ : InMux
    port map (
            O => \N__15416\,
            I => \N__15413\
        );

    \I__1801\ : LocalMux
    port map (
            O => \N__15413\,
            I => \b2v_inst.un4_pix_count_intlto15_1_aZ0Z0\
        );

    \I__1800\ : InMux
    port map (
            O => \N__15410\,
            I => \N__15406\
        );

    \I__1799\ : InMux
    port map (
            O => \N__15409\,
            I => \N__15403\
        );

    \I__1798\ : LocalMux
    port map (
            O => \N__15406\,
            I => \b2v_inst.un4_pix_count_intlt16\
        );

    \I__1797\ : LocalMux
    port map (
            O => \N__15403\,
            I => \b2v_inst.un4_pix_count_intlt16\
        );

    \I__1796\ : CascadeMux
    port map (
            O => \N__15398\,
            I => \N__15393\
        );

    \I__1795\ : InMux
    port map (
            O => \N__15397\,
            I => \N__15387\
        );

    \I__1794\ : InMux
    port map (
            O => \N__15396\,
            I => \N__15387\
        );

    \I__1793\ : InMux
    port map (
            O => \N__15393\,
            I => \N__15384\
        );

    \I__1792\ : InMux
    port map (
            O => \N__15392\,
            I => \N__15381\
        );

    \I__1791\ : LocalMux
    port map (
            O => \N__15387\,
            I => \N__15378\
        );

    \I__1790\ : LocalMux
    port map (
            O => \N__15384\,
            I => \N__15371\
        );

    \I__1789\ : LocalMux
    port map (
            O => \N__15381\,
            I => \N__15371\
        );

    \I__1788\ : Span4Mux_h
    port map (
            O => \N__15378\,
            I => \N__15368\
        );

    \I__1787\ : InMux
    port map (
            O => \N__15377\,
            I => \N__15363\
        );

    \I__1786\ : InMux
    port map (
            O => \N__15376\,
            I => \N__15363\
        );

    \I__1785\ : Odrv4
    port map (
            O => \N__15371\,
            I => \SYNTHESIZED_WIRE_4_12\
        );

    \I__1784\ : Odrv4
    port map (
            O => \N__15368\,
            I => \SYNTHESIZED_WIRE_4_12\
        );

    \I__1783\ : LocalMux
    port map (
            O => \N__15363\,
            I => \SYNTHESIZED_WIRE_4_12\
        );

    \I__1782\ : CascadeMux
    port map (
            O => \N__15356\,
            I => \N__15353\
        );

    \I__1781\ : InMux
    port map (
            O => \N__15353\,
            I => \N__15349\
        );

    \I__1780\ : InMux
    port map (
            O => \N__15352\,
            I => \N__15346\
        );

    \I__1779\ : LocalMux
    port map (
            O => \N__15349\,
            I => \N__15337\
        );

    \I__1778\ : LocalMux
    port map (
            O => \N__15346\,
            I => \N__15337\
        );

    \I__1777\ : InMux
    port map (
            O => \N__15345\,
            I => \N__15332\
        );

    \I__1776\ : InMux
    port map (
            O => \N__15344\,
            I => \N__15332\
        );

    \I__1775\ : InMux
    port map (
            O => \N__15343\,
            I => \N__15327\
        );

    \I__1774\ : InMux
    port map (
            O => \N__15342\,
            I => \N__15327\
        );

    \I__1773\ : Odrv4
    port map (
            O => \N__15337\,
            I => \SYNTHESIZED_WIRE_4_11\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__15332\,
            I => \SYNTHESIZED_WIRE_4_11\
        );

    \I__1771\ : LocalMux
    port map (
            O => \N__15327\,
            I => \SYNTHESIZED_WIRE_4_11\
        );

    \I__1770\ : InMux
    port map (
            O => \N__15320\,
            I => \N__15316\
        );

    \I__1769\ : InMux
    port map (
            O => \N__15319\,
            I => \N__15313\
        );

    \I__1768\ : LocalMux
    port map (
            O => \N__15316\,
            I => \N__15310\
        );

    \I__1767\ : LocalMux
    port map (
            O => \N__15313\,
            I => \N__15307\
        );

    \I__1766\ : Span4Mux_h
    port map (
            O => \N__15310\,
            I => \N__15302\
        );

    \I__1765\ : Span4Mux_v
    port map (
            O => \N__15307\,
            I => \N__15299\
        );

    \I__1764\ : InMux
    port map (
            O => \N__15306\,
            I => \N__15294\
        );

    \I__1763\ : InMux
    port map (
            O => \N__15305\,
            I => \N__15294\
        );

    \I__1762\ : Odrv4
    port map (
            O => \N__15302\,
            I => \SYNTHESIZED_WIRE_4_9_rep1\
        );

    \I__1761\ : Odrv4
    port map (
            O => \N__15299\,
            I => \SYNTHESIZED_WIRE_4_9_rep1\
        );

    \I__1760\ : LocalMux
    port map (
            O => \N__15294\,
            I => \SYNTHESIZED_WIRE_4_9_rep1\
        );

    \I__1759\ : CascadeMux
    port map (
            O => \N__15287\,
            I => \b2v_inst1.r_RX_Bytece_0_4_cascade_\
        );

    \I__1758\ : CascadeMux
    port map (
            O => \N__15284\,
            I => \b2v_inst.un4_pix_count_intlto10_1_d_0_xZ0Z1_cascade_\
        );

    \I__1757\ : InMux
    port map (
            O => \N__15281\,
            I => \N__15277\
        );

    \I__1756\ : InMux
    port map (
            O => \N__15280\,
            I => \N__15274\
        );

    \I__1755\ : LocalMux
    port map (
            O => \N__15277\,
            I => \N__15266\
        );

    \I__1754\ : LocalMux
    port map (
            O => \N__15274\,
            I => \N__15266\
        );

    \I__1753\ : InMux
    port map (
            O => \N__15273\,
            I => \N__15263\
        );

    \I__1752\ : InMux
    port map (
            O => \N__15272\,
            I => \N__15257\
        );

    \I__1751\ : InMux
    port map (
            O => \N__15271\,
            I => \N__15257\
        );

    \I__1750\ : Span4Mux_h
    port map (
            O => \N__15266\,
            I => \N__15254\
        );

    \I__1749\ : LocalMux
    port map (
            O => \N__15263\,
            I => \N__15251\
        );

    \I__1748\ : InMux
    port map (
            O => \N__15262\,
            I => \N__15248\
        );

    \I__1747\ : LocalMux
    port map (
            O => \N__15257\,
            I => \SYNTHESIZED_WIRE_4_0\
        );

    \I__1746\ : Odrv4
    port map (
            O => \N__15254\,
            I => \SYNTHESIZED_WIRE_4_0\
        );

    \I__1745\ : Odrv4
    port map (
            O => \N__15251\,
            I => \SYNTHESIZED_WIRE_4_0\
        );

    \I__1744\ : LocalMux
    port map (
            O => \N__15248\,
            I => \SYNTHESIZED_WIRE_4_0\
        );

    \I__1743\ : CascadeMux
    port map (
            O => \N__15239\,
            I => \N__15233\
        );

    \I__1742\ : InMux
    port map (
            O => \N__15238\,
            I => \N__15230\
        );

    \I__1741\ : InMux
    port map (
            O => \N__15237\,
            I => \N__15227\
        );

    \I__1740\ : InMux
    port map (
            O => \N__15236\,
            I => \N__15220\
        );

    \I__1739\ : InMux
    port map (
            O => \N__15233\,
            I => \N__15220\
        );

    \I__1738\ : LocalMux
    port map (
            O => \N__15230\,
            I => \N__15215\
        );

    \I__1737\ : LocalMux
    port map (
            O => \N__15227\,
            I => \N__15215\
        );

    \I__1736\ : InMux
    port map (
            O => \N__15226\,
            I => \N__15212\
        );

    \I__1735\ : InMux
    port map (
            O => \N__15225\,
            I => \N__15209\
        );

    \I__1734\ : LocalMux
    port map (
            O => \N__15220\,
            I => \SYNTHESIZED_WIRE_4_3\
        );

    \I__1733\ : Odrv12
    port map (
            O => \N__15215\,
            I => \SYNTHESIZED_WIRE_4_3\
        );

    \I__1732\ : LocalMux
    port map (
            O => \N__15212\,
            I => \SYNTHESIZED_WIRE_4_3\
        );

    \I__1731\ : LocalMux
    port map (
            O => \N__15209\,
            I => \SYNTHESIZED_WIRE_4_3\
        );

    \I__1730\ : CascadeMux
    port map (
            O => \N__15200\,
            I => \N__15194\
        );

    \I__1729\ : CascadeMux
    port map (
            O => \N__15199\,
            I => \N__15190\
        );

    \I__1728\ : CascadeMux
    port map (
            O => \N__15198\,
            I => \N__15187\
        );

    \I__1727\ : InMux
    port map (
            O => \N__15197\,
            I => \N__15184\
        );

    \I__1726\ : InMux
    port map (
            O => \N__15194\,
            I => \N__15181\
        );

    \I__1725\ : InMux
    port map (
            O => \N__15193\,
            I => \N__15178\
        );

    \I__1724\ : InMux
    port map (
            O => \N__15190\,
            I => \N__15175\
        );

    \I__1723\ : InMux
    port map (
            O => \N__15187\,
            I => \N__15172\
        );

    \I__1722\ : LocalMux
    port map (
            O => \N__15184\,
            I => \N__15166\
        );

    \I__1721\ : LocalMux
    port map (
            O => \N__15181\,
            I => \N__15166\
        );

    \I__1720\ : LocalMux
    port map (
            O => \N__15178\,
            I => \N__15163\
        );

    \I__1719\ : LocalMux
    port map (
            O => \N__15175\,
            I => \N__15158\
        );

    \I__1718\ : LocalMux
    port map (
            O => \N__15172\,
            I => \N__15158\
        );

    \I__1717\ : InMux
    port map (
            O => \N__15171\,
            I => \N__15155\
        );

    \I__1716\ : Span4Mux_h
    port map (
            O => \N__15166\,
            I => \N__15152\
        );

    \I__1715\ : Span4Mux_v
    port map (
            O => \N__15163\,
            I => \N__15147\
        );

    \I__1714\ : Span4Mux_h
    port map (
            O => \N__15158\,
            I => \N__15147\
        );

    \I__1713\ : LocalMux
    port map (
            O => \N__15155\,
            I => \SYNTHESIZED_WIRE_4_1\
        );

    \I__1712\ : Odrv4
    port map (
            O => \N__15152\,
            I => \SYNTHESIZED_WIRE_4_1\
        );

    \I__1711\ : Odrv4
    port map (
            O => \N__15147\,
            I => \SYNTHESIZED_WIRE_4_1\
        );

    \I__1710\ : InMux
    port map (
            O => \N__15140\,
            I => \N__15136\
        );

    \I__1709\ : InMux
    port map (
            O => \N__15139\,
            I => \N__15133\
        );

    \I__1708\ : LocalMux
    port map (
            O => \N__15136\,
            I => \N__15127\
        );

    \I__1707\ : LocalMux
    port map (
            O => \N__15133\,
            I => \N__15127\
        );

    \I__1706\ : InMux
    port map (
            O => \N__15132\,
            I => \N__15124\
        );

    \I__1705\ : Span4Mux_h
    port map (
            O => \N__15127\,
            I => \N__15118\
        );

    \I__1704\ : LocalMux
    port map (
            O => \N__15124\,
            I => \N__15115\
        );

    \I__1703\ : InMux
    port map (
            O => \N__15123\,
            I => \N__15108\
        );

    \I__1702\ : InMux
    port map (
            O => \N__15122\,
            I => \N__15108\
        );

    \I__1701\ : InMux
    port map (
            O => \N__15121\,
            I => \N__15108\
        );

    \I__1700\ : Odrv4
    port map (
            O => \N__15118\,
            I => \SYNTHESIZED_WIRE_4_2\
        );

    \I__1699\ : Odrv4
    port map (
            O => \N__15115\,
            I => \SYNTHESIZED_WIRE_4_2\
        );

    \I__1698\ : LocalMux
    port map (
            O => \N__15108\,
            I => \SYNTHESIZED_WIRE_4_2\
        );

    \I__1697\ : CascadeMux
    port map (
            O => \N__15101\,
            I => \b2v_inst.dir_mem_316lt6_0_cascade_\
        );

    \I__1696\ : InMux
    port map (
            O => \N__15098\,
            I => \N__15095\
        );

    \I__1695\ : LocalMux
    port map (
            O => \N__15095\,
            I => \b2v_inst.dir_mem_316lt7\
        );

    \I__1694\ : InMux
    port map (
            O => \N__15092\,
            I => \N__15089\
        );

    \I__1693\ : LocalMux
    port map (
            O => \N__15089\,
            I => \N__15084\
        );

    \I__1692\ : InMux
    port map (
            O => \N__15088\,
            I => \N__15081\
        );

    \I__1691\ : InMux
    port map (
            O => \N__15087\,
            I => \N__15078\
        );

    \I__1690\ : Span4Mux_v
    port map (
            O => \N__15084\,
            I => \N__15073\
        );

    \I__1689\ : LocalMux
    port map (
            O => \N__15081\,
            I => \N__15073\
        );

    \I__1688\ : LocalMux
    port map (
            O => \N__15078\,
            I => \b2v_inst.un1_indice_cry_1_c_RNIUSJGZ0\
        );

    \I__1687\ : Odrv4
    port map (
            O => \N__15073\,
            I => \b2v_inst.un1_indice_cry_1_c_RNIUSJGZ0\
        );

    \I__1686\ : InMux
    port map (
            O => \N__15068\,
            I => \N__15065\
        );

    \I__1685\ : LocalMux
    port map (
            O => \N__15065\,
            I => \SYNTHESIZED_WIRE_4_fast_10\
        );

    \I__1684\ : InMux
    port map (
            O => \N__15062\,
            I => \N__15059\
        );

    \I__1683\ : LocalMux
    port map (
            O => \N__15059\,
            I => \N__15056\
        );

    \I__1682\ : Odrv4
    port map (
            O => \N__15056\,
            I => \SYNTHESIZED_WIRE_4_fast_9\
        );

    \I__1681\ : CascadeMux
    port map (
            O => \N__15053\,
            I => \b2v_inst.N_9_cascade_\
        );

    \I__1680\ : InMux
    port map (
            O => \N__15050\,
            I => \N__15047\
        );

    \I__1679\ : LocalMux
    port map (
            O => \N__15047\,
            I => \N__15044\
        );

    \I__1678\ : Span4Mux_h
    port map (
            O => \N__15044\,
            I => \N__15038\
        );

    \I__1677\ : InMux
    port map (
            O => \N__15043\,
            I => \N__15035\
        );

    \I__1676\ : InMux
    port map (
            O => \N__15042\,
            I => \N__15030\
        );

    \I__1675\ : InMux
    port map (
            O => \N__15041\,
            I => \N__15030\
        );

    \I__1674\ : Odrv4
    port map (
            O => \N__15038\,
            I => b2v_inst4_pix_count_int_fast_5
        );

    \I__1673\ : LocalMux
    port map (
            O => \N__15035\,
            I => b2v_inst4_pix_count_int_fast_5
        );

    \I__1672\ : LocalMux
    port map (
            O => \N__15030\,
            I => b2v_inst4_pix_count_int_fast_5
        );

    \I__1671\ : InMux
    port map (
            O => \N__15023\,
            I => \N__15020\
        );

    \I__1670\ : LocalMux
    port map (
            O => \N__15020\,
            I => \N__15014\
        );

    \I__1669\ : InMux
    port map (
            O => \N__15019\,
            I => \N__15007\
        );

    \I__1668\ : InMux
    port map (
            O => \N__15018\,
            I => \N__15007\
        );

    \I__1667\ : InMux
    port map (
            O => \N__15017\,
            I => \N__15007\
        );

    \I__1666\ : Odrv12
    port map (
            O => \N__15014\,
            I => b2v_inst4_pix_count_int_fast_6
        );

    \I__1665\ : LocalMux
    port map (
            O => \N__15007\,
            I => b2v_inst4_pix_count_int_fast_6
        );

    \I__1664\ : InMux
    port map (
            O => \N__15002\,
            I => \N__14999\
        );

    \I__1663\ : LocalMux
    port map (
            O => \N__14999\,
            I => \N__14996\
        );

    \I__1662\ : Odrv12
    port map (
            O => \N__14996\,
            I => \b2v_inst.un4_pix_count_intlto6_1_xZ0Z1\
        );

    \I__1661\ : InMux
    port map (
            O => \N__14993\,
            I => \N__14990\
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__14990\,
            I => \N__14987\
        );

    \I__1659\ : Span4Mux_h
    port map (
            O => \N__14987\,
            I => \N__14984\
        );

    \I__1658\ : Odrv4
    port map (
            O => \N__14984\,
            I => \b2v_inst.un4_pix_count_intlto6_1_xZ0Z0\
        );

    \I__1657\ : InMux
    port map (
            O => \N__14981\,
            I => \N__14978\
        );

    \I__1656\ : LocalMux
    port map (
            O => \N__14978\,
            I => \N__14975\
        );

    \I__1655\ : Span4Mux_h
    port map (
            O => \N__14975\,
            I => \N__14972\
        );

    \I__1654\ : Span4Mux_h
    port map (
            O => \N__14972\,
            I => \N__14969\
        );

    \I__1653\ : Odrv4
    port map (
            O => \N__14969\,
            I => \b2v_inst.un4_pix_count_intlto6_dZ0Z_1\
        );

    \I__1652\ : InMux
    port map (
            O => \N__14966\,
            I => \b2v_inst.un8_dir_mem_1_cry_4\
        );

    \I__1651\ : InMux
    port map (
            O => \N__14963\,
            I => \b2v_inst.un8_dir_mem_1_cry_5\
        );

    \I__1650\ : InMux
    port map (
            O => \N__14960\,
            I => \b2v_inst.un8_dir_mem_1_cry_6\
        );

    \I__1649\ : InMux
    port map (
            O => \N__14957\,
            I => \bfn_7_7_0_\
        );

    \I__1648\ : InMux
    port map (
            O => \N__14954\,
            I => \b2v_inst.un8_dir_mem_1_cry_8\
        );

    \I__1647\ : InMux
    port map (
            O => \N__14951\,
            I => \b2v_inst.un8_dir_mem_1_cry_9\
        );

    \I__1646\ : InMux
    port map (
            O => \N__14948\,
            I => \b2v_inst.un8_dir_mem_1_cry_10\
        );

    \I__1645\ : InMux
    port map (
            O => \N__14945\,
            I => \N__14942\
        );

    \I__1644\ : LocalMux
    port map (
            O => \N__14942\,
            I => \b2v_inst1.N_40\
        );

    \I__1643\ : InMux
    port map (
            O => \N__14939\,
            I => \b2v_inst.un8_dir_mem_1_cry_0\
        );

    \I__1642\ : InMux
    port map (
            O => \N__14936\,
            I => \b2v_inst.un8_dir_mem_1_cry_1\
        );

    \I__1641\ : InMux
    port map (
            O => \N__14933\,
            I => \b2v_inst.un8_dir_mem_1_cry_2\
        );

    \I__1640\ : InMux
    port map (
            O => \N__14930\,
            I => \b2v_inst.un8_dir_mem_1_cry_3\
        );

    \I__1639\ : IoInMux
    port map (
            O => \N__14927\,
            I => \N__14924\
        );

    \I__1638\ : LocalMux
    port map (
            O => \N__14924\,
            I => \N__14921\
        );

    \I__1637\ : Span4Mux_s1_h
    port map (
            O => \N__14921\,
            I => \N__14918\
        );

    \I__1636\ : Span4Mux_h
    port map (
            O => \N__14918\,
            I => \N__14915\
        );

    \I__1635\ : Span4Mux_h
    port map (
            O => \N__14915\,
            I => \N__14912\
        );

    \I__1634\ : Odrv4
    port map (
            O => \N__14912\,
            I => \b2v_inst.N_305_1\
        );

    \I__1633\ : CEMux
    port map (
            O => \N__14909\,
            I => \N__14906\
        );

    \I__1632\ : LocalMux
    port map (
            O => \N__14906\,
            I => \N__14903\
        );

    \I__1631\ : Span4Mux_v
    port map (
            O => \N__14903\,
            I => \N__14900\
        );

    \I__1630\ : Odrv4
    port map (
            O => \N__14900\,
            I => \b2v_inst.un1_state_36_0\
        );

    \I__1629\ : InMux
    port map (
            O => \N__14897\,
            I => \N__14892\
        );

    \I__1628\ : InMux
    port map (
            O => \N__14896\,
            I => \N__14889\
        );

    \I__1627\ : InMux
    port map (
            O => \N__14895\,
            I => \N__14886\
        );

    \I__1626\ : LocalMux
    port map (
            O => \N__14892\,
            I => \N__14881\
        );

    \I__1625\ : LocalMux
    port map (
            O => \N__14889\,
            I => \N__14881\
        );

    \I__1624\ : LocalMux
    port map (
            O => \N__14886\,
            I => \b2v_inst4.stateZ0Z_0\
        );

    \I__1623\ : Odrv12
    port map (
            O => \N__14881\,
            I => \b2v_inst4.stateZ0Z_0\
        );

    \I__1622\ : InMux
    port map (
            O => \N__14876\,
            I => \N__14872\
        );

    \I__1621\ : InMux
    port map (
            O => \N__14875\,
            I => \N__14869\
        );

    \I__1620\ : LocalMux
    port map (
            O => \N__14872\,
            I => \N__14866\
        );

    \I__1619\ : LocalMux
    port map (
            O => \N__14869\,
            I => \N__14861\
        );

    \I__1618\ : Span4Mux_h
    port map (
            O => \N__14866\,
            I => \N__14858\
        );

    \I__1617\ : InMux
    port map (
            O => \N__14865\,
            I => \N__14853\
        );

    \I__1616\ : InMux
    port map (
            O => \N__14864\,
            I => \N__14853\
        );

    \I__1615\ : Odrv12
    port map (
            O => \N__14861\,
            I => \SYNTHESIZED_WIRE_9\
        );

    \I__1614\ : Odrv4
    port map (
            O => \N__14858\,
            I => \SYNTHESIZED_WIRE_9\
        );

    \I__1613\ : LocalMux
    port map (
            O => \N__14853\,
            I => \SYNTHESIZED_WIRE_9\
        );

    \I__1612\ : CascadeMux
    port map (
            O => \N__14846\,
            I => \N__14843\
        );

    \I__1611\ : InMux
    port map (
            O => \N__14843\,
            I => \N__14840\
        );

    \I__1610\ : LocalMux
    port map (
            O => \N__14840\,
            I => \N__14837\
        );

    \I__1609\ : Odrv4
    port map (
            O => \N__14837\,
            I => \b2v_inst.un1_state_36_0_a2_0_1_mbZ0Z_1\
        );

    \I__1608\ : InMux
    port map (
            O => \N__14834\,
            I => \N__14825\
        );

    \I__1607\ : InMux
    port map (
            O => \N__14833\,
            I => \N__14825\
        );

    \I__1606\ : InMux
    port map (
            O => \N__14832\,
            I => \N__14825\
        );

    \I__1605\ : LocalMux
    port map (
            O => \N__14825\,
            I => \N__14822\
        );

    \I__1604\ : Span4Mux_h
    port map (
            O => \N__14822\,
            I => \N__14819\
        );

    \I__1603\ : Odrv4
    port map (
            O => \N__14819\,
            I => \b2v_inst4.un1_pix_count_int_cry_9_c_RNIB86JZ0\
        );

    \I__1602\ : InMux
    port map (
            O => \N__14816\,
            I => \N__14813\
        );

    \I__1601\ : LocalMux
    port map (
            O => \N__14813\,
            I => \N__14808\
        );

    \I__1600\ : InMux
    port map (
            O => \N__14812\,
            I => \N__14803\
        );

    \I__1599\ : InMux
    port map (
            O => \N__14811\,
            I => \N__14803\
        );

    \I__1598\ : Span4Mux_h
    port map (
            O => \N__14808\,
            I => \N__14800\
        );

    \I__1597\ : LocalMux
    port map (
            O => \N__14803\,
            I => \N__14797\
        );

    \I__1596\ : Odrv4
    port map (
            O => \N__14800\,
            I => \b2v_inst4.un1_pix_count_int_cry_8_c_RNI25BIZ0\
        );

    \I__1595\ : Odrv4
    port map (
            O => \N__14797\,
            I => \b2v_inst4.un1_pix_count_int_cry_8_c_RNI25BIZ0\
        );

    \I__1594\ : CascadeMux
    port map (
            O => \N__14792\,
            I => \N__14780\
        );

    \I__1593\ : InMux
    port map (
            O => \N__14791\,
            I => \N__14774\
        );

    \I__1592\ : InMux
    port map (
            O => \N__14790\,
            I => \N__14771\
        );

    \I__1591\ : InMux
    port map (
            O => \N__14789\,
            I => \N__14768\
        );

    \I__1590\ : InMux
    port map (
            O => \N__14788\,
            I => \N__14765\
        );

    \I__1589\ : InMux
    port map (
            O => \N__14787\,
            I => \N__14762\
        );

    \I__1588\ : InMux
    port map (
            O => \N__14786\,
            I => \N__14755\
        );

    \I__1587\ : InMux
    port map (
            O => \N__14785\,
            I => \N__14755\
        );

    \I__1586\ : InMux
    port map (
            O => \N__14784\,
            I => \N__14755\
        );

    \I__1585\ : InMux
    port map (
            O => \N__14783\,
            I => \N__14740\
        );

    \I__1584\ : InMux
    port map (
            O => \N__14780\,
            I => \N__14740\
        );

    \I__1583\ : InMux
    port map (
            O => \N__14779\,
            I => \N__14740\
        );

    \I__1582\ : InMux
    port map (
            O => \N__14778\,
            I => \N__14740\
        );

    \I__1581\ : InMux
    port map (
            O => \N__14777\,
            I => \N__14740\
        );

    \I__1580\ : LocalMux
    port map (
            O => \N__14774\,
            I => \N__14737\
        );

    \I__1579\ : LocalMux
    port map (
            O => \N__14771\,
            I => \N__14734\
        );

    \I__1578\ : LocalMux
    port map (
            O => \N__14768\,
            I => \N__14731\
        );

    \I__1577\ : LocalMux
    port map (
            O => \N__14765\,
            I => \N__14726\
        );

    \I__1576\ : LocalMux
    port map (
            O => \N__14762\,
            I => \N__14726\
        );

    \I__1575\ : LocalMux
    port map (
            O => \N__14755\,
            I => \N__14723\
        );

    \I__1574\ : InMux
    port map (
            O => \N__14754\,
            I => \N__14714\
        );

    \I__1573\ : InMux
    port map (
            O => \N__14753\,
            I => \N__14714\
        );

    \I__1572\ : InMux
    port map (
            O => \N__14752\,
            I => \N__14714\
        );

    \I__1571\ : InMux
    port map (
            O => \N__14751\,
            I => \N__14714\
        );

    \I__1570\ : LocalMux
    port map (
            O => \N__14740\,
            I => \N__14711\
        );

    \I__1569\ : Span4Mux_h
    port map (
            O => \N__14737\,
            I => \N__14708\
        );

    \I__1568\ : Span4Mux_h
    port map (
            O => \N__14734\,
            I => \N__14705\
        );

    \I__1567\ : Span4Mux_h
    port map (
            O => \N__14731\,
            I => \N__14698\
        );

    \I__1566\ : Span4Mux_h
    port map (
            O => \N__14726\,
            I => \N__14698\
        );

    \I__1565\ : Span4Mux_h
    port map (
            O => \N__14723\,
            I => \N__14698\
        );

    \I__1564\ : LocalMux
    port map (
            O => \N__14714\,
            I => \b2v_inst4.un1_pix_count_int_0_sqmuxa_0\
        );

    \I__1563\ : Odrv4
    port map (
            O => \N__14711\,
            I => \b2v_inst4.un1_pix_count_int_0_sqmuxa_0\
        );

    \I__1562\ : Odrv4
    port map (
            O => \N__14708\,
            I => \b2v_inst4.un1_pix_count_int_0_sqmuxa_0\
        );

    \I__1561\ : Odrv4
    port map (
            O => \N__14705\,
            I => \b2v_inst4.un1_pix_count_int_0_sqmuxa_0\
        );

    \I__1560\ : Odrv4
    port map (
            O => \N__14698\,
            I => \b2v_inst4.un1_pix_count_int_0_sqmuxa_0\
        );

    \I__1559\ : InMux
    port map (
            O => \N__14687\,
            I => \N__14684\
        );

    \I__1558\ : LocalMux
    port map (
            O => \N__14684\,
            I => \N__14680\
        );

    \I__1557\ : InMux
    port map (
            O => \N__14683\,
            I => \N__14677\
        );

    \I__1556\ : Span4Mux_h
    port map (
            O => \N__14680\,
            I => \N__14674\
        );

    \I__1555\ : LocalMux
    port map (
            O => \N__14677\,
            I => \N__14671\
        );

    \I__1554\ : Odrv4
    port map (
            O => \N__14674\,
            I => \b2v_inst4.un1_pix_count_int_cry_10_c_RNIKMUJZ0\
        );

    \I__1553\ : Odrv4
    port map (
            O => \N__14671\,
            I => \b2v_inst4.un1_pix_count_int_cry_10_c_RNIKMUJZ0\
        );

    \I__1552\ : InMux
    port map (
            O => \N__14666\,
            I => \N__14663\
        );

    \I__1551\ : LocalMux
    port map (
            O => \N__14663\,
            I => \N__14660\
        );

    \I__1550\ : Odrv4
    port map (
            O => \N__14660\,
            I => \b2v_inst.ignorar_ancho_1_RNOZ0Z_0\
        );

    \I__1549\ : CascadeMux
    port map (
            O => \N__14657\,
            I => \b2v_inst.N_482_cascade_\
        );

    \I__1548\ : CEMux
    port map (
            O => \N__14654\,
            I => \N__14651\
        );

    \I__1547\ : LocalMux
    port map (
            O => \N__14651\,
            I => \N__14648\
        );

    \I__1546\ : Odrv4
    port map (
            O => \N__14648\,
            I => \b2v_inst.un1_state_34_0\
        );

    \I__1545\ : InMux
    port map (
            O => \N__14645\,
            I => \N__14642\
        );

    \I__1544\ : LocalMux
    port map (
            O => \N__14642\,
            I => \N__14637\
        );

    \I__1543\ : InMux
    port map (
            O => \N__14641\,
            I => \N__14632\
        );

    \I__1542\ : InMux
    port map (
            O => \N__14640\,
            I => \N__14632\
        );

    \I__1541\ : Span4Mux_v
    port map (
            O => \N__14637\,
            I => \N__14629\
        );

    \I__1540\ : LocalMux
    port map (
            O => \N__14632\,
            I => \N__14626\
        );

    \I__1539\ : Odrv4
    port map (
            O => \N__14629\,
            I => \b2v_inst.un1_cuenta_pixel_cry_8_c_RNIMU4IZ0\
        );

    \I__1538\ : Odrv4
    port map (
            O => \N__14626\,
            I => \b2v_inst.un1_cuenta_pixel_cry_8_c_RNIMU4IZ0\
        );

    \I__1537\ : InMux
    port map (
            O => \N__14621\,
            I => \N__14618\
        );

    \I__1536\ : LocalMux
    port map (
            O => \N__14618\,
            I => \N__14613\
        );

    \I__1535\ : InMux
    port map (
            O => \N__14617\,
            I => \N__14610\
        );

    \I__1534\ : InMux
    port map (
            O => \N__14616\,
            I => \N__14607\
        );

    \I__1533\ : Span4Mux_h
    port map (
            O => \N__14613\,
            I => \N__14604\
        );

    \I__1532\ : LocalMux
    port map (
            O => \N__14610\,
            I => \N__14601\
        );

    \I__1531\ : LocalMux
    port map (
            O => \N__14607\,
            I => \b2v_inst.cuenta_pixel_RNIVBL9Z0Z_10\
        );

    \I__1530\ : Odrv4
    port map (
            O => \N__14604\,
            I => \b2v_inst.cuenta_pixel_RNIVBL9Z0Z_10\
        );

    \I__1529\ : Odrv4
    port map (
            O => \N__14601\,
            I => \b2v_inst.cuenta_pixel_RNIVBL9Z0Z_10\
        );

    \I__1528\ : CascadeMux
    port map (
            O => \N__14594\,
            I => \N__14591\
        );

    \I__1527\ : InMux
    port map (
            O => \N__14591\,
            I => \N__14587\
        );

    \I__1526\ : CascadeMux
    port map (
            O => \N__14590\,
            I => \N__14584\
        );

    \I__1525\ : LocalMux
    port map (
            O => \N__14587\,
            I => \N__14580\
        );

    \I__1524\ : InMux
    port map (
            O => \N__14584\,
            I => \N__14577\
        );

    \I__1523\ : InMux
    port map (
            O => \N__14583\,
            I => \N__14574\
        );

    \I__1522\ : Span4Mux_h
    port map (
            O => \N__14580\,
            I => \N__14571\
        );

    \I__1521\ : LocalMux
    port map (
            O => \N__14577\,
            I => \N__14568\
        );

    \I__1520\ : LocalMux
    port map (
            O => \N__14574\,
            I => \b2v_inst.un1_cuenta_pixel_cry_7_c_RNIKR3IZ0\
        );

    \I__1519\ : Odrv4
    port map (
            O => \N__14571\,
            I => \b2v_inst.un1_cuenta_pixel_cry_7_c_RNIKR3IZ0\
        );

    \I__1518\ : Odrv4
    port map (
            O => \N__14568\,
            I => \b2v_inst.un1_cuenta_pixel_cry_7_c_RNIKR3IZ0\
        );

    \I__1517\ : InMux
    port map (
            O => \N__14561\,
            I => \N__14558\
        );

    \I__1516\ : LocalMux
    port map (
            O => \N__14558\,
            I => \N__14554\
        );

    \I__1515\ : InMux
    port map (
            O => \N__14557\,
            I => \N__14551\
        );

    \I__1514\ : Span4Mux_h
    port map (
            O => \N__14554\,
            I => \N__14548\
        );

    \I__1513\ : LocalMux
    port map (
            O => \N__14551\,
            I => \b2v_inst.cuenta_pixel_5_i_a2_1_1_0_5\
        );

    \I__1512\ : Odrv4
    port map (
            O => \N__14548\,
            I => \b2v_inst.cuenta_pixel_5_i_a2_1_1_0_5\
        );

    \I__1511\ : InMux
    port map (
            O => \N__14543\,
            I => \N__14540\
        );

    \I__1510\ : LocalMux
    port map (
            O => \N__14540\,
            I => \N__14536\
        );

    \I__1509\ : InMux
    port map (
            O => \N__14539\,
            I => \N__14533\
        );

    \I__1508\ : Odrv4
    port map (
            O => \N__14536\,
            I => \b2v_inst.N_325\
        );

    \I__1507\ : LocalMux
    port map (
            O => \N__14533\,
            I => \b2v_inst.N_325\
        );

    \I__1506\ : InMux
    port map (
            O => \N__14528\,
            I => \N__14525\
        );

    \I__1505\ : LocalMux
    port map (
            O => \N__14525\,
            I => \N__14522\
        );

    \I__1504\ : Odrv4
    port map (
            O => \N__14522\,
            I => \b2v_inst.un1_state_36_0_rn_1\
        );

    \I__1503\ : InMux
    port map (
            O => \N__14519\,
            I => \N__14516\
        );

    \I__1502\ : LocalMux
    port map (
            O => \N__14516\,
            I => \N__14513\
        );

    \I__1501\ : Odrv4
    port map (
            O => \N__14513\,
            I => \b2v_inst.un1_state_36_0_sn\
        );

    \I__1500\ : CascadeMux
    port map (
            O => \N__14510\,
            I => \b2v_inst.N_325_cascade_\
        );

    \I__1499\ : InMux
    port map (
            O => \N__14507\,
            I => \b2v_inst.un1_indice_cry_6\
        );

    \I__1498\ : InMux
    port map (
            O => \N__14504\,
            I => \b2v_inst.un1_indice_cry_7\
        );

    \I__1497\ : InMux
    port map (
            O => \N__14501\,
            I => \bfn_6_7_0_\
        );

    \I__1496\ : InMux
    port map (
            O => \N__14498\,
            I => \b2v_inst.un1_indice_cry_9\
        );

    \I__1495\ : InMux
    port map (
            O => \N__14495\,
            I => \b2v_inst.un1_indice_cry_10\
        );

    \I__1494\ : InMux
    port map (
            O => \N__14492\,
            I => \N__14489\
        );

    \I__1493\ : LocalMux
    port map (
            O => \N__14489\,
            I => \b2v_inst.ignorar_ancho_1_RNOZ0Z_1\
        );

    \I__1492\ : InMux
    port map (
            O => \N__14486\,
            I => \N__14483\
        );

    \I__1491\ : LocalMux
    port map (
            O => \N__14483\,
            I => \b2v_inst.ignorar_ancho_1_RNOZ0Z_2\
        );

    \I__1490\ : InMux
    port map (
            O => \N__14480\,
            I => \b2v_inst.un2_dir_mem_3_cry_2\
        );

    \I__1489\ : InMux
    port map (
            O => \N__14477\,
            I => \b2v_inst.un2_dir_mem_3_cry_3\
        );

    \I__1488\ : InMux
    port map (
            O => \N__14474\,
            I => \b2v_inst.un2_dir_mem_3_cry_4\
        );

    \I__1487\ : InMux
    port map (
            O => \N__14471\,
            I => \b2v_inst.un1_indice_cry_1\
        );

    \I__1486\ : InMux
    port map (
            O => \N__14468\,
            I => \b2v_inst.un1_indice_cry_2\
        );

    \I__1485\ : InMux
    port map (
            O => \N__14465\,
            I => \b2v_inst.un1_indice_cry_3\
        );

    \I__1484\ : InMux
    port map (
            O => \N__14462\,
            I => \b2v_inst.un1_indice_cry_4\
        );

    \I__1483\ : InMux
    port map (
            O => \N__14459\,
            I => \b2v_inst.un1_indice_cry_5\
        );

    \I__1482\ : InMux
    port map (
            O => \N__14456\,
            I => \b2v_inst4.un1_pix_count_int_cry_18\
        );

    \I__1481\ : CascadeMux
    port map (
            O => \N__14453\,
            I => \N__14449\
        );

    \I__1480\ : CascadeMux
    port map (
            O => \N__14452\,
            I => \N__14446\
        );

    \I__1479\ : CascadeBuf
    port map (
            O => \N__14449\,
            I => \N__14443\
        );

    \I__1478\ : CascadeBuf
    port map (
            O => \N__14446\,
            I => \N__14440\
        );

    \I__1477\ : CascadeMux
    port map (
            O => \N__14443\,
            I => \N__14437\
        );

    \I__1476\ : CascadeMux
    port map (
            O => \N__14440\,
            I => \N__14434\
        );

    \I__1475\ : CascadeBuf
    port map (
            O => \N__14437\,
            I => \N__14431\
        );

    \I__1474\ : CascadeBuf
    port map (
            O => \N__14434\,
            I => \N__14428\
        );

    \I__1473\ : CascadeMux
    port map (
            O => \N__14431\,
            I => \N__14425\
        );

    \I__1472\ : CascadeMux
    port map (
            O => \N__14428\,
            I => \N__14422\
        );

    \I__1471\ : CascadeBuf
    port map (
            O => \N__14425\,
            I => \N__14419\
        );

    \I__1470\ : CascadeBuf
    port map (
            O => \N__14422\,
            I => \N__14416\
        );

    \I__1469\ : CascadeMux
    port map (
            O => \N__14419\,
            I => \N__14413\
        );

    \I__1468\ : CascadeMux
    port map (
            O => \N__14416\,
            I => \N__14410\
        );

    \I__1467\ : CascadeBuf
    port map (
            O => \N__14413\,
            I => \N__14407\
        );

    \I__1466\ : CascadeBuf
    port map (
            O => \N__14410\,
            I => \N__14404\
        );

    \I__1465\ : CascadeMux
    port map (
            O => \N__14407\,
            I => \N__14401\
        );

    \I__1464\ : CascadeMux
    port map (
            O => \N__14404\,
            I => \N__14398\
        );

    \I__1463\ : CascadeBuf
    port map (
            O => \N__14401\,
            I => \N__14395\
        );

    \I__1462\ : CascadeBuf
    port map (
            O => \N__14398\,
            I => \N__14392\
        );

    \I__1461\ : CascadeMux
    port map (
            O => \N__14395\,
            I => \N__14389\
        );

    \I__1460\ : CascadeMux
    port map (
            O => \N__14392\,
            I => \N__14386\
        );

    \I__1459\ : CascadeBuf
    port map (
            O => \N__14389\,
            I => \N__14383\
        );

    \I__1458\ : CascadeBuf
    port map (
            O => \N__14386\,
            I => \N__14380\
        );

    \I__1457\ : CascadeMux
    port map (
            O => \N__14383\,
            I => \N__14377\
        );

    \I__1456\ : CascadeMux
    port map (
            O => \N__14380\,
            I => \N__14374\
        );

    \I__1455\ : InMux
    port map (
            O => \N__14377\,
            I => \N__14371\
        );

    \I__1454\ : InMux
    port map (
            O => \N__14374\,
            I => \N__14368\
        );

    \I__1453\ : LocalMux
    port map (
            O => \N__14371\,
            I => \N__14365\
        );

    \I__1452\ : LocalMux
    port map (
            O => \N__14368\,
            I => \SYNTHESIZED_WIRE_12_1\
        );

    \I__1451\ : Odrv4
    port map (
            O => \N__14365\,
            I => \SYNTHESIZED_WIRE_12_1\
        );

    \I__1450\ : CascadeMux
    port map (
            O => \N__14360\,
            I => \N__14357\
        );

    \I__1449\ : CascadeBuf
    port map (
            O => \N__14357\,
            I => \N__14353\
        );

    \I__1448\ : CascadeMux
    port map (
            O => \N__14356\,
            I => \N__14350\
        );

    \I__1447\ : CascadeMux
    port map (
            O => \N__14353\,
            I => \N__14347\
        );

    \I__1446\ : CascadeBuf
    port map (
            O => \N__14350\,
            I => \N__14344\
        );

    \I__1445\ : CascadeBuf
    port map (
            O => \N__14347\,
            I => \N__14341\
        );

    \I__1444\ : CascadeMux
    port map (
            O => \N__14344\,
            I => \N__14338\
        );

    \I__1443\ : CascadeMux
    port map (
            O => \N__14341\,
            I => \N__14335\
        );

    \I__1442\ : CascadeBuf
    port map (
            O => \N__14338\,
            I => \N__14332\
        );

    \I__1441\ : CascadeBuf
    port map (
            O => \N__14335\,
            I => \N__14329\
        );

    \I__1440\ : CascadeMux
    port map (
            O => \N__14332\,
            I => \N__14326\
        );

    \I__1439\ : CascadeMux
    port map (
            O => \N__14329\,
            I => \N__14323\
        );

    \I__1438\ : CascadeBuf
    port map (
            O => \N__14326\,
            I => \N__14320\
        );

    \I__1437\ : CascadeBuf
    port map (
            O => \N__14323\,
            I => \N__14317\
        );

    \I__1436\ : CascadeMux
    port map (
            O => \N__14320\,
            I => \N__14314\
        );

    \I__1435\ : CascadeMux
    port map (
            O => \N__14317\,
            I => \N__14311\
        );

    \I__1434\ : CascadeBuf
    port map (
            O => \N__14314\,
            I => \N__14308\
        );

    \I__1433\ : CascadeBuf
    port map (
            O => \N__14311\,
            I => \N__14305\
        );

    \I__1432\ : CascadeMux
    port map (
            O => \N__14308\,
            I => \N__14302\
        );

    \I__1431\ : CascadeMux
    port map (
            O => \N__14305\,
            I => \N__14299\
        );

    \I__1430\ : CascadeBuf
    port map (
            O => \N__14302\,
            I => \N__14296\
        );

    \I__1429\ : CascadeBuf
    port map (
            O => \N__14299\,
            I => \N__14293\
        );

    \I__1428\ : CascadeMux
    port map (
            O => \N__14296\,
            I => \N__14290\
        );

    \I__1427\ : CascadeMux
    port map (
            O => \N__14293\,
            I => \N__14287\
        );

    \I__1426\ : CascadeBuf
    port map (
            O => \N__14290\,
            I => \N__14284\
        );

    \I__1425\ : InMux
    port map (
            O => \N__14287\,
            I => \N__14281\
        );

    \I__1424\ : CascadeMux
    port map (
            O => \N__14284\,
            I => \N__14278\
        );

    \I__1423\ : LocalMux
    port map (
            O => \N__14281\,
            I => \N__14275\
        );

    \I__1422\ : InMux
    port map (
            O => \N__14278\,
            I => \N__14272\
        );

    \I__1421\ : Span4Mux_h
    port map (
            O => \N__14275\,
            I => \N__14269\
        );

    \I__1420\ : LocalMux
    port map (
            O => \N__14272\,
            I => \SYNTHESIZED_WIRE_12_7\
        );

    \I__1419\ : Odrv4
    port map (
            O => \N__14269\,
            I => \SYNTHESIZED_WIRE_12_7\
        );

    \I__1418\ : CascadeMux
    port map (
            O => \N__14264\,
            I => \N__14260\
        );

    \I__1417\ : CascadeMux
    port map (
            O => \N__14263\,
            I => \N__14257\
        );

    \I__1416\ : CascadeBuf
    port map (
            O => \N__14260\,
            I => \N__14254\
        );

    \I__1415\ : CascadeBuf
    port map (
            O => \N__14257\,
            I => \N__14251\
        );

    \I__1414\ : CascadeMux
    port map (
            O => \N__14254\,
            I => \N__14248\
        );

    \I__1413\ : CascadeMux
    port map (
            O => \N__14251\,
            I => \N__14245\
        );

    \I__1412\ : CascadeBuf
    port map (
            O => \N__14248\,
            I => \N__14242\
        );

    \I__1411\ : CascadeBuf
    port map (
            O => \N__14245\,
            I => \N__14239\
        );

    \I__1410\ : CascadeMux
    port map (
            O => \N__14242\,
            I => \N__14236\
        );

    \I__1409\ : CascadeMux
    port map (
            O => \N__14239\,
            I => \N__14233\
        );

    \I__1408\ : CascadeBuf
    port map (
            O => \N__14236\,
            I => \N__14230\
        );

    \I__1407\ : CascadeBuf
    port map (
            O => \N__14233\,
            I => \N__14227\
        );

    \I__1406\ : CascadeMux
    port map (
            O => \N__14230\,
            I => \N__14224\
        );

    \I__1405\ : CascadeMux
    port map (
            O => \N__14227\,
            I => \N__14221\
        );

    \I__1404\ : CascadeBuf
    port map (
            O => \N__14224\,
            I => \N__14218\
        );

    \I__1403\ : CascadeBuf
    port map (
            O => \N__14221\,
            I => \N__14215\
        );

    \I__1402\ : CascadeMux
    port map (
            O => \N__14218\,
            I => \N__14212\
        );

    \I__1401\ : CascadeMux
    port map (
            O => \N__14215\,
            I => \N__14209\
        );

    \I__1400\ : CascadeBuf
    port map (
            O => \N__14212\,
            I => \N__14206\
        );

    \I__1399\ : CascadeBuf
    port map (
            O => \N__14209\,
            I => \N__14203\
        );

    \I__1398\ : CascadeMux
    port map (
            O => \N__14206\,
            I => \N__14200\
        );

    \I__1397\ : CascadeMux
    port map (
            O => \N__14203\,
            I => \N__14197\
        );

    \I__1396\ : CascadeBuf
    port map (
            O => \N__14200\,
            I => \N__14194\
        );

    \I__1395\ : CascadeBuf
    port map (
            O => \N__14197\,
            I => \N__14191\
        );

    \I__1394\ : CascadeMux
    port map (
            O => \N__14194\,
            I => \N__14188\
        );

    \I__1393\ : CascadeMux
    port map (
            O => \N__14191\,
            I => \N__14185\
        );

    \I__1392\ : InMux
    port map (
            O => \N__14188\,
            I => \N__14182\
        );

    \I__1391\ : InMux
    port map (
            O => \N__14185\,
            I => \N__14179\
        );

    \I__1390\ : LocalMux
    port map (
            O => \N__14182\,
            I => \N__14176\
        );

    \I__1389\ : LocalMux
    port map (
            O => \N__14179\,
            I => \SYNTHESIZED_WIRE_12_0\
        );

    \I__1388\ : Odrv4
    port map (
            O => \N__14176\,
            I => \SYNTHESIZED_WIRE_12_0\
        );

    \I__1387\ : CascadeMux
    port map (
            O => \N__14171\,
            I => \N__14167\
        );

    \I__1386\ : CascadeMux
    port map (
            O => \N__14170\,
            I => \N__14164\
        );

    \I__1385\ : CascadeBuf
    port map (
            O => \N__14167\,
            I => \N__14161\
        );

    \I__1384\ : CascadeBuf
    port map (
            O => \N__14164\,
            I => \N__14158\
        );

    \I__1383\ : CascadeMux
    port map (
            O => \N__14161\,
            I => \N__14155\
        );

    \I__1382\ : CascadeMux
    port map (
            O => \N__14158\,
            I => \N__14152\
        );

    \I__1381\ : CascadeBuf
    port map (
            O => \N__14155\,
            I => \N__14149\
        );

    \I__1380\ : CascadeBuf
    port map (
            O => \N__14152\,
            I => \N__14146\
        );

    \I__1379\ : CascadeMux
    port map (
            O => \N__14149\,
            I => \N__14143\
        );

    \I__1378\ : CascadeMux
    port map (
            O => \N__14146\,
            I => \N__14140\
        );

    \I__1377\ : CascadeBuf
    port map (
            O => \N__14143\,
            I => \N__14137\
        );

    \I__1376\ : CascadeBuf
    port map (
            O => \N__14140\,
            I => \N__14134\
        );

    \I__1375\ : CascadeMux
    port map (
            O => \N__14137\,
            I => \N__14131\
        );

    \I__1374\ : CascadeMux
    port map (
            O => \N__14134\,
            I => \N__14128\
        );

    \I__1373\ : CascadeBuf
    port map (
            O => \N__14131\,
            I => \N__14125\
        );

    \I__1372\ : CascadeBuf
    port map (
            O => \N__14128\,
            I => \N__14122\
        );

    \I__1371\ : CascadeMux
    port map (
            O => \N__14125\,
            I => \N__14119\
        );

    \I__1370\ : CascadeMux
    port map (
            O => \N__14122\,
            I => \N__14116\
        );

    \I__1369\ : CascadeBuf
    port map (
            O => \N__14119\,
            I => \N__14113\
        );

    \I__1368\ : CascadeBuf
    port map (
            O => \N__14116\,
            I => \N__14110\
        );

    \I__1367\ : CascadeMux
    port map (
            O => \N__14113\,
            I => \N__14107\
        );

    \I__1366\ : CascadeMux
    port map (
            O => \N__14110\,
            I => \N__14104\
        );

    \I__1365\ : CascadeBuf
    port map (
            O => \N__14107\,
            I => \N__14101\
        );

    \I__1364\ : CascadeBuf
    port map (
            O => \N__14104\,
            I => \N__14098\
        );

    \I__1363\ : CascadeMux
    port map (
            O => \N__14101\,
            I => \N__14095\
        );

    \I__1362\ : CascadeMux
    port map (
            O => \N__14098\,
            I => \N__14092\
        );

    \I__1361\ : InMux
    port map (
            O => \N__14095\,
            I => \N__14089\
        );

    \I__1360\ : InMux
    port map (
            O => \N__14092\,
            I => \N__14086\
        );

    \I__1359\ : LocalMux
    port map (
            O => \N__14089\,
            I => \SYNTHESIZED_WIRE_12_8\
        );

    \I__1358\ : LocalMux
    port map (
            O => \N__14086\,
            I => \SYNTHESIZED_WIRE_12_8\
        );

    \I__1357\ : InMux
    port map (
            O => \N__14081\,
            I => \b2v_inst.un2_dir_mem_3_cry_0\
        );

    \I__1356\ : InMux
    port map (
            O => \N__14078\,
            I => \b2v_inst.un2_dir_mem_3_cry_1\
        );

    \I__1355\ : InMux
    port map (
            O => \N__14075\,
            I => \b2v_inst4.un1_pix_count_int_cry_9\
        );

    \I__1354\ : InMux
    port map (
            O => \N__14072\,
            I => \b2v_inst4.un1_pix_count_int_cry_10\
        );

    \I__1353\ : InMux
    port map (
            O => \N__14069\,
            I => \N__14063\
        );

    \I__1352\ : InMux
    port map (
            O => \N__14068\,
            I => \N__14063\
        );

    \I__1351\ : LocalMux
    port map (
            O => \N__14063\,
            I => \N__14060\
        );

    \I__1350\ : Odrv4
    port map (
            O => \N__14060\,
            I => \b2v_inst4.un1_pix_count_int_cry_11_c_RNIMPVJZ0\
        );

    \I__1349\ : InMux
    port map (
            O => \N__14057\,
            I => \b2v_inst4.un1_pix_count_int_cry_11\
        );

    \I__1348\ : InMux
    port map (
            O => \N__14054\,
            I => \b2v_inst4.un1_pix_count_int_cry_12\
        );

    \I__1347\ : InMux
    port map (
            O => \N__14051\,
            I => \b2v_inst4.un1_pix_count_int_cry_13\
        );

    \I__1346\ : InMux
    port map (
            O => \N__14048\,
            I => \b2v_inst4.un1_pix_count_int_cry_14\
        );

    \I__1345\ : InMux
    port map (
            O => \N__14045\,
            I => \bfn_5_15_0_\
        );

    \I__1344\ : InMux
    port map (
            O => \N__14042\,
            I => \b2v_inst4.un1_pix_count_int_cry_16\
        );

    \I__1343\ : InMux
    port map (
            O => \N__14039\,
            I => \b2v_inst4.un1_pix_count_int_cry_17\
        );

    \I__1342\ : InMux
    port map (
            O => \N__14036\,
            I => \N__14033\
        );

    \I__1341\ : LocalMux
    port map (
            O => \N__14033\,
            I => \N__14029\
        );

    \I__1340\ : InMux
    port map (
            O => \N__14032\,
            I => \N__14026\
        );

    \I__1339\ : Span4Mux_v
    port map (
            O => \N__14029\,
            I => \N__14021\
        );

    \I__1338\ : LocalMux
    port map (
            O => \N__14026\,
            I => \N__14021\
        );

    \I__1337\ : Span4Mux_h
    port map (
            O => \N__14021\,
            I => \N__14018\
        );

    \I__1336\ : Odrv4
    port map (
            O => \N__14018\,
            I => \b2v_inst4.un1_pix_count_int_cry_0_c_RNIIC2IZ0\
        );

    \I__1335\ : InMux
    port map (
            O => \N__14015\,
            I => \b2v_inst4.un1_pix_count_int_cry_0\
        );

    \I__1334\ : InMux
    port map (
            O => \N__14012\,
            I => \N__14009\
        );

    \I__1333\ : LocalMux
    port map (
            O => \N__14009\,
            I => \N__14005\
        );

    \I__1332\ : InMux
    port map (
            O => \N__14008\,
            I => \N__14002\
        );

    \I__1331\ : Span4Mux_v
    port map (
            O => \N__14005\,
            I => \N__13997\
        );

    \I__1330\ : LocalMux
    port map (
            O => \N__14002\,
            I => \N__13997\
        );

    \I__1329\ : Span4Mux_h
    port map (
            O => \N__13997\,
            I => \N__13994\
        );

    \I__1328\ : Odrv4
    port map (
            O => \N__13994\,
            I => \b2v_inst4.un1_pix_count_int_cry_1_c_RNIKF3IZ0\
        );

    \I__1327\ : InMux
    port map (
            O => \N__13991\,
            I => \b2v_inst4.un1_pix_count_int_cry_1\
        );

    \I__1326\ : InMux
    port map (
            O => \N__13988\,
            I => \N__13982\
        );

    \I__1325\ : InMux
    port map (
            O => \N__13987\,
            I => \N__13982\
        );

    \I__1324\ : LocalMux
    port map (
            O => \N__13982\,
            I => \N__13979\
        );

    \I__1323\ : Odrv12
    port map (
            O => \N__13979\,
            I => \b2v_inst4.un1_pix_count_int_cry_2_c_RNIMI4IZ0\
        );

    \I__1322\ : InMux
    port map (
            O => \N__13976\,
            I => \b2v_inst4.un1_pix_count_int_cry_2\
        );

    \I__1321\ : InMux
    port map (
            O => \N__13973\,
            I => \b2v_inst4.un1_pix_count_int_cry_3\
        );

    \I__1320\ : InMux
    port map (
            O => \N__13970\,
            I => \N__13964\
        );

    \I__1319\ : InMux
    port map (
            O => \N__13969\,
            I => \N__13964\
        );

    \I__1318\ : LocalMux
    port map (
            O => \N__13964\,
            I => \N__13961\
        );

    \I__1317\ : Span4Mux_h
    port map (
            O => \N__13961\,
            I => \N__13958\
        );

    \I__1316\ : Odrv4
    port map (
            O => \N__13958\,
            I => \b2v_inst4.un1_pix_count_int_cry_4_c_RNIQO6IZ0\
        );

    \I__1315\ : InMux
    port map (
            O => \N__13955\,
            I => \b2v_inst4.un1_pix_count_int_cry_4\
        );

    \I__1314\ : InMux
    port map (
            O => \N__13952\,
            I => \N__13949\
        );

    \I__1313\ : LocalMux
    port map (
            O => \N__13949\,
            I => \N__13945\
        );

    \I__1312\ : InMux
    port map (
            O => \N__13948\,
            I => \N__13942\
        );

    \I__1311\ : Span4Mux_v
    port map (
            O => \N__13945\,
            I => \N__13937\
        );

    \I__1310\ : LocalMux
    port map (
            O => \N__13942\,
            I => \N__13937\
        );

    \I__1309\ : Span4Mux_h
    port map (
            O => \N__13937\,
            I => \N__13934\
        );

    \I__1308\ : Odrv4
    port map (
            O => \N__13934\,
            I => \b2v_inst4.un1_pix_count_int_cry_5_c_RNISR7IZ0\
        );

    \I__1307\ : InMux
    port map (
            O => \N__13931\,
            I => \b2v_inst4.un1_pix_count_int_cry_5\
        );

    \I__1306\ : InMux
    port map (
            O => \N__13928\,
            I => \b2v_inst4.un1_pix_count_int_cry_6\
        );

    \I__1305\ : InMux
    port map (
            O => \N__13925\,
            I => \bfn_5_14_0_\
        );

    \I__1304\ : InMux
    port map (
            O => \N__13922\,
            I => \b2v_inst4.un1_pix_count_int_cry_8\
        );

    \I__1303\ : CascadeMux
    port map (
            O => \N__13919\,
            I => \N__13915\
        );

    \I__1302\ : InMux
    port map (
            O => \N__13918\,
            I => \N__13907\
        );

    \I__1301\ : InMux
    port map (
            O => \N__13915\,
            I => \N__13907\
        );

    \I__1300\ : InMux
    port map (
            O => \N__13914\,
            I => \N__13907\
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__13907\,
            I => \N__13904\
        );

    \I__1298\ : Odrv12
    port map (
            O => \N__13904\,
            I => \b2v_inst.un1_cuenta_pixel_cry_3_c_RNICFVHZ0\
        );

    \I__1297\ : CascadeMux
    port map (
            O => \N__13901\,
            I => \N__13898\
        );

    \I__1296\ : InMux
    port map (
            O => \N__13898\,
            I => \N__13895\
        );

    \I__1295\ : LocalMux
    port map (
            O => \N__13895\,
            I => \N__13892\
        );

    \I__1294\ : Odrv4
    port map (
            O => \N__13892\,
            I => \b2v_inst.cuenta_pixelZ0Z_4\
        );

    \I__1293\ : CascadeMux
    port map (
            O => \N__13889\,
            I => \N__13886\
        );

    \I__1292\ : InMux
    port map (
            O => \N__13886\,
            I => \N__13883\
        );

    \I__1291\ : LocalMux
    port map (
            O => \N__13883\,
            I => \N__13880\
        );

    \I__1290\ : Odrv12
    port map (
            O => \N__13880\,
            I => \b2v_inst.un7_pix_count_int_0_I_9_c_RNOZ0\
        );

    \I__1289\ : InMux
    port map (
            O => \N__13877\,
            I => \N__13874\
        );

    \I__1288\ : LocalMux
    port map (
            O => \N__13874\,
            I => \b2v_inst.pix_count_anteriorZ0Z_10\
        );

    \I__1287\ : CascadeMux
    port map (
            O => \N__13871\,
            I => \N__13868\
        );

    \I__1286\ : InMux
    port map (
            O => \N__13868\,
            I => \N__13865\
        );

    \I__1285\ : LocalMux
    port map (
            O => \N__13865\,
            I => \b2v_inst.pix_count_anteriorZ0Z_11\
        );

    \I__1284\ : InMux
    port map (
            O => \N__13862\,
            I => \N__13859\
        );

    \I__1283\ : LocalMux
    port map (
            O => \N__13859\,
            I => \N__13856\
        );

    \I__1282\ : Odrv4
    port map (
            O => \N__13856\,
            I => \b2v_inst.pix_count_anteriorZ0Z_17\
        );

    \I__1281\ : CEMux
    port map (
            O => \N__13853\,
            I => \N__13823\
        );

    \I__1280\ : CEMux
    port map (
            O => \N__13852\,
            I => \N__13823\
        );

    \I__1279\ : CEMux
    port map (
            O => \N__13851\,
            I => \N__13823\
        );

    \I__1278\ : CEMux
    port map (
            O => \N__13850\,
            I => \N__13823\
        );

    \I__1277\ : CEMux
    port map (
            O => \N__13849\,
            I => \N__13823\
        );

    \I__1276\ : CEMux
    port map (
            O => \N__13848\,
            I => \N__13823\
        );

    \I__1275\ : CEMux
    port map (
            O => \N__13847\,
            I => \N__13823\
        );

    \I__1274\ : CEMux
    port map (
            O => \N__13846\,
            I => \N__13823\
        );

    \I__1273\ : CEMux
    port map (
            O => \N__13845\,
            I => \N__13823\
        );

    \I__1272\ : CEMux
    port map (
            O => \N__13844\,
            I => \N__13823\
        );

    \I__1271\ : GlobalMux
    port map (
            O => \N__13823\,
            I => \N__13820\
        );

    \I__1270\ : gio2CtrlBuf
    port map (
            O => \N__13820\,
            I => \b2v_inst.N_305_1_g\
        );

    \I__1269\ : InMux
    port map (
            O => \N__13817\,
            I => \N__13814\
        );

    \I__1268\ : LocalMux
    port map (
            O => \N__13814\,
            I => \N__13811\
        );

    \I__1267\ : Odrv4
    port map (
            O => \N__13811\,
            I => \b2v_inst.N_4_i_i_a6_1\
        );

    \I__1266\ : InMux
    port map (
            O => \N__13808\,
            I => \N__13805\
        );

    \I__1265\ : LocalMux
    port map (
            O => \N__13805\,
            I => \N__13802\
        );

    \I__1264\ : Span4Mux_v
    port map (
            O => \N__13802\,
            I => \N__13798\
        );

    \I__1263\ : InMux
    port map (
            O => \N__13801\,
            I => \N__13795\
        );

    \I__1262\ : Sp12to4
    port map (
            O => \N__13798\,
            I => \N__13790\
        );

    \I__1261\ : LocalMux
    port map (
            O => \N__13795\,
            I => \N__13790\
        );

    \I__1260\ : Odrv12
    port map (
            O => \N__13790\,
            I => \b2v_inst4.pix_count_int_RNI0EPTZ0Z_0\
        );

    \I__1259\ : InMux
    port map (
            O => \N__13787\,
            I => \N__13784\
        );

    \I__1258\ : LocalMux
    port map (
            O => \N__13784\,
            I => \b2v_inst4.un1_pix_count_int_0_sqmuxa_10\
        );

    \I__1257\ : InMux
    port map (
            O => \N__13781\,
            I => \N__13778\
        );

    \I__1256\ : LocalMux
    port map (
            O => \N__13778\,
            I => \N__13775\
        );

    \I__1255\ : Span4Mux_v
    port map (
            O => \N__13775\,
            I => \N__13771\
        );

    \I__1254\ : InMux
    port map (
            O => \N__13774\,
            I => \N__13768\
        );

    \I__1253\ : Span4Mux_h
    port map (
            O => \N__13771\,
            I => \N__13763\
        );

    \I__1252\ : LocalMux
    port map (
            O => \N__13768\,
            I => \N__13763\
        );

    \I__1251\ : Odrv4
    port map (
            O => \N__13763\,
            I => \b2v_inst.cuenta_pixel_RNIT0FMZ0Z_1\
        );

    \I__1250\ : InMux
    port map (
            O => \N__13760\,
            I => \N__13755\
        );

    \I__1249\ : InMux
    port map (
            O => \N__13759\,
            I => \N__13752\
        );

    \I__1248\ : CascadeMux
    port map (
            O => \N__13758\,
            I => \N__13749\
        );

    \I__1247\ : LocalMux
    port map (
            O => \N__13755\,
            I => \N__13744\
        );

    \I__1246\ : LocalMux
    port map (
            O => \N__13752\,
            I => \N__13740\
        );

    \I__1245\ : InMux
    port map (
            O => \N__13749\,
            I => \N__13737\
        );

    \I__1244\ : InMux
    port map (
            O => \N__13748\,
            I => \N__13732\
        );

    \I__1243\ : InMux
    port map (
            O => \N__13747\,
            I => \N__13732\
        );

    \I__1242\ : Span4Mux_h
    port map (
            O => \N__13744\,
            I => \N__13729\
        );

    \I__1241\ : InMux
    port map (
            O => \N__13743\,
            I => \N__13726\
        );

    \I__1240\ : Span4Mux_h
    port map (
            O => \N__13740\,
            I => \N__13721\
        );

    \I__1239\ : LocalMux
    port map (
            O => \N__13737\,
            I => \N__13721\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__13732\,
            I => \b2v_inst.cuenta_pixelZ0Z_0\
        );

    \I__1237\ : Odrv4
    port map (
            O => \N__13729\,
            I => \b2v_inst.cuenta_pixelZ0Z_0\
        );

    \I__1236\ : LocalMux
    port map (
            O => \N__13726\,
            I => \b2v_inst.cuenta_pixelZ0Z_0\
        );

    \I__1235\ : Odrv4
    port map (
            O => \N__13721\,
            I => \b2v_inst.cuenta_pixelZ0Z_0\
        );

    \I__1234\ : CascadeMux
    port map (
            O => \N__13712\,
            I => \b2v_inst.cuenta_pixel_5_i_a2_0_2_5_cascade_\
        );

    \I__1233\ : InMux
    port map (
            O => \N__13709\,
            I => \N__13706\
        );

    \I__1232\ : LocalMux
    port map (
            O => \N__13706\,
            I => \N__13703\
        );

    \I__1231\ : Odrv4
    port map (
            O => \N__13703\,
            I => \b2v_inst.cuenta_pixelZ0Z_2\
        );

    \I__1230\ : InMux
    port map (
            O => \N__13700\,
            I => \N__13697\
        );

    \I__1229\ : LocalMux
    port map (
            O => \N__13697\,
            I => \N__13694\
        );

    \I__1228\ : Odrv4
    port map (
            O => \N__13694\,
            I => \b2v_inst.cuenta_pixelZ0Z_3\
        );

    \I__1227\ : InMux
    port map (
            O => \N__13691\,
            I => \N__13682\
        );

    \I__1226\ : InMux
    port map (
            O => \N__13690\,
            I => \N__13682\
        );

    \I__1225\ : InMux
    port map (
            O => \N__13689\,
            I => \N__13682\
        );

    \I__1224\ : LocalMux
    port map (
            O => \N__13682\,
            I => \N__13679\
        );

    \I__1223\ : Odrv4
    port map (
            O => \N__13679\,
            I => \b2v_inst.un1_cuenta_pixel_cry_1_c_RNI89THZ0\
        );

    \I__1222\ : CascadeMux
    port map (
            O => \N__13676\,
            I => \N__13672\
        );

    \I__1221\ : InMux
    port map (
            O => \N__13675\,
            I => \N__13664\
        );

    \I__1220\ : InMux
    port map (
            O => \N__13672\,
            I => \N__13664\
        );

    \I__1219\ : InMux
    port map (
            O => \N__13671\,
            I => \N__13664\
        );

    \I__1218\ : LocalMux
    port map (
            O => \N__13664\,
            I => \N__13661\
        );

    \I__1217\ : Odrv12
    port map (
            O => \N__13661\,
            I => \b2v_inst.un1_cuenta_pixel_cry_2_c_RNIACUHZ0\
        );

    \I__1216\ : InMux
    port map (
            O => \N__13658\,
            I => \N__13652\
        );

    \I__1215\ : InMux
    port map (
            O => \N__13657\,
            I => \N__13645\
        );

    \I__1214\ : InMux
    port map (
            O => \N__13656\,
            I => \N__13645\
        );

    \I__1213\ : InMux
    port map (
            O => \N__13655\,
            I => \N__13645\
        );

    \I__1212\ : LocalMux
    port map (
            O => \N__13652\,
            I => \N__13642\
        );

    \I__1211\ : LocalMux
    port map (
            O => \N__13645\,
            I => \N__13639\
        );

    \I__1210\ : Odrv4
    port map (
            O => \N__13642\,
            I => \b2v_inst.un1_cuenta_pixel_cry_4_c_RNIEI0IZ0\
        );

    \I__1209\ : Odrv4
    port map (
            O => \N__13639\,
            I => \b2v_inst.un1_cuenta_pixel_cry_4_c_RNIEI0IZ0\
        );

    \I__1208\ : InMux
    port map (
            O => \N__13634\,
            I => \N__13631\
        );

    \I__1207\ : LocalMux
    port map (
            O => \N__13631\,
            I => \N__13627\
        );

    \I__1206\ : InMux
    port map (
            O => \N__13630\,
            I => \N__13624\
        );

    \I__1205\ : Span4Mux_h
    port map (
            O => \N__13627\,
            I => \N__13621\
        );

    \I__1204\ : LocalMux
    port map (
            O => \N__13624\,
            I => \b2v_inst.cuenta_pixel_5_i_a2_0_2_5\
        );

    \I__1203\ : Odrv4
    port map (
            O => \N__13621\,
            I => \b2v_inst.cuenta_pixel_5_i_a2_0_2_5\
        );

    \I__1202\ : InMux
    port map (
            O => \N__13616\,
            I => \N__13613\
        );

    \I__1201\ : LocalMux
    port map (
            O => \N__13613\,
            I => \N__13609\
        );

    \I__1200\ : CascadeMux
    port map (
            O => \N__13612\,
            I => \N__13606\
        );

    \I__1199\ : Span4Mux_v
    port map (
            O => \N__13609\,
            I => \N__13602\
        );

    \I__1198\ : InMux
    port map (
            O => \N__13606\,
            I => \N__13597\
        );

    \I__1197\ : InMux
    port map (
            O => \N__13605\,
            I => \N__13597\
        );

    \I__1196\ : Odrv4
    port map (
            O => \N__13602\,
            I => \b2v_inst.cuenta_pixel_5_i_a2_0_1_5\
        );

    \I__1195\ : LocalMux
    port map (
            O => \N__13597\,
            I => \b2v_inst.cuenta_pixel_5_i_a2_0_1_5\
        );

    \I__1194\ : CascadeMux
    port map (
            O => \N__13592\,
            I => \N__13589\
        );

    \I__1193\ : InMux
    port map (
            O => \N__13589\,
            I => \N__13586\
        );

    \I__1192\ : LocalMux
    port map (
            O => \N__13586\,
            I => \N__13583\
        );

    \I__1191\ : Odrv4
    port map (
            O => \N__13583\,
            I => \b2v_inst.cuenta_pixelZ0Z_5\
        );

    \I__1190\ : InMux
    port map (
            O => \N__13580\,
            I => \N__13577\
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__13577\,
            I => \N__13574\
        );

    \I__1188\ : Odrv4
    port map (
            O => \N__13574\,
            I => \b2v_inst4.un1_pix_count_int_0_sqmuxa_7\
        );

    \I__1187\ : InMux
    port map (
            O => \N__13571\,
            I => \N__13568\
        );

    \I__1186\ : LocalMux
    port map (
            O => \N__13568\,
            I => \b2v_inst4.un1_pix_count_int_0_sqmuxa_13\
        );

    \I__1185\ : CascadeMux
    port map (
            O => \N__13565\,
            I => \b2v_inst4.un1_pix_count_int_0_sqmuxa_8_cascade_\
        );

    \I__1184\ : InMux
    port map (
            O => \N__13562\,
            I => \N__13559\
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__13559\,
            I => \b2v_inst4.un1_pix_count_int_0_sqmuxa_14\
        );

    \I__1182\ : InMux
    port map (
            O => \N__13556\,
            I => \N__13553\
        );

    \I__1181\ : LocalMux
    port map (
            O => \N__13553\,
            I => \N__13550\
        );

    \I__1180\ : Span4Mux_v
    port map (
            O => \N__13550\,
            I => \N__13547\
        );

    \I__1179\ : Odrv4
    port map (
            O => \N__13547\,
            I => \b2v_inst.pix_count_anteriorZ0Z_9\
        );

    \I__1178\ : CascadeMux
    port map (
            O => \N__13544\,
            I => \N__13541\
        );

    \I__1177\ : InMux
    port map (
            O => \N__13541\,
            I => \N__13538\
        );

    \I__1176\ : LocalMux
    port map (
            O => \N__13538\,
            I => \b2v_inst.un7_pix_count_int_0_I_51_c_RNOZ0\
        );

    \I__1175\ : CascadeMux
    port map (
            O => \N__13535\,
            I => \b2v_inst.N_1_0_0_cascade_\
        );

    \I__1174\ : CascadeMux
    port map (
            O => \N__13532\,
            I => \b2v_inst.N_4_i_i_o6_2_cascade_\
        );

    \I__1173\ : InMux
    port map (
            O => \N__13529\,
            I => \N__13526\
        );

    \I__1172\ : LocalMux
    port map (
            O => \N__13526\,
            I => \N__13523\
        );

    \I__1171\ : Span4Mux_h
    port map (
            O => \N__13523\,
            I => \N__13520\
        );

    \I__1170\ : Odrv4
    port map (
            O => \N__13520\,
            I => \b2v_inst.N_7\
        );

    \I__1169\ : CascadeMux
    port map (
            O => \N__13517\,
            I => \N__13514\
        );

    \I__1168\ : InMux
    port map (
            O => \N__13514\,
            I => \N__13511\
        );

    \I__1167\ : LocalMux
    port map (
            O => \N__13511\,
            I => \N__13508\
        );

    \I__1166\ : Odrv4
    port map (
            O => \N__13508\,
            I => \b2v_inst.un7_pix_count_int_0_I_21_c_RNOZ0\
        );

    \I__1165\ : InMux
    port map (
            O => \N__13505\,
            I => \N__13502\
        );

    \I__1164\ : LocalMux
    port map (
            O => \N__13502\,
            I => \b2v_inst.pix_count_anteriorZ0Z_6\
        );

    \I__1163\ : InMux
    port map (
            O => \N__13499\,
            I => \N__13496\
        );

    \I__1162\ : LocalMux
    port map (
            O => \N__13496\,
            I => \b2v_inst.pix_count_anteriorZ0Z_7\
        );

    \I__1161\ : CascadeMux
    port map (
            O => \N__13493\,
            I => \N__13490\
        );

    \I__1160\ : InMux
    port map (
            O => \N__13490\,
            I => \N__13487\
        );

    \I__1159\ : LocalMux
    port map (
            O => \N__13487\,
            I => \b2v_inst.pix_count_anteriorZ0Z_8\
        );

    \I__1158\ : InMux
    port map (
            O => \N__13484\,
            I => \b2v_inst.un1_cuenta_pixel_cry_3\
        );

    \I__1157\ : InMux
    port map (
            O => \N__13481\,
            I => \b2v_inst.un1_cuenta_pixel_cry_4\
        );

    \I__1156\ : InMux
    port map (
            O => \N__13478\,
            I => \N__13475\
        );

    \I__1155\ : LocalMux
    port map (
            O => \N__13475\,
            I => \N__13472\
        );

    \I__1154\ : Odrv4
    port map (
            O => \N__13472\,
            I => \b2v_inst.cuenta_pixelZ0Z_6\
        );

    \I__1153\ : InMux
    port map (
            O => \N__13469\,
            I => \N__13466\
        );

    \I__1152\ : LocalMux
    port map (
            O => \N__13466\,
            I => \N__13462\
        );

    \I__1151\ : InMux
    port map (
            O => \N__13465\,
            I => \N__13459\
        );

    \I__1150\ : Odrv4
    port map (
            O => \N__13462\,
            I => \b2v_inst.un1_cuenta_pixel_cry_5_c_RNIGL1IZ0\
        );

    \I__1149\ : LocalMux
    port map (
            O => \N__13459\,
            I => \b2v_inst.un1_cuenta_pixel_cry_5_c_RNIGL1IZ0\
        );

    \I__1148\ : InMux
    port map (
            O => \N__13454\,
            I => \b2v_inst.un1_cuenta_pixel_cry_5\
        );

    \I__1147\ : InMux
    port map (
            O => \N__13451\,
            I => \N__13448\
        );

    \I__1146\ : LocalMux
    port map (
            O => \N__13448\,
            I => \b2v_inst.cuenta_pixelZ0Z_7\
        );

    \I__1145\ : InMux
    port map (
            O => \N__13445\,
            I => \N__13441\
        );

    \I__1144\ : InMux
    port map (
            O => \N__13444\,
            I => \N__13438\
        );

    \I__1143\ : LocalMux
    port map (
            O => \N__13441\,
            I => \b2v_inst.un1_cuenta_pixel_cry_6_c_RNIIO2IZ0\
        );

    \I__1142\ : LocalMux
    port map (
            O => \N__13438\,
            I => \b2v_inst.un1_cuenta_pixel_cry_6_c_RNIIO2IZ0\
        );

    \I__1141\ : InMux
    port map (
            O => \N__13433\,
            I => \b2v_inst.un1_cuenta_pixel_cry_6\
        );

    \I__1140\ : InMux
    port map (
            O => \N__13430\,
            I => \N__13427\
        );

    \I__1139\ : LocalMux
    port map (
            O => \N__13427\,
            I => \b2v_inst.cuenta_pixelZ0Z_8\
        );

    \I__1138\ : InMux
    port map (
            O => \N__13424\,
            I => \b2v_inst.un1_cuenta_pixel_cry_7\
        );

    \I__1137\ : InMux
    port map (
            O => \N__13421\,
            I => \N__13418\
        );

    \I__1136\ : LocalMux
    port map (
            O => \N__13418\,
            I => \N__13415\
        );

    \I__1135\ : Odrv12
    port map (
            O => \N__13415\,
            I => \b2v_inst.cuenta_pixelZ0Z_9\
        );

    \I__1134\ : InMux
    port map (
            O => \N__13412\,
            I => \bfn_3_11_0_\
        );

    \I__1133\ : InMux
    port map (
            O => \N__13409\,
            I => \b2v_inst.un1_cuenta_pixel_cry_9\
        );

    \I__1132\ : InMux
    port map (
            O => \N__13406\,
            I => \N__13403\
        );

    \I__1131\ : LocalMux
    port map (
            O => \N__13403\,
            I => \b2v_inst.cuenta_pixelZ0Z_10\
        );

    \I__1130\ : CascadeMux
    port map (
            O => \N__13400\,
            I => \b2v_inst.un1_state_36_0_a2_0_2_1_cascade_\
        );

    \I__1129\ : InMux
    port map (
            O => \N__13397\,
            I => \N__13394\
        );

    \I__1128\ : LocalMux
    port map (
            O => \N__13394\,
            I => \N__13389\
        );

    \I__1127\ : InMux
    port map (
            O => \N__13393\,
            I => \N__13384\
        );

    \I__1126\ : InMux
    port map (
            O => \N__13392\,
            I => \N__13384\
        );

    \I__1125\ : Odrv4
    port map (
            O => \N__13389\,
            I => \b2v_inst.N_305_2\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__13384\,
            I => \b2v_inst.N_305_2\
        );

    \I__1123\ : CascadeMux
    port map (
            O => \N__13379\,
            I => \b2v_inst.N_305_2_cascade_\
        );

    \I__1122\ : InMux
    port map (
            O => \N__13376\,
            I => \N__13371\
        );

    \I__1121\ : InMux
    port map (
            O => \N__13375\,
            I => \N__13368\
        );

    \I__1120\ : InMux
    port map (
            O => \N__13374\,
            I => \N__13365\
        );

    \I__1119\ : LocalMux
    port map (
            O => \N__13371\,
            I => \N__13362\
        );

    \I__1118\ : LocalMux
    port map (
            O => \N__13368\,
            I => \b2v_inst.cuenta_pixelZ0Z_1\
        );

    \I__1117\ : LocalMux
    port map (
            O => \N__13365\,
            I => \b2v_inst.cuenta_pixelZ0Z_1\
        );

    \I__1116\ : Odrv4
    port map (
            O => \N__13362\,
            I => \b2v_inst.cuenta_pixelZ0Z_1\
        );

    \I__1115\ : InMux
    port map (
            O => \N__13355\,
            I => \b2v_inst.un1_cuenta_pixel_cry_1\
        );

    \I__1114\ : InMux
    port map (
            O => \N__13352\,
            I => \b2v_inst.un1_cuenta_pixel_cry_2\
        );

    \I__1113\ : InMux
    port map (
            O => \N__13349\,
            I => \N__13346\
        );

    \I__1112\ : LocalMux
    port map (
            O => \N__13346\,
            I => \b2v_inst.pix_count_anteriorZ0Z_13\
        );

    \I__1111\ : CascadeMux
    port map (
            O => \N__13343\,
            I => \N__13340\
        );

    \I__1110\ : InMux
    port map (
            O => \N__13340\,
            I => \N__13337\
        );

    \I__1109\ : LocalMux
    port map (
            O => \N__13337\,
            I => \N__13334\
        );

    \I__1108\ : Odrv4
    port map (
            O => \N__13334\,
            I => \b2v_inst.un7_pix_count_int_0_I_45_c_RNOZ0\
        );

    \I__1107\ : CascadeMux
    port map (
            O => \N__13331\,
            I => \N__13328\
        );

    \I__1106\ : InMux
    port map (
            O => \N__13328\,
            I => \N__13325\
        );

    \I__1105\ : LocalMux
    port map (
            O => \N__13325\,
            I => \b2v_inst.pix_count_anteriorZ0Z_14\
        );

    \I__1104\ : CascadeMux
    port map (
            O => \N__13322\,
            I => \b2v_inst4.un1_pix_count_int_0_sqmuxa_5_cascade_\
        );

    \I__1103\ : InMux
    port map (
            O => \N__13319\,
            I => \N__13316\
        );

    \I__1102\ : LocalMux
    port map (
            O => \N__13316\,
            I => \b2v_inst.pix_count_anteriorZ0Z_15\
        );

    \I__1101\ : CascadeMux
    port map (
            O => \N__13313\,
            I => \N__13310\
        );

    \I__1100\ : InMux
    port map (
            O => \N__13310\,
            I => \N__13307\
        );

    \I__1099\ : LocalMux
    port map (
            O => \N__13307\,
            I => \N__13304\
        );

    \I__1098\ : Odrv4
    port map (
            O => \N__13304\,
            I => \b2v_inst.pix_count_anteriorZ0Z_19\
        );

    \I__1097\ : CascadeMux
    port map (
            O => \N__13301\,
            I => \N__13298\
        );

    \I__1096\ : InMux
    port map (
            O => \N__13298\,
            I => \N__13295\
        );

    \I__1095\ : LocalMux
    port map (
            O => \N__13295\,
            I => \N__13292\
        );

    \I__1094\ : Span4Mux_h
    port map (
            O => \N__13292\,
            I => \N__13289\
        );

    \I__1093\ : Odrv4
    port map (
            O => \N__13289\,
            I => \b2v_inst.pix_count_anteriorZ0Z_16\
        );

    \I__1092\ : InMux
    port map (
            O => \N__13286\,
            I => \N__13283\
        );

    \I__1091\ : LocalMux
    port map (
            O => \N__13283\,
            I => \b2v_inst.pix_count_anteriorZ0Z_2\
        );

    \I__1090\ : CascadeMux
    port map (
            O => \N__13280\,
            I => \N__13277\
        );

    \I__1089\ : InMux
    port map (
            O => \N__13277\,
            I => \N__13274\
        );

    \I__1088\ : LocalMux
    port map (
            O => \N__13274\,
            I => \b2v_inst.pix_count_anteriorZ0Z_3\
        );

    \I__1087\ : InMux
    port map (
            O => \N__13271\,
            I => \N__13268\
        );

    \I__1086\ : LocalMux
    port map (
            O => \N__13268\,
            I => \b2v_inst.pix_count_anteriorZ0Z_0\
        );

    \I__1085\ : InMux
    port map (
            O => \N__13265\,
            I => \N__13262\
        );

    \I__1084\ : LocalMux
    port map (
            O => \N__13262\,
            I => \N__13259\
        );

    \I__1083\ : Odrv4
    port map (
            O => \N__13259\,
            I => \b2v_inst.pix_count_anteriorZ0Z_5\
        );

    \I__1082\ : CascadeMux
    port map (
            O => \N__13256\,
            I => \N__13253\
        );

    \I__1081\ : InMux
    port map (
            O => \N__13253\,
            I => \N__13250\
        );

    \I__1080\ : LocalMux
    port map (
            O => \N__13250\,
            I => \b2v_inst.un7_pix_count_int_0_I_33_c_RNOZ0\
        );

    \I__1079\ : InMux
    port map (
            O => \N__13247\,
            I => \N__13244\
        );

    \I__1078\ : LocalMux
    port map (
            O => \N__13244\,
            I => \b2v_inst.pix_count_anteriorZ0Z_18\
        );

    \I__1077\ : CascadeMux
    port map (
            O => \N__13241\,
            I => \N__13238\
        );

    \I__1076\ : InMux
    port map (
            O => \N__13238\,
            I => \N__13235\
        );

    \I__1075\ : LocalMux
    port map (
            O => \N__13235\,
            I => \N__13232\
        );

    \I__1074\ : Odrv4
    port map (
            O => \N__13232\,
            I => \b2v_inst.un7_pix_count_int_0_I_39_c_RNOZ0\
        );

    \I__1073\ : CascadeMux
    port map (
            O => \N__13229\,
            I => \N__13226\
        );

    \I__1072\ : InMux
    port map (
            O => \N__13226\,
            I => \N__13223\
        );

    \I__1071\ : LocalMux
    port map (
            O => \N__13223\,
            I => \b2v_inst.pix_count_anteriorZ0Z_12\
        );

    \I__1070\ : InMux
    port map (
            O => \N__13220\,
            I => \b2v_inst.un7_pix_count_int_0_N_2\
        );

    \I__1069\ : CascadeMux
    port map (
            O => \N__13217\,
            I => \N__13214\
        );

    \I__1068\ : InMux
    port map (
            O => \N__13214\,
            I => \N__13211\
        );

    \I__1067\ : LocalMux
    port map (
            O => \N__13211\,
            I => \b2v_inst.un7_pix_count_int_0_I_57_c_RNOZ0\
        );

    \I__1066\ : InMux
    port map (
            O => \N__13208\,
            I => \N__13205\
        );

    \I__1065\ : LocalMux
    port map (
            O => \N__13205\,
            I => \N__13202\
        );

    \I__1064\ : Span4Mux_h
    port map (
            O => \N__13202\,
            I => \N__13199\
        );

    \I__1063\ : Odrv4
    port map (
            O => \N__13199\,
            I => \b2v_inst4.un1_pix_count_int_0_sqmuxa_6\
        );

    \I__1062\ : CascadeMux
    port map (
            O => \N__13196\,
            I => \N__13193\
        );

    \I__1061\ : InMux
    port map (
            O => \N__13193\,
            I => \N__13190\
        );

    \I__1060\ : LocalMux
    port map (
            O => \N__13190\,
            I => \N__13187\
        );

    \I__1059\ : Odrv4
    port map (
            O => \N__13187\,
            I => \b2v_inst.un7_pix_count_int_0_I_27_c_RNOZ0\
        );

    \I__1058\ : InMux
    port map (
            O => \N__13184\,
            I => \N__13181\
        );

    \I__1057\ : LocalMux
    port map (
            O => \N__13181\,
            I => \b2v_inst.pix_count_anteriorZ0Z_4\
        );

    \I__1056\ : InMux
    port map (
            O => \N__13178\,
            I => \N__13175\
        );

    \I__1055\ : LocalMux
    port map (
            O => \N__13175\,
            I => \b2v_inst.un7_pix_count_int_0_I_1_c_RNOZ0\
        );

    \I__1054\ : CascadeMux
    port map (
            O => \N__13172\,
            I => \N__13169\
        );

    \I__1053\ : InMux
    port map (
            O => \N__13169\,
            I => \N__13166\
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__13166\,
            I => \b2v_inst.un7_pix_count_int_0_I_15_c_RNOZ0\
        );

    \I__1051\ : InMux
    port map (
            O => \N__13163\,
            I => \N__13156\
        );

    \I__1050\ : InMux
    port map (
            O => \N__13162\,
            I => \N__13156\
        );

    \I__1049\ : InMux
    port map (
            O => \N__13161\,
            I => \N__13153\
        );

    \I__1048\ : LocalMux
    port map (
            O => \N__13156\,
            I => b2v_inst4_pix_count_int_fast_0
        );

    \I__1047\ : LocalMux
    port map (
            O => \N__13153\,
            I => b2v_inst4_pix_count_int_fast_0
        );

    \I__1046\ : InMux
    port map (
            O => \N__13148\,
            I => \N__13145\
        );

    \I__1045\ : LocalMux
    port map (
            O => \N__13145\,
            I => \b2v_inst.N_13\
        );

    \I__1044\ : InMux
    port map (
            O => \N__13142\,
            I => \N__13133\
        );

    \I__1043\ : InMux
    port map (
            O => \N__13141\,
            I => \N__13133\
        );

    \I__1042\ : InMux
    port map (
            O => \N__13140\,
            I => \N__13133\
        );

    \I__1041\ : LocalMux
    port map (
            O => \N__13133\,
            I => b2v_inst4_pix_count_int_fast_2
        );

    \I__1040\ : CascadeMux
    port map (
            O => \N__13130\,
            I => \N__13126\
        );

    \I__1039\ : CascadeMux
    port map (
            O => \N__13129\,
            I => \N__13122\
        );

    \I__1038\ : InMux
    port map (
            O => \N__13126\,
            I => \N__13115\
        );

    \I__1037\ : InMux
    port map (
            O => \N__13125\,
            I => \N__13115\
        );

    \I__1036\ : InMux
    port map (
            O => \N__13122\,
            I => \N__13115\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__13115\,
            I => b2v_inst4_pix_count_int_fast_3
        );

    \I__1034\ : CascadeMux
    port map (
            O => \N__13112\,
            I => \N__13109\
        );

    \I__1033\ : InMux
    port map (
            O => \N__13109\,
            I => \N__13106\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__13106\,
            I => \N__13103\
        );

    \I__1031\ : Odrv4
    port map (
            O => \N__13103\,
            I => \b2v_inst.pix_count_anteriorZ0Z_1\
        );

    \I__1030\ : CascadeMux
    port map (
            O => \N__13100\,
            I => \b2v_inst.un4_pix_count_intlto6_d_1_1_cascade_\
        );

    \I__1029\ : InMux
    port map (
            O => \N__13097\,
            I => \N__13088\
        );

    \I__1028\ : InMux
    port map (
            O => \N__13096\,
            I => \N__13088\
        );

    \I__1027\ : InMux
    port map (
            O => \N__13095\,
            I => \N__13088\
        );

    \I__1026\ : LocalMux
    port map (
            O => \N__13088\,
            I => b2v_inst4_pix_count_int_fast_1
        );

    \I__1025\ : CascadeMux
    port map (
            O => \N__13085\,
            I => \b2v_inst.N_4_i_i_a3_0_0_cascade_\
        );

    \IN_MUX_bfv_17_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_13_0_\
        );

    \IN_MUX_bfv_9_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_5_0_\
        );

    \IN_MUX_bfv_9_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst.un8_dir_mem_2_cry_8\,
            carryinitout => \bfn_9_6_0_\
        );

    \IN_MUX_bfv_7_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_6_0_\
        );

    \IN_MUX_bfv_7_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst.un8_dir_mem_1_cry_7\,
            carryinitout => \bfn_7_7_0_\
        );

    \IN_MUX_bfv_2_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_11_0_\
        );

    \IN_MUX_bfv_2_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst.un7_pix_count_int_0_data_tmp_7\,
            carryinitout => \bfn_2_12_0_\
        );

    \IN_MUX_bfv_13_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_12_0_\
        );

    \IN_MUX_bfv_13_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst.un4_cuenta_cry_8\,
            carryinitout => \bfn_13_13_0_\
        );

    \IN_MUX_bfv_8_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_9_0_\
        );

    \IN_MUX_bfv_8_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst.un3_dir_mem_cry_7\,
            carryinitout => \bfn_8_10_0_\
        );

    \IN_MUX_bfv_6_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_5_0_\
        );

    \IN_MUX_bfv_6_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_6_0_\
        );

    \IN_MUX_bfv_6_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst.un1_indice_cry_8\,
            carryinitout => \bfn_6_7_0_\
        );

    \IN_MUX_bfv_3_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_10_0_\
        );

    \IN_MUX_bfv_3_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst.un1_cuenta_pixel_cry_8\,
            carryinitout => \bfn_3_11_0_\
        );

    \IN_MUX_bfv_19_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_19_14_0_\
        );

    \IN_MUX_bfv_17_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_8_0_\
        );

    \IN_MUX_bfv_17_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst.valor_max_final4_3_cry_7\,
            carryinitout => \bfn_17_9_0_\
        );

    \IN_MUX_bfv_17_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_5_0_\
        );

    \IN_MUX_bfv_17_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst.valor_max_final4_2_cry_7\,
            carryinitout => \bfn_17_6_0_\
        );

    \IN_MUX_bfv_18_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_6_0_\
        );

    \IN_MUX_bfv_18_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst.un2_valor_max2_cry_7\,
            carryinitout => \bfn_18_7_0_\
        );

    \IN_MUX_bfv_13_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_16_0_\
        );

    \IN_MUX_bfv_13_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst.dir_energia_cry_7\,
            carryinitout => \bfn_13_17_0_\
        );

    \IN_MUX_bfv_15_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_8_0_\
        );

    \IN_MUX_bfv_15_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst.data_a_escribir11_7\,
            carryinitout => \bfn_15_9_0_\
        );

    \IN_MUX_bfv_17_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_16_0_\
        );

    \IN_MUX_bfv_5_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_13_0_\
        );

    \IN_MUX_bfv_5_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst4.un1_pix_count_int_cry_7\,
            carryinitout => \bfn_5_14_0_\
        );

    \IN_MUX_bfv_5_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst4.un1_pix_count_int_cry_15\,
            carryinitout => \bfn_5_15_0_\
        );

    \IN_MUX_bfv_14_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_14_0_\
        );

    \IN_MUX_bfv_14_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst.un14_data_ram_energia_o_cry_7\,
            carryinitout => \bfn_14_15_0_\
        );

    \IN_MUX_bfv_13_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_6_0_\
        );

    \IN_MUX_bfv_13_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst.un2_dir_mem_2_cry_7\,
            carryinitout => \bfn_13_7_0_\
        );

    \IN_MUX_bfv_8_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_5_0_\
        );

    \IN_MUX_bfv_8_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst.un2_dir_mem_1_cry_7\,
            carryinitout => \bfn_8_6_0_\
        );

    \IN_MUX_bfv_15_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_10_0_\
        );

    \IN_MUX_bfv_15_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst.eventos_cry_7\,
            carryinitout => \bfn_15_11_0_\
        );

    \IN_MUX_bfv_17_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_10_0_\
        );

    \IN_MUX_bfv_17_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst.valor_max_final4_1_cry_7\,
            carryinitout => \bfn_17_11_0_\
        );

    \IN_MUX_bfv_18_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_8_0_\
        );

    \IN_MUX_bfv_18_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst.valor_max_final4_0_cry_7\,
            carryinitout => \bfn_18_9_0_\
        );

    \IN_MUX_bfv_16_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_6_0_\
        );

    \IN_MUX_bfv_16_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst.un2_valor_max1_cry_7\,
            carryinitout => \bfn_16_7_0_\
        );

    \b2v_inst.state_RNI9A7V8_0_29\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__14927\,
            GLOBALBUFFEROUTPUT => \b2v_inst.N_305_1_g\
        );

    \reset_ibuf_RNI8255_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__24088\,
            GLOBALBUFFEROUTPUT => reset_c_i_g
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \reset_ibuf_RNI8255_LC_1_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27787\,
            lcout => reset_c_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un4_pix_count_intlto6_1_x1_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__16747\,
            in1 => \N__15018\,
            in2 => \N__16852\,
            in3 => \N__15043\,
            lcout => \b2v_inst.un4_pix_count_intlto6_1_xZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNO_27_29_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__15019\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15042\,
            lcout => OPEN,
            ltout => \b2v_inst.N_4_i_i_a3_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNO_19_29_LC_1_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011101100"
        )
    port map (
            in0 => \N__16748\,
            in1 => \N__16847\,
            in2 => \N__13085\,
            in3 => \N__13148\,
            lcout => \b2v_inst.N_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un4_pix_count_intlto6_1_x0_LC_1_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110111"
        )
    port map (
            in0 => \N__15017\,
            in1 => \N__15041\,
            in2 => \_gnd_net_\,
            in3 => \N__16843\,
            lcout => \b2v_inst.un4_pix_count_intlto6_1_xZ0Z0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst4.pix_count_int_fast_5_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__14786\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13970\,
            lcout => b2v_inst4_pix_count_int_fast_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34509\,
            ce => 'H',
            sr => \N__38041\
        );

    \b2v_inst4.pix_count_int_fast_6_LC_1_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14784\,
            in2 => \_gnd_net_\,
            in3 => \N__13952\,
            lcout => b2v_inst4_pix_count_int_fast_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34509\,
            ce => 'H',
            sr => \N__38041\
        );

    \b2v_inst4.pix_count_int_5_LC_1_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__14785\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13969\,
            lcout => \SYNTHESIZED_WIRE_4_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34509\,
            ce => 'H',
            sr => \N__38041\
        );

    \b2v_inst.un7_pix_count_int_0_I_15_c_RNO_LC_1_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__13265\,
            in1 => \N__16746\,
            in2 => \N__15807\,
            in3 => \N__13184\,
            lcout => \b2v_inst.un7_pix_count_int_0_I_15_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.g0_3_LC_1_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111101111111"
        )
    port map (
            in0 => \N__13142\,
            in1 => \N__13097\,
            in2 => \N__13130\,
            in3 => \N__13163\,
            lcout => OPEN,
            ltout => \b2v_inst.un4_pix_count_intlto6_d_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.g2_1_LC_1_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111110111"
        )
    port map (
            in0 => \N__15878\,
            in1 => \N__15801\,
            in2 => \N__13100\,
            in3 => \N__16756\,
            lcout => \b2v_inst.g2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un4_pix_count_intlto6_d_1_LC_1_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111101111111"
        )
    port map (
            in0 => \N__13140\,
            in1 => \N__13096\,
            in2 => \N__13129\,
            in3 => \N__13162\,
            lcout => \b2v_inst.un4_pix_count_intlto6_dZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst4.pix_count_int_fast_1_LC_1_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14036\,
            lcout => b2v_inst4_pix_count_int_fast_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34514\,
            ce => 'H',
            sr => \N__38042\
        );

    \b2v_inst.un7_pix_count_int_0_I_1_c_RNO_LC_1_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__13161\,
            in1 => \N__13095\,
            in2 => \N__13112\,
            in3 => \N__13271\,
            lcout => \b2v_inst.un7_pix_count_int_0_I_1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst4.pix_count_int_fast_0_LC_1_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13808\,
            in2 => \_gnd_net_\,
            in3 => \N__14791\,
            lcout => b2v_inst4_pix_count_int_fast_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34514\,
            ce => 'H',
            sr => \N__38042\
        );

    \b2v_inst.state_RNO_28_29_LC_1_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000000000"
        )
    port map (
            in0 => \N__15273\,
            in1 => \N__13141\,
            in2 => \N__15199\,
            in3 => \N__13125\,
            lcout => \b2v_inst.N_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst4.pix_count_int_fast_2_LC_1_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__14778\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14012\,
            lcout => b2v_inst4_pix_count_int_fast_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34523\,
            ce => 'H',
            sr => \N__38043\
        );

    \b2v_inst4.pix_count_int_0_LC_1_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13801\,
            in2 => \_gnd_net_\,
            in3 => \N__14783\,
            lcout => \SYNTHESIZED_WIRE_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34523\,
            ce => 'H',
            sr => \N__38043\
        );

    \b2v_inst4.pix_count_int_fast_3_LC_1_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101000001010"
        )
    port map (
            in0 => \N__13988\,
            in1 => \_gnd_net_\,
            in2 => \N__14792\,
            in3 => \_gnd_net_\,
            lcout => b2v_inst4_pix_count_int_fast_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34523\,
            ce => 'H',
            sr => \N__38043\
        );

    \b2v_inst4.pix_count_int_3_LC_1_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14779\,
            in2 => \_gnd_net_\,
            in3 => \N__13987\,
            lcout => \SYNTHESIZED_WIRE_4_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34523\,
            ce => 'H',
            sr => \N__38043\
        );

    \b2v_inst4.pix_count_int_fast_11_LC_1_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__14777\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14687\,
            lcout => b2v_inst4_pix_count_int_fast_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34523\,
            ce => 'H',
            sr => \N__38043\
        );

    \b2v_inst4.state_RNI8N511_0_LC_1_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__14897\,
            in1 => \N__15503\,
            in2 => \_gnd_net_\,
            in3 => \N__15875\,
            lcout => \b2v_inst4.un1_pix_count_int_0_sqmuxa_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.pix_count_anterior_1_LC_2_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15193\,
            lcout => \b2v_inst.pix_count_anteriorZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34511\,
            ce => \N__13845\,
            sr => \N__38040\
        );

    \b2v_inst.pix_count_anterior_4_LC_2_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16757\,
            lcout => \b2v_inst.pix_count_anteriorZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34511\,
            ce => \N__13845\,
            sr => \N__38040\
        );

    \b2v_inst.pix_count_anterior_9_LC_2_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15566\,
            lcout => \b2v_inst.pix_count_anteriorZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34511\,
            ce => \N__13845\,
            sr => \N__38040\
        );

    \b2v_inst.cuenta_pixel_7_LC_2_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13445\,
            lcout => \b2v_inst.cuenta_pixelZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34511\,
            ce => \N__13845\,
            sr => \N__38040\
        );

    \b2v_inst.cuenta_pixel_8_LC_2_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__13397\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14583\,
            lcout => \b2v_inst.cuenta_pixelZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34511\,
            ce => \N__13845\,
            sr => \N__38040\
        );

    \b2v_inst.un7_pix_count_int_0_I_1_c_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13178\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_11_0_\,
            carryout => \b2v_inst.un7_pix_count_int_0_data_tmp_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un7_pix_count_int_0_I_27_c_LC_2_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37300\,
            in2 => \N__13196\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.un7_pix_count_int_0_data_tmp_0\,
            carryout => \b2v_inst.un7_pix_count_int_0_data_tmp_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un7_pix_count_int_0_I_15_c_LC_2_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37296\,
            in2 => \N__13172\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.un7_pix_count_int_0_data_tmp_1\,
            carryout => \b2v_inst.un7_pix_count_int_0_data_tmp_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un7_pix_count_int_0_I_21_c_LC_2_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37299\,
            in2 => \N__13517\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.un7_pix_count_int_0_data_tmp_2\,
            carryout => \b2v_inst.un7_pix_count_int_0_data_tmp_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un7_pix_count_int_0_I_51_c_LC_2_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37298\,
            in2 => \N__13544\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.un7_pix_count_int_0_data_tmp_3\,
            carryout => \b2v_inst.un7_pix_count_int_0_data_tmp_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un7_pix_count_int_0_I_9_c_LC_2_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37302\,
            in2 => \N__13889\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.un7_pix_count_int_0_data_tmp_4\,
            carryout => \b2v_inst.un7_pix_count_int_0_data_tmp_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un7_pix_count_int_0_I_39_c_LC_2_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37297\,
            in2 => \N__13241\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.un7_pix_count_int_0_data_tmp_5\,
            carryout => \b2v_inst.un7_pix_count_int_0_data_tmp_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un7_pix_count_int_0_I_45_c_LC_2_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37301\,
            in2 => \N__13343\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.un7_pix_count_int_0_data_tmp_6\,
            carryout => \b2v_inst.un7_pix_count_int_0_data_tmp_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un7_pix_count_int_0_I_57_c_LC_2_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37265\,
            in2 => \N__13217\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_12_0_\,
            carryout => \b2v_inst.un7_pix_count_int_0_data_tmp_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un7_pix_count_int_0_I_33_c_LC_2_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37264\,
            in2 => \N__13256\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.un7_pix_count_int_0_data_tmp_8\,
            carryout => \b2v_inst.un7_pix_count_int_0_N_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un7_pix_count_int_0_N_2_THRU_LUT4_0_LC_2_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13220\,
            lcout => \b2v_inst.un7_pix_count_int_0_N_2_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un7_pix_count_int_0_I_57_c_RNO_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__17610\,
            in1 => \N__17445\,
            in2 => \N__13301\,
            in3 => \N__13862\,
            lcout => \b2v_inst.un7_pix_count_int_0_I_57_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.g0_5_LC_2_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011111111111"
        )
    port map (
            in0 => \N__15262\,
            in1 => \N__15226\,
            in2 => \N__15198\,
            in3 => \N__15132\,
            lcout => \b2v_inst.un4_pix_count_intlto6_d_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst4.state_RNI9BF02_0_LC_2_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__13208\,
            in1 => \N__14876\,
            in2 => \_gnd_net_\,
            in3 => \N__15641\,
            lcout => \b2v_inst4.un1_pix_count_int_0_sqmuxa_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un7_pix_count_int_0_I_27_c_RNO_LC_2_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__15225\,
            in1 => \N__13286\,
            in2 => \N__13280\,
            in3 => \N__15121\,
            lcout => \b2v_inst.un7_pix_count_int_0_I_27_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.pix_count_anterior_2_LC_2_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__15123\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst.pix_count_anteriorZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34515\,
            ce => \N__13846\,
            sr => \N__38046\
        );

    \b2v_inst.pix_count_anterior_3_LC_2_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15236\,
            lcout => \b2v_inst.pix_count_anteriorZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34515\,
            ce => \N__13846\,
            sr => \N__38046\
        );

    \b2v_inst4.pix_count_int_RNIQK3K1_0_LC_2_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__15122\,
            in1 => \N__15271\,
            in2 => \N__15239\,
            in3 => \N__15824\,
            lcout => \b2v_inst4.un1_pix_count_int_0_sqmuxa_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.pix_count_anterior_0_LC_2_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__15272\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst.pix_count_anteriorZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34515\,
            ce => \N__13846\,
            sr => \N__38046\
        );

    \b2v_inst.pix_count_anterior_5_LC_2_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15825\,
            lcout => \b2v_inst.pix_count_anteriorZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34515\,
            ce => \N__13846\,
            sr => \N__38046\
        );

    \b2v_inst.un7_pix_count_int_0_I_33_c_RNO_LC_2_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__17500\,
            in1 => \N__17722\,
            in2 => \N__13313\,
            in3 => \N__13247\,
            lcout => \b2v_inst.un7_pix_count_int_0_I_33_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.pix_count_anterior_18_LC_2_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17501\,
            lcout => \b2v_inst.pix_count_anteriorZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34515\,
            ce => \N__13846\,
            sr => \N__38046\
        );

    \b2v_inst.un7_pix_count_int_0_I_39_c_RNO_LC_2_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__15376\,
            in1 => \N__16474\,
            in2 => \N__13229\,
            in3 => \N__13349\,
            lcout => \b2v_inst.un7_pix_count_int_0_I_39_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.pix_count_anterior_12_LC_2_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15377\,
            lcout => \b2v_inst.pix_count_anteriorZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34524\,
            ce => \N__13848\,
            sr => \N__38049\
        );

    \b2v_inst.pix_count_anterior_13_LC_2_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16475\,
            lcout => \b2v_inst.pix_count_anteriorZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34524\,
            ce => \N__13848\,
            sr => \N__38049\
        );

    \b2v_inst.un7_pix_count_int_0_I_45_c_RNO_LC_2_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__16408\,
            in1 => \N__16338\,
            in2 => \N__13331\,
            in3 => \N__13319\,
            lcout => \b2v_inst.un7_pix_count_int_0_I_45_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.pix_count_anterior_14_LC_2_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__16340\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst.pix_count_anteriorZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34524\,
            ce => \N__13848\,
            sr => \N__38049\
        );

    \b2v_inst4.pix_count_int_RNIDQ1Q_1_LC_2_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15171\,
            in2 => \_gnd_net_\,
            in3 => \N__16752\,
            lcout => OPEN,
            ltout => \b2v_inst4.un1_pix_count_int_0_sqmuxa_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst4.pix_count_int_RNII16D3_14_LC_2_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__16339\,
            in1 => \N__16409\,
            in2 => \N__13322\,
            in3 => \N__13787\,
            lcout => \b2v_inst4.un1_pix_count_int_0_sqmuxa_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.pix_count_anterior_15_LC_2_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__16410\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst.pix_count_anteriorZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34524\,
            ce => \N__13848\,
            sr => \N__38049\
        );

    \b2v_inst.pix_count_anterior_19_LC_2_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17705\,
            lcout => \b2v_inst.pix_count_anteriorZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34525\,
            ce => \N__13850\,
            sr => \N__38053\
        );

    \b2v_inst.pix_count_anterior_16_LC_2_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17612\,
            lcout => \b2v_inst.pix_count_anteriorZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34525\,
            ce => \N__13850\,
            sr => \N__38053\
        );

    \b2v_inst.cuenta_pixel_9_LC_3_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__13393\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14641\,
            lcout => \b2v_inst.cuenta_pixelZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34516\,
            ce => \N__13851\,
            sr => \N__38047\
        );

    \b2v_inst.cuenta_pixel_0_LC_3_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13392\,
            in2 => \_gnd_net_\,
            in3 => \N__13747\,
            lcout => \b2v_inst.cuenta_pixelZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34516\,
            ce => \N__13851\,
            sr => \N__38047\
        );

    \b2v_inst.cuenta_pixel_RNINOUV1_10_LC_3_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__14640\,
            in1 => \N__14617\,
            in2 => \N__14590\,
            in3 => \N__13658\,
            lcout => OPEN,
            ltout => \b2v_inst.un1_state_36_0_a2_0_2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.cuenta_pixel_RNIISKR5_0_LC_3_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__13634\,
            in1 => \N__13616\,
            in2 => \N__13400\,
            in3 => \N__14557\,
            lcout => \b2v_inst.N_305_2\,
            ltout => \b2v_inst.N_305_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.cuenta_pixel_6_LC_3_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13469\,
            in2 => \N__13379\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst.cuenta_pixelZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34516\,
            ce => \N__13851\,
            sr => \N__38047\
        );

    \b2v_inst.cuenta_pixel_1_LC_3_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__13748\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13375\,
            lcout => \b2v_inst.cuenta_pixelZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34516\,
            ce => \N__13851\,
            sr => \N__38047\
        );

    \b2v_inst.cuenta_pixel_RNIT0FM_1_LC_3_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13743\,
            in2 => \_gnd_net_\,
            in3 => \N__13374\,
            lcout => \b2v_inst.cuenta_pixel_RNIT0FMZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un1_cuenta_pixel_cry_5_c_RNI2E441_LC_3_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__13444\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13465\,
            lcout => \b2v_inst.cuenta_pixel_5_i_a2_1_1_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un1_cuenta_pixel_cry_1_c_LC_3_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13376\,
            in2 => \N__13758\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_3_10_0_\,
            carryout => \b2v_inst.un1_cuenta_pixel_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un1_cuenta_pixel_cry_1_c_RNI89TH_LC_3_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13709\,
            in2 => \_gnd_net_\,
            in3 => \N__13355\,
            lcout => \b2v_inst.un1_cuenta_pixel_cry_1_c_RNI89THZ0\,
            ltout => OPEN,
            carryin => \b2v_inst.un1_cuenta_pixel_cry_1\,
            carryout => \b2v_inst.un1_cuenta_pixel_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un1_cuenta_pixel_cry_2_c_RNIACUH_LC_3_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13700\,
            in2 => \_gnd_net_\,
            in3 => \N__13352\,
            lcout => \b2v_inst.un1_cuenta_pixel_cry_2_c_RNIACUHZ0\,
            ltout => OPEN,
            carryin => \b2v_inst.un1_cuenta_pixel_cry_2\,
            carryout => \b2v_inst.un1_cuenta_pixel_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un1_cuenta_pixel_cry_3_c_RNICFVH_LC_3_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13901\,
            in3 => \N__13484\,
            lcout => \b2v_inst.un1_cuenta_pixel_cry_3_c_RNICFVHZ0\,
            ltout => OPEN,
            carryin => \b2v_inst.un1_cuenta_pixel_cry_3\,
            carryout => \b2v_inst.un1_cuenta_pixel_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un1_cuenta_pixel_cry_4_c_RNIEI0I_LC_3_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13592\,
            in3 => \N__13481\,
            lcout => \b2v_inst.un1_cuenta_pixel_cry_4_c_RNIEI0IZ0\,
            ltout => OPEN,
            carryin => \b2v_inst.un1_cuenta_pixel_cry_4\,
            carryout => \b2v_inst.un1_cuenta_pixel_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un1_cuenta_pixel_cry_5_c_RNIGL1I_LC_3_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13478\,
            in2 => \_gnd_net_\,
            in3 => \N__13454\,
            lcout => \b2v_inst.un1_cuenta_pixel_cry_5_c_RNIGL1IZ0\,
            ltout => OPEN,
            carryin => \b2v_inst.un1_cuenta_pixel_cry_5\,
            carryout => \b2v_inst.un1_cuenta_pixel_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un1_cuenta_pixel_cry_6_c_RNIIO2I_LC_3_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13451\,
            in2 => \_gnd_net_\,
            in3 => \N__13433\,
            lcout => \b2v_inst.un1_cuenta_pixel_cry_6_c_RNIIO2IZ0\,
            ltout => OPEN,
            carryin => \b2v_inst.un1_cuenta_pixel_cry_6\,
            carryout => \b2v_inst.un1_cuenta_pixel_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un1_cuenta_pixel_cry_7_c_RNIKR3I_LC_3_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13430\,
            in2 => \_gnd_net_\,
            in3 => \N__13424\,
            lcout => \b2v_inst.un1_cuenta_pixel_cry_7_c_RNIKR3IZ0\,
            ltout => OPEN,
            carryin => \b2v_inst.un1_cuenta_pixel_cry_7\,
            carryout => \b2v_inst.un1_cuenta_pixel_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un1_cuenta_pixel_cry_8_c_RNIMU4I_LC_3_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13421\,
            in2 => \_gnd_net_\,
            in3 => \N__13412\,
            lcout => \b2v_inst.un1_cuenta_pixel_cry_8_c_RNIMU4IZ0\,
            ltout => OPEN,
            carryin => \bfn_3_11_0_\,
            carryout => \b2v_inst.un1_cuenta_pixel_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.cuenta_pixel_RNIVBL9_10_LC_3_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13406\,
            in2 => \_gnd_net_\,
            in3 => \N__13409\,
            lcout => \b2v_inst.cuenta_pixel_RNIVBL9Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.cuenta_pixel_10_LC_3_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14616\,
            lcout => \b2v_inst.cuenta_pixelZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34497\,
            ce => \N__13844\,
            sr => \N__38044\
        );

    \b2v_inst4.pix_count_int_9_rep1_LC_3_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14816\,
            lcout => \SYNTHESIZED_WIRE_4_9_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34503\,
            ce => 'H',
            sr => \N__38048\
        );

    \b2v_inst.un7_pix_count_int_0_I_51_c_RNO_LC_3_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__13556\,
            in1 => \N__15495\,
            in2 => \N__13493\,
            in3 => \N__15305\,
            lcout => \b2v_inst.un7_pix_count_int_0_I_51_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNO_26_29_LC_3_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000000000"
        )
    port map (
            in0 => \N__15306\,
            in1 => \N__15725\,
            in2 => \N__15779\,
            in3 => \N__15674\,
            lcout => OPEN,
            ltout => \b2v_inst.N_1_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNO_18_29_LC_3_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__16429\,
            in1 => \N__16362\,
            in2 => \N__13535\,
            in3 => \N__16499\,
            lcout => OPEN,
            ltout => \b2v_inst.N_4_i_i_o6_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNO_7_29_LC_3_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001010100000"
        )
    port map (
            in0 => \N__13817\,
            in1 => \N__16271\,
            in2 => \N__13532\,
            in3 => \N__13529\,
            lcout => \b2v_inst.N_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un7_pix_count_int_0_I_21_c_RNO_LC_3_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__13505\,
            in1 => \N__16822\,
            in2 => \N__15859\,
            in3 => \N__13499\,
            lcout => \b2v_inst.un7_pix_count_int_0_I_21_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.pix_count_anterior_6_LC_3_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15848\,
            lcout => \b2v_inst.pix_count_anteriorZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34512\,
            ce => \N__13849\,
            sr => \N__38050\
        );

    \b2v_inst.pix_count_anterior_7_LC_3_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16824\,
            lcout => \b2v_inst.pix_count_anteriorZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34512\,
            ce => \N__13849\,
            sr => \N__38050\
        );

    \b2v_inst.pix_count_anterior_8_LC_3_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15502\,
            lcout => \b2v_inst.pix_count_anteriorZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34512\,
            ce => \N__13849\,
            sr => \N__38050\
        );

    \b2v_inst4.pix_count_int_RNI5JOL1_9_LC_3_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__16823\,
            in1 => \N__16500\,
            in2 => \N__15565\,
            in3 => \N__15617\,
            lcout => OPEN,
            ltout => \b2v_inst4.un1_pix_count_int_0_sqmuxa_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst4.pix_count_int_RNIQKHN8_0_LC_3_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__13580\,
            in1 => \N__13571\,
            in2 => \N__13565\,
            in3 => \N__13562\,
            lcout => \b2v_inst4.un1_pix_count_int_0_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst4.pix_count_int_12_LC_3_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__14752\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14068\,
            lcout => \SYNTHESIZED_WIRE_4_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34517\,
            ce => 'H',
            sr => \N__38054\
        );

    \b2v_inst4.pix_count_int_fast_12_LC_3_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__14069\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14753\,
            lcout => b2v_inst4_pix_count_int_fast_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34517\,
            ce => 'H',
            sr => \N__38054\
        );

    \b2v_inst4.pix_count_int_2_LC_3_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__14754\,
            in1 => \N__14008\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \SYNTHESIZED_WIRE_4_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34517\,
            ce => 'H',
            sr => \N__38054\
        );

    \b2v_inst4.pix_count_int_6_LC_3_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14751\,
            in2 => \_gnd_net_\,
            in3 => \N__13948\,
            lcout => \SYNTHESIZED_WIRE_4_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34517\,
            ce => 'H',
            sr => \N__38054\
        );

    \b2v_inst.state_19_LC_3_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30977\,
            lcout => \b2v_inst.stateZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34517\,
            ce => 'H',
            sr => \N__38054\
        );

    \b2v_inst.state_32_rep1_LC_3_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21269\,
            lcout => \b2v_inst.state_32_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34517\,
            ce => 'H',
            sr => \N__38054\
        );

    \b2v_inst4.state_0_LC_3_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14895\,
            in2 => \_gnd_net_\,
            in3 => \N__14875\,
            lcout => \b2v_inst4.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34517\,
            ce => 'H',
            sr => \N__38054\
        );

    \b2v_inst4.pix_count_int_1_LC_3_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14032\,
            lcout => \SYNTHESIZED_WIRE_4_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34517\,
            ce => 'H',
            sr => \N__38054\
        );

    \b2v_inst4.pix_count_int_RNIIJDN1_17_LC_3_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__17490\,
            in1 => \N__17594\,
            in2 => \N__17723\,
            in3 => \N__17444\,
            lcout => \b2v_inst4.un1_pix_count_int_0_sqmuxa_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.ignorar_ancho_1_RNO_1_LC_5_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13774\,
            in2 => \_gnd_net_\,
            in3 => \N__13760\,
            lcout => \b2v_inst.ignorar_ancho_1_RNOZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.cuenta_pixel_RNI70MJ1_0_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__13781\,
            in1 => \_gnd_net_\,
            in2 => \N__13919\,
            in3 => \N__13759\,
            lcout => \b2v_inst.cuenta_pixel_5_i_a2_0_2_5\,
            ltout => \b2v_inst.cuenta_pixel_5_i_a2_0_2_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.ignorar_anterior_RNO_1_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__28205\,
            in1 => \N__13605\,
            in2 => \N__13712\,
            in3 => \N__13656\,
            lcout => \b2v_inst.un1_state_36_0_sn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un1_cuenta_pixel_cry_1_c_RNIILR31_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13689\,
            in2 => \_gnd_net_\,
            in3 => \N__13671\,
            lcout => \b2v_inst.cuenta_pixel_5_i_a2_0_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.cuenta_pixel_2_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__13691\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst.cuenta_pixelZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34495\,
            ce => \N__13852\,
            sr => \N__38045\
        );

    \b2v_inst.cuenta_pixel_3_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13675\,
            lcout => \b2v_inst.cuenta_pixelZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34495\,
            ce => \N__13852\,
            sr => \N__38045\
        );

    \b2v_inst.ignorar_ancho_1_RNO_2_LC_5_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__13690\,
            in1 => \N__13914\,
            in2 => \N__13676\,
            in3 => \N__13655\,
            lcout => \b2v_inst.ignorar_ancho_1_RNOZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.cuenta_pixel_5_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010101010101010"
        )
    port map (
            in0 => \N__13657\,
            in1 => \N__13630\,
            in2 => \N__13612\,
            in3 => \N__14543\,
            lcout => \b2v_inst.cuenta_pixelZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34495\,
            ce => \N__13852\,
            sr => \N__38045\
        );

    \b2v_inst.cuenta_pixel_4_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13918\,
            lcout => \b2v_inst.cuenta_pixelZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34495\,
            ce => \N__13852\,
            sr => \N__38045\
        );

    \b2v_inst.un7_pix_count_int_0_I_9_c_RNO_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__15596\,
            in1 => \N__15342\,
            in2 => \N__13871\,
            in3 => \N__13877\,
            lcout => \b2v_inst.un7_pix_count_int_0_I_9_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.pix_count_anterior_10_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15597\,
            lcout => \b2v_inst.pix_count_anteriorZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34477\,
            ce => \N__13847\,
            sr => \N__38051\
        );

    \b2v_inst.pix_count_anterior_11_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15343\,
            lcout => \b2v_inst.pix_count_anteriorZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34477\,
            ce => \N__13847\,
            sr => \N__38051\
        );

    \b2v_inst1.r_Clk_Count_RNIGMPV1_0_2_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__22634\,
            in1 => \N__22893\,
            in2 => \N__16913\,
            in3 => \N__16541\,
            lcout => \b2v_inst1.r_RX_Byte_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.pix_count_anterior_17_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__17437\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst.pix_count_anteriorZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34496\,
            ce => \N__13853\,
            sr => \N__38055\
        );

    \b2v_inst.state_RNO_17_29_LC_5_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__28202\,
            in1 => \N__17713\,
            in2 => \_gnd_net_\,
            in3 => \N__17592\,
            lcout => \b2v_inst.N_4_i_i_a6_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.ignorar_anterior_RNO_0_LC_5_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__28203\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26004\,
            lcout => \b2v_inst.un1_state_36_0_rn_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst4.pix_count_int_RNI0EPT_0_LC_5_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15281\,
            in2 => \N__28760\,
            in3 => \N__28751\,
            lcout => \b2v_inst4.pix_count_int_RNI0EPTZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_5_13_0_\,
            carryout => \b2v_inst4.un1_pix_count_int_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst4.un1_pix_count_int_cry_0_c_RNIIC2I_LC_5_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15197\,
            in2 => \_gnd_net_\,
            in3 => \N__14015\,
            lcout => \b2v_inst4.un1_pix_count_int_cry_0_c_RNIIC2IZ0\,
            ltout => OPEN,
            carryin => \b2v_inst4.un1_pix_count_int_cry_0\,
            carryout => \b2v_inst4.un1_pix_count_int_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst4.un1_pix_count_int_cry_1_c_RNIKF3I_LC_5_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15140\,
            in2 => \_gnd_net_\,
            in3 => \N__13991\,
            lcout => \b2v_inst4.un1_pix_count_int_cry_1_c_RNIKF3IZ0\,
            ltout => OPEN,
            carryin => \b2v_inst4.un1_pix_count_int_cry_1\,
            carryout => \b2v_inst4.un1_pix_count_int_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst4.un1_pix_count_int_cry_2_c_RNIMI4I_LC_5_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15238\,
            in2 => \_gnd_net_\,
            in3 => \N__13976\,
            lcout => \b2v_inst4.un1_pix_count_int_cry_2_c_RNIMI4IZ0\,
            ltout => OPEN,
            carryin => \b2v_inst4.un1_pix_count_int_cry_2\,
            carryout => \b2v_inst4.un1_pix_count_int_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst4.pix_count_int_4_LC_5_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16727\,
            in2 => \_gnd_net_\,
            in3 => \N__13973\,
            lcout => \SYNTHESIZED_WIRE_4_4\,
            ltout => OPEN,
            carryin => \b2v_inst4.un1_pix_count_int_cry_3\,
            carryout => \b2v_inst4.un1_pix_count_int_cry_4\,
            clk => \N__34502\,
            ce => 'H',
            sr => \N__38059\
        );

    \b2v_inst4.un1_pix_count_int_cry_4_c_RNIQO6I_LC_5_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15827\,
            in2 => \_gnd_net_\,
            in3 => \N__13955\,
            lcout => \b2v_inst4.un1_pix_count_int_cry_4_c_RNIQO6IZ0\,
            ltout => OPEN,
            carryin => \b2v_inst4.un1_pix_count_int_cry_4\,
            carryout => \b2v_inst4.un1_pix_count_int_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst4.un1_pix_count_int_cry_5_c_RNISR7I_LC_5_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15877\,
            in2 => \_gnd_net_\,
            in3 => \N__13931\,
            lcout => \b2v_inst4.un1_pix_count_int_cry_5_c_RNISR7IZ0\,
            ltout => OPEN,
            carryin => \b2v_inst4.un1_pix_count_int_cry_5\,
            carryout => \b2v_inst4.un1_pix_count_int_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst4.pix_count_int_7_LC_5_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16821\,
            in2 => \_gnd_net_\,
            in3 => \N__13928\,
            lcout => \SYNTHESIZED_WIRE_4_7\,
            ltout => OPEN,
            carryin => \b2v_inst4.un1_pix_count_int_cry_6\,
            carryout => \b2v_inst4.un1_pix_count_int_cry_7\,
            clk => \N__34502\,
            ce => 'H',
            sr => \N__38059\
        );

    \b2v_inst4.pix_count_int_8_LC_5_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__14790\,
            in1 => \N__15477\,
            in2 => \_gnd_net_\,
            in3 => \N__13925\,
            lcout => \SYNTHESIZED_WIRE_4_8\,
            ltout => OPEN,
            carryin => \bfn_5_14_0_\,
            carryout => \b2v_inst4.un1_pix_count_int_cry_8\,
            clk => \N__34508\,
            ce => 'H',
            sr => \N__38062\
        );

    \b2v_inst4.un1_pix_count_int_cry_8_c_RNI25BI_LC_5_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15564\,
            in2 => \_gnd_net_\,
            in3 => \N__13922\,
            lcout => \b2v_inst4.un1_pix_count_int_cry_8_c_RNI25BIZ0\,
            ltout => OPEN,
            carryin => \b2v_inst4.un1_pix_count_int_cry_8\,
            carryout => \b2v_inst4.un1_pix_count_int_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst4.un1_pix_count_int_cry_9_c_RNIB86J_LC_5_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15616\,
            in2 => \_gnd_net_\,
            in3 => \N__14075\,
            lcout => \b2v_inst4.un1_pix_count_int_cry_9_c_RNIB86JZ0\,
            ltout => OPEN,
            carryin => \b2v_inst4.un1_pix_count_int_cry_9\,
            carryout => \b2v_inst4.un1_pix_count_int_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst4.un1_pix_count_int_cry_10_c_RNIKMUJ_LC_5_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15356\,
            in3 => \N__14072\,
            lcout => \b2v_inst4.un1_pix_count_int_cry_10_c_RNIKMUJZ0\,
            ltout => OPEN,
            carryin => \b2v_inst4.un1_pix_count_int_cry_10\,
            carryout => \b2v_inst4.un1_pix_count_int_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst4.un1_pix_count_int_cry_11_c_RNIMPVJ_LC_5_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15398\,
            in3 => \N__14057\,
            lcout => \b2v_inst4.un1_pix_count_int_cry_11_c_RNIMPVJZ0\,
            ltout => OPEN,
            carryin => \b2v_inst4.un1_pix_count_int_cry_11\,
            carryout => \b2v_inst4.un1_pix_count_int_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst4.pix_count_int_13_LC_5_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16473\,
            in2 => \_gnd_net_\,
            in3 => \N__14054\,
            lcout => \SYNTHESIZED_WIRE_4_13\,
            ltout => OPEN,
            carryin => \b2v_inst4.un1_pix_count_int_cry_12\,
            carryout => \b2v_inst4.un1_pix_count_int_cry_13\,
            clk => \N__34508\,
            ce => 'H',
            sr => \N__38062\
        );

    \b2v_inst4.pix_count_int_14_LC_5_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16354\,
            in2 => \_gnd_net_\,
            in3 => \N__14051\,
            lcout => \SYNTHESIZED_WIRE_4_14\,
            ltout => OPEN,
            carryin => \b2v_inst4.un1_pix_count_int_cry_13\,
            carryout => \b2v_inst4.un1_pix_count_int_cry_14\,
            clk => \N__34508\,
            ce => 'H',
            sr => \N__38062\
        );

    \b2v_inst4.pix_count_int_15_LC_5_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16407\,
            in2 => \_gnd_net_\,
            in3 => \N__14048\,
            lcout => \SYNTHESIZED_WIRE_4_15\,
            ltout => OPEN,
            carryin => \b2v_inst4.un1_pix_count_int_cry_14\,
            carryout => \b2v_inst4.un1_pix_count_int_cry_15\,
            clk => \N__34508\,
            ce => 'H',
            sr => \N__38062\
        );

    \b2v_inst4.pix_count_int_16_LC_5_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__14788\,
            in1 => \N__17598\,
            in2 => \_gnd_net_\,
            in3 => \N__14045\,
            lcout => \SYNTHESIZED_WIRE_4_16\,
            ltout => OPEN,
            carryin => \bfn_5_15_0_\,
            carryout => \b2v_inst4.un1_pix_count_int_cry_16\,
            clk => \N__34513\,
            ce => 'H',
            sr => \N__38065\
        );

    \b2v_inst4.pix_count_int_17_LC_5_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17432\,
            in2 => \_gnd_net_\,
            in3 => \N__14042\,
            lcout => \SYNTHESIZED_WIRE_4_17\,
            ltout => OPEN,
            carryin => \b2v_inst4.un1_pix_count_int_cry_16\,
            carryout => \b2v_inst4.un1_pix_count_int_cry_17\,
            clk => \N__34513\,
            ce => 'H',
            sr => \N__38065\
        );

    \b2v_inst4.pix_count_int_18_LC_5_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17484\,
            in2 => \_gnd_net_\,
            in3 => \N__14039\,
            lcout => \SYNTHESIZED_WIRE_4_18\,
            ltout => OPEN,
            carryin => \b2v_inst4.un1_pix_count_int_cry_17\,
            carryout => \b2v_inst4.un1_pix_count_int_cry_18\,
            clk => \N__34513\,
            ce => 'H',
            sr => \N__38065\
        );

    \b2v_inst4.pix_count_int_19_LC_5_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__14787\,
            in1 => \N__17695\,
            in2 => \_gnd_net_\,
            in3 => \N__14456\,
            lcout => \SYNTHESIZED_WIRE_4_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34513\,
            ce => 'H',
            sr => \N__38065\
        );

    \b2v_inst1.r_RX_Byte_1_LC_5_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__27018\,
            in1 => \N__17299\,
            in2 => \_gnd_net_\,
            in3 => \N__14945\,
            lcout => \SYNTHESIZED_WIRE_10_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34522\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_RNI2OT15_1_LC_5_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__21663\,
            in1 => \N__35217\,
            in2 => \N__20168\,
            in3 => \N__38665\,
            lcout => \SYNTHESIZED_WIRE_12_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_RNIKAU15_7_LC_5_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__35218\,
            in1 => \N__21664\,
            in2 => \N__18893\,
            in3 => \N__38870\,
            lcout => \SYNTHESIZED_WIRE_12_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_RNIVKT15_0_LC_5_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__21665\,
            in1 => \N__39317\,
            in2 => \N__20384\,
            in3 => \N__35219\,
            lcout => \SYNTHESIZED_WIRE_12_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_RNINDU15_8_LC_5_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__35237\,
            in1 => \N__18569\,
            in2 => \N__39101\,
            in3 => \N__21662\,
            lcout => \SYNTHESIZED_WIRE_12_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un2_dir_mem_3_cry_0_c_LC_6_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35701\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_5_0_\,
            carryout => \b2v_inst.un2_dir_mem_3_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_3_RNO_0_6_LC_6_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38337\,
            in2 => \_gnd_net_\,
            in3 => \N__14081\,
            lcout => \b2v_inst.dir_mem_3_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \b2v_inst.un2_dir_mem_3_cry_0\,
            carryout => \b2v_inst.un2_dir_mem_3_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_3_RNO_0_7_LC_6_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38836\,
            in2 => \N__37303\,
            in3 => \N__14078\,
            lcout => \b2v_inst.dir_mem_3_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \b2v_inst.un2_dir_mem_3_cry_1\,
            carryout => \b2v_inst.un2_dir_mem_3_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_3_RNO_0_8_LC_6_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39058\,
            in2 => \_gnd_net_\,
            in3 => \N__14480\,
            lcout => \b2v_inst.dir_mem_3_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \b2v_inst.un2_dir_mem_3_cry_2\,
            carryout => \b2v_inst.un2_dir_mem_3_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_3_RNO_0_9_LC_6_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35915\,
            in2 => \_gnd_net_\,
            in3 => \N__14477\,
            lcout => \b2v_inst.dir_mem_3_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \b2v_inst.un2_dir_mem_3_cry_3\,
            carryout => \b2v_inst.un2_dir_mem_3_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_3_RNO_0_10_LC_6_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__36747\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14474\,
            lcout => \b2v_inst.dir_mem_3_RNO_0Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un1_indice_cry_1_c_LC_6_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39273\,
            in2 => \N__38603\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_6_0_\,
            carryout => \b2v_inst.un1_indice_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un1_indice_cry_1_c_RNIUSJG_LC_6_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36043\,
            in2 => \_gnd_net_\,
            in3 => \N__14471\,
            lcout => \b2v_inst.un1_indice_cry_1_c_RNIUSJGZ0\,
            ltout => OPEN,
            carryin => \b2v_inst.un1_indice_cry_1\,
            carryout => \b2v_inst.un1_indice_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un1_indice_cry_2_c_RNI00LG_LC_6_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36512\,
            in2 => \_gnd_net_\,
            in3 => \N__14468\,
            lcout => \b2v_inst.un1_indice_cry_2_c_RNI00LGZ0\,
            ltout => OPEN,
            carryin => \b2v_inst.un1_indice_cry_2\,
            carryout => \b2v_inst.un1_indice_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un1_indice_cry_3_c_RNI23MG_LC_6_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36363\,
            in2 => \_gnd_net_\,
            in3 => \N__14465\,
            lcout => \b2v_inst.un1_indice_cry_3_c_RNI23MGZ0\,
            ltout => OPEN,
            carryin => \b2v_inst.un1_indice_cry_3\,
            carryout => \b2v_inst.un1_indice_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un1_indice_cry_4_c_RNI46NG_LC_6_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35710\,
            in2 => \_gnd_net_\,
            in3 => \N__14462\,
            lcout => \b2v_inst.un1_indice_cry_4_c_RNI46NGZ0\,
            ltout => OPEN,
            carryin => \b2v_inst.un1_indice_cry_4\,
            carryout => \b2v_inst.un1_indice_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un1_indice_cry_5_c_RNI69OG_LC_6_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38326\,
            in2 => \_gnd_net_\,
            in3 => \N__14459\,
            lcout => \b2v_inst.un1_indice_cry_5_c_RNI69OGZ0\,
            ltout => OPEN,
            carryin => \b2v_inst.un1_indice_cry_5\,
            carryout => \b2v_inst.un1_indice_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un1_indice_cry_6_c_RNI8CPG_LC_6_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38861\,
            in2 => \_gnd_net_\,
            in3 => \N__14507\,
            lcout => \b2v_inst.dir_mem_316lto7\,
            ltout => OPEN,
            carryin => \b2v_inst.un1_indice_cry_6\,
            carryout => \b2v_inst.un1_indice_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un1_indice_cry_7_c_RNIAFQG_LC_6_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39079\,
            in2 => \_gnd_net_\,
            in3 => \N__14504\,
            lcout => \b2v_inst.un1_indice_cry_7_c_RNIAFQGZ0\,
            ltout => OPEN,
            carryin => \b2v_inst.un1_indice_cry_7\,
            carryout => \b2v_inst.un1_indice_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un1_indice_cry_8_c_RNICIRG_LC_6_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35938\,
            in2 => \_gnd_net_\,
            in3 => \N__14501\,
            lcout => \b2v_inst.un1_indice_cry_8_c_RNICIRGZ0\,
            ltout => OPEN,
            carryin => \bfn_6_7_0_\,
            carryout => \b2v_inst.un1_indice_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un1_indice_cry_9_c_RNILAJP_LC_6_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__36746\,
            in3 => \N__14498\,
            lcout => \b2v_inst.un1_indice_cry_9_c_RNILAJPZ0\,
            ltout => OPEN,
            carryin => \b2v_inst.un1_indice_cry_9\,
            carryout => \b2v_inst.un1_indice_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un1_indice_cry_10_THRU_LUT4_0_LC_6_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14495\,
            lcout => \b2v_inst.un1_indice_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.pix_data_reg_4_LC_6_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27086\,
            lcout => \b2v_inst.pix_data_regZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34498\,
            ce => \N__30243\,
            sr => \N__38057\
        );

    \b2v_inst.ignorar_ancho_1_RNO_0_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011111001111"
        )
    port map (
            in0 => \N__14492\,
            in1 => \N__28204\,
            in2 => \N__26033\,
            in3 => \N__14486\,
            lcout => \b2v_inst.ignorar_ancho_1_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst4.pix_count_int_9_LC_6_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14811\,
            lcout => \SYNTHESIZED_WIRE_4_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34468\,
            ce => 'H',
            sr => \N__38052\
        );

    \b2v_inst4.pix_count_int_fast_10_LC_6_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__14834\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \SYNTHESIZED_WIRE_4_fast_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34468\,
            ce => 'H',
            sr => \N__38052\
        );

    \b2v_inst4.pix_count_int_10_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14832\,
            lcout => \SYNTHESIZED_WIRE_4_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34468\,
            ce => 'H',
            sr => \N__38052\
        );

    \b2v_inst4.pix_count_int_10_rep1_LC_6_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14833\,
            lcout => \SYNTHESIZED_WIRE_4_10_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34468\,
            ce => 'H',
            sr => \N__38052\
        );

    \b2v_inst4.pix_count_int_fast_9_LC_6_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14812\,
            lcout => \SYNTHESIZED_WIRE_4_fast_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34468\,
            ce => 'H',
            sr => \N__38052\
        );

    \b2v_inst4.pix_count_int_11_LC_6_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14789\,
            in2 => \_gnd_net_\,
            in3 => \N__14683\,
            lcout => \SYNTHESIZED_WIRE_4_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34468\,
            ce => 'H',
            sr => \N__38052\
        );

    \b2v_inst.un7_pix_count_int_0_I_33_c_RNIGJGQ8_LC_6_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011110000"
        )
    port map (
            in0 => \N__17709\,
            in1 => \N__15410\,
            in2 => \N__17222\,
            in3 => \N__17593\,
            lcout => \b2v_inst.N_482\,
            ltout => \b2v_inst.N_482_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.ignorar_ancho_1_RNO_LC_6_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100010001"
        )
    port map (
            in0 => \N__28184\,
            in1 => \N__14666\,
            in2 => \N__14657\,
            in3 => \N__14539\,
            lcout => \b2v_inst.un1_state_34_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.ignorar_ancho_1_LC_6_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28185\,
            lcout => \b2v_inst.ignorar_anchoZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34478\,
            ce => \N__14654\,
            sr => \N__38058\
        );

    \b2v_inst.cuenta_pixel_RNIBK2I2_10_LC_6_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__14645\,
            in1 => \N__14621\,
            in2 => \N__14594\,
            in3 => \N__14561\,
            lcout => \b2v_inst.N_325\,
            ltout => \b2v_inst.N_325_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.ignorar_anterior_RNO_LC_6_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__14528\,
            in1 => \N__14519\,
            in2 => \N__14510\,
            in3 => \N__28514\,
            lcout => \b2v_inst.un1_state_36_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un7_pix_count_int_0_I_33_c_RNIMVIF1_LC_6_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000011111111"
        )
    port map (
            in0 => \N__17502\,
            in1 => \N__17436\,
            in2 => \N__17727\,
            in3 => \N__17104\,
            lcout => \b2v_inst.un4_pix_count_intlto19_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNI9A7V8_29_LC_6_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101000"
        )
    port map (
            in0 => \N__28183\,
            in1 => \N__15409\,
            in2 => \N__14846\,
            in3 => \N__17217\,
            lcout => \b2v_inst.N_305_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.ignorar_anterior_LC_6_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28174\,
            lcout => \b2v_inst.ignorar_anteriorZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34488\,
            ce => \N__14909\,
            sr => \N__38060\
        );

    \b2v_inst1.r_RX_Byte_RNO_0_0_LC_6_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100011101"
        )
    port map (
            in0 => \N__22832\,
            in1 => \N__16638\,
            in2 => \N__26716\,
            in3 => \N__15434\,
            lcout => \b2v_inst1.N_42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.g1_0_a4_0_LC_6_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010000000"
        )
    port map (
            in0 => \N__15392\,
            in1 => \N__15352\,
            in2 => \N__15774\,
            in3 => \N__15319\,
            lcout => \b2v_inst.N_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst4.state_RNICJOG_0_LC_6_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__14896\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14864\,
            lcout => \b2v_inst4.pix_count_int_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_RX_DV_LC_6_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011100000"
        )
    port map (
            in0 => \N__14865\,
            in1 => \N__22642\,
            in2 => \N__22925\,
            in3 => \N__21165\,
            lcout => \SYNTHESIZED_WIRE_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34499\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un1_state_36_0_a2_0_1_mb_1_LC_6_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17685\,
            in2 => \_gnd_net_\,
            in3 => \N__17565\,
            lcout => \b2v_inst.un1_state_36_0_a2_0_1_mbZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un4_pix_count_intlto18_0_LC_6_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17483\,
            in2 => \_gnd_net_\,
            in3 => \N__17431\,
            lcout => \b2v_inst.un4_pix_count_intlto18Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_RX_Byte_RNO_0_1_LC_6_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100011011"
        )
    port map (
            in0 => \N__16628\,
            in1 => \N__22829\,
            in2 => \N__27022\,
            in3 => \N__15983\,
            lcout => \b2v_inst1.N_40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_1_LC_7_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22106\,
            in2 => \_gnd_net_\,
            in3 => \N__16245\,
            lcout => \b2v_inst.indiceZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34510\,
            ce => \N__22033\,
            sr => \N__38068\
        );

    \b2v_inst.indice_2_LC_7_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__22107\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15087\,
            lcout => \b2v_inst.indiceZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34510\,
            ce => \N__22033\,
            sr => \N__38068\
        );

    \b2v_inst.indice_6_LC_7_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22109\,
            in2 => \_gnd_net_\,
            in3 => \N__16215\,
            lcout => \b2v_inst.indiceZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34510\,
            ce => \N__22033\,
            sr => \N__38068\
        );

    \b2v_inst.indice_3_LC_7_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22108\,
            in2 => \_gnd_net_\,
            in3 => \N__16071\,
            lcout => \b2v_inst.indiceZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34510\,
            ce => \N__22033\,
            sr => \N__38068\
        );

    \b2v_inst.un8_dir_mem_1_cry_0_c_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39304\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_6_0_\,
            carryout => \b2v_inst.un8_dir_mem_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un8_dir_mem_1_cry_0_c_RNI4SNC_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38573\,
            in2 => \N__37288\,
            in3 => \N__14939\,
            lcout => \b2v_inst.un8_dir_mem_1_cry_0_c_RNI4SNCZ0\,
            ltout => OPEN,
            carryin => \b2v_inst.un8_dir_mem_1_cry_0\,
            carryout => \b2v_inst.un8_dir_mem_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un8_dir_mem_1_cry_1_c_RNI6VOC_LC_7_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36050\,
            in2 => \_gnd_net_\,
            in3 => \N__14936\,
            lcout => \b2v_inst.un8_dir_mem_1_cry_1_c_RNI6VOCZ0\,
            ltout => OPEN,
            carryin => \b2v_inst.un8_dir_mem_1_cry_1\,
            carryout => \b2v_inst.un8_dir_mem_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un8_dir_mem_1_cry_2_c_RNI82QC_LC_7_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36499\,
            in2 => \_gnd_net_\,
            in3 => \N__14933\,
            lcout => \b2v_inst.un8_dir_mem_1_cry_2_c_RNI82QCZ0\,
            ltout => OPEN,
            carryin => \b2v_inst.un8_dir_mem_1_cry_2\,
            carryout => \b2v_inst.un8_dir_mem_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un8_dir_mem_1_cry_3_c_RNIA5RC_LC_7_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36357\,
            in2 => \_gnd_net_\,
            in3 => \N__14930\,
            lcout => \b2v_inst.un8_dir_mem_1_cry_3_c_RNIA5RCZ0\,
            ltout => OPEN,
            carryin => \b2v_inst.un8_dir_mem_1_cry_3\,
            carryout => \b2v_inst.un8_dir_mem_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un8_dir_mem_1_cry_4_c_RNIC8SC_LC_7_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35690\,
            in2 => \_gnd_net_\,
            in3 => \N__14966\,
            lcout => \b2v_inst.un8_dir_mem_1_cry_4_c_RNIC8SCZ0\,
            ltout => OPEN,
            carryin => \b2v_inst.un8_dir_mem_1_cry_4\,
            carryout => \b2v_inst.un8_dir_mem_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un8_dir_mem_1_cry_5_c_RNIEBTC_LC_7_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38327\,
            in2 => \_gnd_net_\,
            in3 => \N__14963\,
            lcout => \b2v_inst.un8_dir_mem_1_cry_5_c_RNIEBTCZ0\,
            ltout => OPEN,
            carryin => \b2v_inst.un8_dir_mem_1_cry_5\,
            carryout => \b2v_inst.un8_dir_mem_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un8_dir_mem_1_cry_6_c_RNIGEUC_LC_7_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38860\,
            in3 => \N__14960\,
            lcout => \b2v_inst.dir_mem_115lto7\,
            ltout => OPEN,
            carryin => \b2v_inst.un8_dir_mem_1_cry_6\,
            carryout => \b2v_inst.un8_dir_mem_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un8_dir_mem_1_cry_7_c_RNIIHVC_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39080\,
            in2 => \_gnd_net_\,
            in3 => \N__14957\,
            lcout => \b2v_inst.un8_dir_mem_1_cry_7_c_RNIIHVCZ0\,
            ltout => OPEN,
            carryin => \bfn_7_7_0_\,
            carryout => \b2v_inst.un8_dir_mem_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un8_dir_mem_1_cry_8_c_RNIKK0D_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35939\,
            in2 => \_gnd_net_\,
            in3 => \N__14954\,
            lcout => \b2v_inst.un8_dir_mem_1_cry_8_c_RNIKK0DZ0\,
            ltout => OPEN,
            carryin => \b2v_inst.un8_dir_mem_1_cry_8\,
            carryout => \b2v_inst.un8_dir_mem_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un8_dir_mem_1_cry_9_c_RNITCOL_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36710\,
            in2 => \_gnd_net_\,
            in3 => \N__14951\,
            lcout => \b2v_inst.un8_dir_mem_1_cry_9_c_RNITCOLZ0\,
            ltout => OPEN,
            carryin => \b2v_inst.un8_dir_mem_1_cry_9\,
            carryout => \b2v_inst.un8_dir_mem_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un8_dir_mem_1_cry_10_THRU_LUT4_0_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14948\,
            lcout => \b2v_inst.un8_dir_mem_1_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un1_indice_cry_6_c_RNIRCFH4_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010000000"
        )
    port map (
            in0 => \N__20310\,
            in1 => \N__18796\,
            in2 => \N__18780\,
            in3 => \N__15098\,
            lcout => \b2v_inst.dir_mem_316lt11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un1_indice_cry_10_c_RNIO00U_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16150\,
            in2 => \_gnd_net_\,
            in3 => \N__20337\,
            lcout => \b2v_inst.dir_mem_316lto11_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_RNIJFGT1_0_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__15088\,
            in1 => \N__16072\,
            in2 => \N__16250\,
            in3 => \N__18351\,
            lcout => OPEN,
            ltout => \b2v_inst.dir_mem_316lt6_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un1_indice_cry_4_c_RNITUVU2_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__16216\,
            in1 => \_gnd_net_\,
            in2 => \N__15101\,
            in3 => \N__18834\,
            lcout => \b2v_inst.dir_mem_316lt7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_3_2_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111100100000"
        )
    port map (
            in0 => \N__15092\,
            in1 => \N__18262\,
            in2 => \N__18323\,
            in3 => \N__36092\,
            lcout => \b2v_inst.dir_mem_3Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34479\,
            ce => \N__18208\,
            sr => \_gnd_net_\
        );

    \b2v_inst.g0_0_i_a4_0_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000000000"
        )
    port map (
            in0 => \N__15068\,
            in1 => \N__15062\,
            in2 => \N__15734\,
            in3 => \N__15681\,
            lcout => OPEN,
            ltout => \b2v_inst.N_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.g0_0_i_2_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__16430\,
            in1 => \N__16363\,
            in2 => \N__15053\,
            in3 => \N__16502\,
            lcout => \b2v_inst.g0_0_iZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un4_pix_count_intlto10_1_0_0_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__16424\,
            in1 => \N__16358\,
            in2 => \_gnd_net_\,
            in3 => \N__16494\,
            lcout => \b2v_inst.un4_pix_count_intlto10_1_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.g0_1_1_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__15050\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15023\,
            lcout => \b2v_inst.g0_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un4_pix_count_intlto15_1_a0_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010000000"
        )
    port map (
            in0 => \N__15344\,
            in1 => \N__15396\,
            in2 => \N__15546\,
            in3 => \N__15599\,
            lcout => \b2v_inst.un4_pix_count_intlto15_1_aZ0Z0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un4_pix_count_intlto6_1_ns_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__15002\,
            in1 => \N__14993\,
            in2 => \_gnd_net_\,
            in3 => \N__14981\,
            lcout => OPEN,
            ltout => \b2v_inst.un4_pix_count_intlt8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un4_pix_count_intlto10_1_0_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001000"
        )
    port map (
            in0 => \N__16266\,
            in1 => \N__15425\,
            in2 => \N__15419\,
            in3 => \N__15416\,
            lcout => \b2v_inst.un4_pix_count_intlt16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNO_25_29_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010000000"
        )
    port map (
            in0 => \N__15397\,
            in1 => \N__15345\,
            in2 => \N__15778\,
            in3 => \N__15320\,
            lcout => \b2v_inst.state_RNO_25Z0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_RX_Byte_RNO_0_4_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__17011\,
            in1 => \_gnd_net_\,
            in2 => \N__17060\,
            in3 => \N__16640\,
            lcout => OPEN,
            ltout => \b2v_inst1.r_RX_Bytece_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_RX_Byte_4_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110011001100"
        )
    port map (
            in0 => \N__22831\,
            in1 => \N__26773\,
            in2 => \N__15287\,
            in3 => \N__17285\,
            lcout => \SYNTHESIZED_WIRE_10_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34469\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_SM_Main_RNIHNPV1_2_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__16904\,
            in1 => \N__22627\,
            in2 => \N__22733\,
            in3 => \N__16536\,
            lcout => \b2v_inst1.N_47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un4_pix_count_intlto10_1_d_0_x1_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100011111"
        )
    port map (
            in0 => \N__15529\,
            in1 => \N__15598\,
            in2 => \N__15682\,
            in3 => \N__15499\,
            lcout => OPEN,
            ltout => \b2v_inst.un4_pix_count_intlto10_1_d_0_xZ0Z1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un4_pix_count_intlto10_1_d_0_ns_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__37217\,
            in1 => \_gnd_net_\,
            in2 => \N__15284\,
            in3 => \N__15730\,
            lcout => \b2v_inst.un4_pix_count_intlto10_1_d_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_RX_Byte_RNO_0_6_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__16639\,
            in1 => \N__17056\,
            in2 => \_gnd_net_\,
            in3 => \N__17010\,
            lcout => \b2v_inst1.r_RX_Bytece_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNO_24_29_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011111111111"
        )
    port map (
            in0 => \N__15280\,
            in1 => \N__15237\,
            in2 => \N__15200\,
            in3 => \N__15139\,
            lcout => OPEN,
            ltout => \b2v_inst.un4_pix_count_intlto6_d_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNO_13_29_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111110111"
        )
    port map (
            in0 => \N__15876\,
            in1 => \N__15826\,
            in2 => \N__15782\,
            in3 => \N__16744\,
            lcout => \b2v_inst.g2_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.g0_0_i_a4_0_1_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__15773\,
            in1 => \N__15547\,
            in2 => \N__15634\,
            in3 => \N__15500\,
            lcout => \b2v_inst.g0_0_i_a4Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un4_pix_count_intlto12_0_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__15729\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15683\,
            lcout => b2v_inst_un4_pix_count_intlto12_0,
            ltout => \b2v_inst_un4_pix_count_intlto12_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.g1_0_a4_0_1_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__15609\,
            in1 => \N__15548\,
            in2 => \N__15506\,
            in3 => \N__15501\,
            lcout => \b2v_inst.g1_0_a4Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_SM_Main_ns_2_0__m13_i_o2_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__16632\,
            in1 => \N__17041\,
            in2 => \_gnd_net_\,
            in3 => \N__16995\,
            lcout => \b2v_inst1.N_49\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNIB55E1_6_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__37789\,
            in1 => \N__24740\,
            in2 => \N__35322\,
            in3 => \N__37496\,
            lcout => \N_457_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_RX_Byte_RNO_1_0_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17042\,
            in2 => \_gnd_net_\,
            in3 => \N__16996\,
            lcout => \b2v_inst1.N_48\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_Bit_Index_RNIBK4I_1_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111101011111"
        )
    port map (
            in0 => \N__16997\,
            in1 => \_gnd_net_\,
            in2 => \N__17055\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst1.N_44\,
            ltout => \b2v_inst1.N_44_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_Bit_Index_2_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001001"
        )
    port map (
            in0 => \N__16003\,
            in1 => \N__16630\,
            in2 => \N__15428\,
            in3 => \N__16019\,
            lcout => \b2v_inst1.r_Bit_IndexZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34489\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.g1_0_0_2_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__16423\,
            in1 => \N__16350\,
            in2 => \N__16034\,
            in3 => \N__16498\,
            lcout => \b2v_inst.g1_0_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_RX_Byte_0_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__26712\,
            in1 => \N__17289\,
            in2 => \_gnd_net_\,
            in3 => \N__16025\,
            lcout => \SYNTHESIZED_WIRE_10_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34489\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_Bit_Index_0_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000010001"
        )
    port map (
            in0 => \N__16998\,
            in1 => \N__16015\,
            in2 => \_gnd_net_\,
            in3 => \N__16002\,
            lcout => \b2v_inst1.r_Bit_IndexZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34489\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNI75II_29_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28197\,
            in2 => \_gnd_net_\,
            in3 => \N__17714\,
            lcout => \b2v_inst.g3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_SM_Main_RNIC98H_2_LC_7_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__22908\,
            in1 => \N__22720\,
            in2 => \_gnd_net_\,
            in3 => \N__22638\,
            lcout => \b2v_inst1.r_SM_Main_d_4\,
            ltout => \b2v_inst1.r_SM_Main_d_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_Bit_Index_1_LC_7_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100100001010"
        )
    port map (
            in0 => \N__17048\,
            in1 => \N__16004\,
            in2 => \N__15986\,
            in3 => \N__17012\,
            lcout => \b2v_inst1.r_Bit_IndexZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34500\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_RX_Byte_RNO_1_1_LC_7_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17046\,
            in2 => \_gnd_net_\,
            in3 => \N__16999\,
            lcout => \b2v_inst1.N_51\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_RNIQGU15_9_LC_7_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__16649\,
            in1 => \N__21654\,
            in2 => \N__35952\,
            in3 => \N__35216\,
            lcout => \SYNTHESIZED_WIRE_12_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_RX_Byte_RNO_0_5_LC_7_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__16627\,
            in1 => \N__17047\,
            in2 => \_gnd_net_\,
            in3 => \N__17000\,
            lcout => \b2v_inst1.r_RX_Bytece_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_RNIJFHB_0_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38574\,
            in2 => \_gnd_net_\,
            in3 => \N__39303\,
            lcout => \b2v_inst.indice_RNIJFHBZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_8_5_0_\,
            carryout => \b2v_inst.un2_dir_mem_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_RNILHHB_2_LC_8_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__38575\,
            in1 => \N__36044\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst.indice_RNILHHBZ0Z_2\,
            ltout => OPEN,
            carryin => \b2v_inst.un2_dir_mem_1_cry_0\,
            carryout => \b2v_inst.un2_dir_mem_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un2_dir_mem_1_cry_2_c_LC_8_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36527\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.un2_dir_mem_1_cry_1\,
            carryout => \b2v_inst.un2_dir_mem_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un2_dir_mem_1_cry_3_c_LC_8_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36337\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.un2_dir_mem_1_cry_2\,
            carryout => \b2v_inst.un2_dir_mem_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_1_RNO_0_5_LC_8_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35700\,
            in2 => \N__37158\,
            in3 => \N__16049\,
            lcout => \b2v_inst.dir_mem_1_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \b2v_inst.un2_dir_mem_1_cry_3\,
            carryout => \b2v_inst.un2_dir_mem_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_1_RNO_0_6_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38338\,
            in2 => \_gnd_net_\,
            in3 => \N__16046\,
            lcout => \b2v_inst.dir_mem_1_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \b2v_inst.un2_dir_mem_1_cry_4\,
            carryout => \b2v_inst.un2_dir_mem_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_1_RNO_0_7_LC_8_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38829\,
            in2 => \N__37159\,
            in3 => \N__16043\,
            lcout => \b2v_inst.dir_mem_1_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \b2v_inst.un2_dir_mem_1_cry_5\,
            carryout => \b2v_inst.un2_dir_mem_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_1_RNO_0_8_LC_8_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39068\,
            in2 => \_gnd_net_\,
            in3 => \N__16040\,
            lcout => \b2v_inst.dir_mem_1_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \b2v_inst.un2_dir_mem_1_cry_6\,
            carryout => \b2v_inst.un2_dir_mem_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_1_RNO_0_9_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35920\,
            in2 => \_gnd_net_\,
            in3 => \N__16037\,
            lcout => \b2v_inst.dir_mem_1_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_8_6_0_\,
            carryout => \b2v_inst.un2_dir_mem_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_1_RNO_0_10_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__36728\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16163\,
            lcout => \b2v_inst.dir_mem_1_RNO_0Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un8_dir_mem_1_cry_1_c_RNIS26J1_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__19123\,
            in1 => \N__18013\,
            in2 => \N__19275\,
            in3 => \N__17998\,
            lcout => \b2v_inst.dir_mem_115lt6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_RNIEPAH_4_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__35919\,
            in1 => \N__38313\,
            in2 => \_gnd_net_\,
            in3 => \N__36358\,
            lcout => \b2v_inst.indice_4_i_a2_0_7_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNI3UC9_11_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__25952\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26032\,
            lcout => \b2v_inst.N_442_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_3_0_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000001"
        )
    port map (
            in0 => \N__18254\,
            in1 => \N__20349\,
            in2 => \N__16160\,
            in3 => \N__39306\,
            lcout => \b2v_inst.dir_mem_3Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34490\,
            ce => \N__18209\,
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_3_10_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__20350\,
            in1 => \N__16159\,
            in2 => \N__16139\,
            in3 => \N__18255\,
            lcout => \b2v_inst.dir_mem_3Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34490\,
            ce => \N__18209\,
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_3_7_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010111000"
        )
    port map (
            in0 => \N__18784\,
            in1 => \N__18313\,
            in2 => \N__16121\,
            in3 => \N__18253\,
            lcout => \b2v_inst.dir_mem_3Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34490\,
            ce => \N__18209\,
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_3_8_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011110000"
        )
    port map (
            in0 => \N__18258\,
            in1 => \N__20320\,
            in2 => \N__16106\,
            in3 => \N__18318\,
            lcout => \b2v_inst.dir_mem_3Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34490\,
            ce => \N__18209\,
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_3_9_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010111000"
        )
    port map (
            in0 => \N__18808\,
            in1 => \N__18314\,
            in2 => \N__16091\,
            in3 => \N__18259\,
            lcout => \b2v_inst.dir_mem_3Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34490\,
            ce => \N__18209\,
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_3_3_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111101000000"
        )
    port map (
            in0 => \N__18256\,
            in1 => \N__16076\,
            in2 => \N__18324\,
            in3 => \N__36565\,
            lcout => \b2v_inst.dir_mem_3Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34490\,
            ce => \N__18209\,
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_3_5_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010111000101"
        )
    port map (
            in0 => \N__35705\,
            in1 => \N__18841\,
            in2 => \N__18325\,
            in3 => \N__18257\,
            lcout => \b2v_inst.dir_mem_3Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34490\,
            ce => \N__18209\,
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_3_1_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111100100000"
        )
    port map (
            in0 => \N__16246\,
            in1 => \N__18260\,
            in2 => \N__18322\,
            in3 => \N__38640\,
            lcout => \b2v_inst.dir_mem_3Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34480\,
            ce => \N__18204\,
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_3_6_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__18306\,
            in1 => \N__16220\,
            in2 => \N__16193\,
            in3 => \N__18261\,
            lcout => \b2v_inst.dir_mem_3Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34480\,
            ce => \N__18204\,
            sr => \_gnd_net_\
        );

    \b2v_inst.un3_dir_mem_cry_0_c_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39305\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_9_0_\,
            carryout => \b2v_inst.un3_dir_mem_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un3_dir_mem_cry_1_c_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38642\,
            in2 => \N__37157\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.un3_dir_mem_cry_0\,
            carryout => \b2v_inst.un3_dir_mem_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_2_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36103\,
            in2 => \N__37152\,
            in3 => \N__16175\,
            lcout => \b2v_inst.dir_memZ0Z_2\,
            ltout => OPEN,
            carryin => \b2v_inst.un3_dir_mem_cry_1\,
            carryout => \b2v_inst.un3_dir_mem_cry_2\,
            clk => \N__34470\,
            ce => \N__22170\,
            sr => \N__38061\
        );

    \b2v_inst.dir_mem_3_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36570\,
            in2 => \N__37155\,
            in3 => \N__16172\,
            lcout => \b2v_inst.dir_memZ0Z_3\,
            ltout => OPEN,
            carryin => \b2v_inst.un3_dir_mem_cry_2\,
            carryout => \b2v_inst.un3_dir_mem_cry_3\,
            clk => \N__34470\,
            ce => \N__22170\,
            sr => \N__38061\
        );

    \b2v_inst.dir_mem_4_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36359\,
            in2 => \N__37153\,
            in3 => \N__16169\,
            lcout => \b2v_inst.dir_memZ0Z_4\,
            ltout => OPEN,
            carryin => \b2v_inst.un3_dir_mem_cry_3\,
            carryout => \b2v_inst.un3_dir_mem_cry_4\,
            clk => \N__34470\,
            ce => \N__22170\,
            sr => \N__38061\
        );

    \b2v_inst.dir_mem_RNO_0_5_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37063\,
            in2 => \N__35715\,
            in3 => \N__16166\,
            lcout => \b2v_inst.dir_mem_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \b2v_inst.un3_dir_mem_cry_4\,
            carryout => \b2v_inst.un3_dir_mem_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_RNO_0_6_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38359\,
            in2 => \N__37154\,
            in3 => \N__16517\,
            lcout => \b2v_inst.dir_mem_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \b2v_inst.un3_dir_mem_cry_5\,
            carryout => \b2v_inst.un3_dir_mem_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_7_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38847\,
            in2 => \N__37156\,
            in3 => \N__16514\,
            lcout => \b2v_inst.dir_memZ0Z_7\,
            ltout => OPEN,
            carryin => \b2v_inst.un3_dir_mem_cry_6\,
            carryout => \b2v_inst.un3_dir_mem_cry_7\,
            clk => \N__34470\,
            ce => \N__22170\,
            sr => \N__38061\
        );

    \b2v_inst.dir_mem_RNO_0_8_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39069\,
            in2 => \N__37151\,
            in3 => \N__16511\,
            lcout => \b2v_inst.dir_mem_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \bfn_8_10_0_\,
            carryout => \b2v_inst.un3_dir_mem_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_RNO_0_9_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37056\,
            in2 => \N__35954\,
            in3 => \N__16508\,
            lcout => \b2v_inst.dir_mem_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \b2v_inst.un3_dir_mem_cry_8\,
            carryout => \b2v_inst.un3_dir_mem_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_10_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36745\,
            in2 => \_gnd_net_\,
            in3 => \N__16505\,
            lcout => \b2v_inst.dir_memZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34458\,
            ce => \N__22187\,
            sr => \N__38056\
        );

    \b2v_inst.state_RNO_14_29_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__16501\,
            in1 => \N__16425\,
            in2 => \N__16364\,
            in3 => \N__16289\,
            lcout => OPEN,
            ltout => \b2v_inst.m29_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNO_5_29_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001000000"
        )
    port map (
            in0 => \N__16853\,
            in1 => \N__16283\,
            in2 => \N__16274\,
            in3 => \N__16267\,
            lcout => \b2v_inst.o2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_Clk_Count_RNI64771_0_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__16905\,
            in1 => \N__21077\,
            in2 => \_gnd_net_\,
            in3 => \N__21108\,
            lcout => \b2v_inst1.un22_r_clk_count_ac0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNO_20_29_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__25686\,
            in1 => \N__26075\,
            in2 => \N__25742\,
            in3 => \N__25439\,
            lcout => \b2v_inst.N_618_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_Clk_Count_RNI4O4Q_0_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__21109\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16906\,
            lcout => \b2v_inst1.N_119\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNO_22_29_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__30875\,
            in1 => \N__24658\,
            in2 => \N__28201\,
            in3 => \N__25827\,
            lcout => \b2v_inst.G_40_i_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_SM_Main_ns_2_0__m13_i_a3_2_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__22643\,
            in1 => \N__21181\,
            in2 => \N__22924\,
            in3 => \N__21082\,
            lcout => \b2v_inst1.N_96\,
            ltout => \b2v_inst1.N_96_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_Clk_Count_0_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001000001100"
        )
    port map (
            in0 => \N__22724\,
            in1 => \N__21150\,
            in2 => \N__16577\,
            in3 => \N__21112\,
            lcout => \b2v_inst1.r_Clk_CountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34459\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.g0_0_i_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011001110"
        )
    port map (
            in0 => \N__16574\,
            in1 => \N__16568\,
            in2 => \N__16559\,
            in3 => \N__16848\,
            lcout => \b2v_inst.N_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_Clk_Count_RNO_0_2_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001001100110011"
        )
    port map (
            in0 => \N__21111\,
            in1 => \N__16902\,
            in2 => \N__21083\,
            in3 => \N__21145\,
            lcout => OPEN,
            ltout => \b2v_inst1.N_58_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_Clk_Count_2_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100001010"
        )
    port map (
            in0 => \N__21146\,
            in1 => \_gnd_net_\,
            in2 => \N__16544\,
            in3 => \N__22713\,
            lcout => \b2v_inst1.r_Clk_CountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34471\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_SM_Main_2_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__22626\,
            in1 => \N__20902\,
            in2 => \_gnd_net_\,
            in3 => \N__22916\,
            lcout => \b2v_inst1.r_SM_MainZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34471\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_Clk_Count_RNIGMPV1_2_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110011111100"
        )
    port map (
            in0 => \N__16540\,
            in1 => \N__22624\,
            in2 => \N__22923\,
            in3 => \N__16903\,
            lcout => \b2v_inst1.N_43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_RX_Byte_6_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__16919\,
            in1 => \N__22830\,
            in2 => \N__26761\,
            in3 => \N__17290\,
            lcout => \SYNTHESIZED_WIRE_10_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34471\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_SM_Main_ns_2_0__m16_0_o2_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101110111"
        )
    port map (
            in0 => \N__16901\,
            in1 => \N__21078\,
            in2 => \_gnd_net_\,
            in3 => \N__21110\,
            lcout => \b2v_inst1.m16_0_o2\,
            ltout => \b2v_inst1.m16_0_o2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_SM_Main_ns_2_0__m13_i_2_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110001001000"
        )
    port map (
            in0 => \N__22625\,
            in1 => \N__22915\,
            in2 => \N__16865\,
            in3 => \N__17314\,
            lcout => \b2v_inst1.m13_i_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.g1_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000110010"
        )
    port map (
            in0 => \N__16862\,
            in1 => \N__16842\,
            in2 => \N__16775\,
            in3 => \N__16745\,
            lcout => \b2v_inst.g1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.g0_1_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110000000000"
        )
    port map (
            in0 => \N__16688\,
            in1 => \N__16682\,
            in2 => \N__16676\,
            in3 => \N__17611\,
            lcout => \b2v_inst.g3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_energia_RNID0NB2_9_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__16667\,
            in1 => \N__21718\,
            in2 => \_gnd_net_\,
            in3 => \N__35819\,
            lcout => \b2v_inst.addr_ram_energia_m0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_RX_Byte_RNO_0_2_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000011111"
        )
    port map (
            in0 => \N__16964\,
            in1 => \N__16631\,
            in2 => \N__26986\,
            in3 => \N__22826\,
            lcout => OPEN,
            ltout => \b2v_inst1.N_38_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_RX_Byte_2_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111100001010"
        )
    port map (
            in0 => \N__17302\,
            in1 => \_gnd_net_\,
            in2 => \N__16643\,
            in3 => \N__26982\,
            lcout => \SYNTHESIZED_WIRE_10_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34481\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_RX_Byte_RNO_0_3_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100011011"
        )
    port map (
            in0 => \N__16629\,
            in1 => \N__22827\,
            in2 => \N__26800\,
            in3 => \N__16583\,
            lcout => OPEN,
            ltout => \b2v_inst1.N_36_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_RX_Byte_3_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111100001010"
        )
    port map (
            in0 => \N__17303\,
            in1 => \_gnd_net_\,
            in2 => \N__17063\,
            in3 => \N__26796\,
            lcout => \SYNTHESIZED_WIRE_10_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34481\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_RX_Byte_RNO_1_2_LC_8_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17054\,
            in2 => \_gnd_net_\,
            in3 => \N__17009\,
            lcout => \b2v_inst1.N_50\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_RX_Byte_5_LC_8_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__17300\,
            in1 => \N__28813\,
            in2 => \N__16958\,
            in3 => \N__22816\,
            lcout => \SYNTHESIZED_WIRE_10_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34491\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNIAD041_9_LC_8_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__37467\,
            in1 => \N__37791\,
            in2 => \N__32872\,
            in3 => \N__24677\,
            lcout => \N_460_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNI79V31_8_LC_8_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__37790\,
            in1 => \N__24692\,
            in2 => \N__33398\,
            in3 => \N__37466\,
            lcout => \N_459_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un8_dir_mem_2_cry_1_c_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38587\,
            in2 => \N__36076\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_5_0_\,
            carryout => \b2v_inst.un8_dir_mem_2_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un8_dir_mem_2_cry_1_c_RNI88LL_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36523\,
            in2 => \_gnd_net_\,
            in3 => \N__16928\,
            lcout => \b2v_inst.un8_dir_mem_2_cry_1_c_RNI88LLZ0\,
            ltout => OPEN,
            carryin => \b2v_inst.un8_dir_mem_2_cry_1\,
            carryout => \b2v_inst.un8_dir_mem_2_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un8_dir_mem_2_cry_2_c_RNIABML_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36309\,
            in2 => \_gnd_net_\,
            in3 => \N__16925\,
            lcout => \b2v_inst.un8_dir_mem_2_cry_2_c_RNIABMLZ0\,
            ltout => OPEN,
            carryin => \b2v_inst.un8_dir_mem_2_cry_2\,
            carryout => \b2v_inst.un8_dir_mem_2_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un8_dir_mem_2_cry_3_c_RNICENL_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35669\,
            in2 => \_gnd_net_\,
            in3 => \N__16922\,
            lcout => \b2v_inst.un8_dir_mem_2_cry_3_c_RNICENLZ0\,
            ltout => OPEN,
            carryin => \b2v_inst.un8_dir_mem_2_cry_3\,
            carryout => \b2v_inst.un8_dir_mem_2_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un8_dir_mem_2_cry_4_c_RNIEHOL_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38342\,
            in2 => \_gnd_net_\,
            in3 => \N__17087\,
            lcout => \b2v_inst.un8_dir_mem_2_cry_4_c_RNIEHOLZ0\,
            ltout => OPEN,
            carryin => \b2v_inst.un8_dir_mem_2_cry_4\,
            carryout => \b2v_inst.un8_dir_mem_2_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un8_dir_mem_2_cry_5_c_RNIGKP5_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38828\,
            in2 => \_gnd_net_\,
            in3 => \N__17084\,
            lcout => \b2v_inst.dir_mem_215lto7\,
            ltout => OPEN,
            carryin => \b2v_inst.un8_dir_mem_2_cry_5\,
            carryout => \b2v_inst.un8_dir_mem_2_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un8_dir_mem_2_cry_6_c_RNIINQ5_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39034\,
            in2 => \_gnd_net_\,
            in3 => \N__17081\,
            lcout => \b2v_inst.un8_dir_mem_2_cry_6_c_RNIINQZ0Z5\,
            ltout => OPEN,
            carryin => \b2v_inst.un8_dir_mem_2_cry_6\,
            carryout => \b2v_inst.un8_dir_mem_2_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un8_dir_mem_2_cry_7_c_RNIKQR5_LC_9_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35911\,
            in2 => \_gnd_net_\,
            in3 => \N__17078\,
            lcout => \b2v_inst.un8_dir_mem_2_cry_7_c_RNIKQRZ0Z5\,
            ltout => OPEN,
            carryin => \b2v_inst.un8_dir_mem_2_cry_7\,
            carryout => \b2v_inst.un8_dir_mem_2_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un8_dir_mem_2_cry_8_c_RNITIJE_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36727\,
            in2 => \_gnd_net_\,
            in3 => \N__17075\,
            lcout => \b2v_inst.un8_dir_mem_2_cry_8_c_RNITIJEZ0\,
            ltout => OPEN,
            carryin => \bfn_9_6_0_\,
            carryout => \b2v_inst.un8_dir_mem_2_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un8_dir_mem_2_cry_9_THRU_LUT4_0_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17072\,
            lcout => \b2v_inst.un8_dir_mem_2_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_RNIHTLS1_1_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__19059\,
            in1 => \N__19035\,
            in2 => \N__19200\,
            in3 => \N__38625\,
            lcout => \b2v_inst.dir_mem_215lt6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un8_dir_mem_2_cry_9_c_RNI1HOE_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20260\,
            in2 => \_gnd_net_\,
            in3 => \N__20241\,
            lcout => \b2v_inst.dir_mem_215lto11_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_RNIBT583_1_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__18997\,
            in1 => \N__18979\,
            in2 => \_gnd_net_\,
            in3 => \N__17069\,
            lcout => \b2v_inst.dir_mem_215lt7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.energia_temp_4_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17185\,
            lcout => b2v_inst_energia_temp_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34482\,
            ce => \N__26144\,
            sr => \N__38069\
        );

    \b2v_inst.energia_temp_5_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17149\,
            lcout => b2v_inst_energia_temp_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34482\,
            ce => \N__26144\,
            sr => \N__38069\
        );

    \b2v_inst.data_a_escribir_RNO_2_5_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__27398\,
            in1 => \N__29560\,
            in2 => \_gnd_net_\,
            in3 => \N__32535\,
            lcout => \b2v_inst.N_273\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un8_dir_mem_1_cry_4_c_RNIMMVC2_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__18112\,
            in1 => \N__17987\,
            in2 => \_gnd_net_\,
            in3 => \N__17120\,
            lcout => \b2v_inst.dir_mem_115lt7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNIQHR9_22_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27837\,
            in2 => \_gnd_net_\,
            in3 => \N__20972\,
            lcout => \b2v_inst.N_362_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_27_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111010101010"
        )
    port map (
            in0 => \N__22150\,
            in1 => \N__31622\,
            in2 => \_gnd_net_\,
            in3 => \N__23016\,
            lcout => \b2v_inst.stateZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34460\,
            ce => 'H',
            sr => \N__38064\
        );

    \b2v_inst.state_28_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32051\,
            in2 => \_gnd_net_\,
            in3 => \N__23017\,
            lcout => \b2v_inst.stateZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34460\,
            ce => 'H',
            sr => \N__38064\
        );

    \b2v_inst.state_RNO_29_29_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__31613\,
            in1 => \N__20947\,
            in2 => \N__22169\,
            in3 => \N__26449\,
            lcout => \b2v_inst.N_618_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNO_23_29_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26074\,
            in2 => \_gnd_net_\,
            in3 => \N__25438\,
            lcout => OPEN,
            ltout => \b2v_inst.g0_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNO_11_29_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__25738\,
            in1 => \N__25685\,
            in2 => \N__17114\,
            in3 => \N__17111\,
            lcout => OPEN,
            ltout => \b2v_inst.g0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNO_4_29_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011111"
        )
    port map (
            in0 => \N__17333\,
            in1 => \N__38259\,
            in2 => \N__17345\,
            in3 => \N__17738\,
            lcout => OPEN,
            ltout => \b2v_inst.G_40_i_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNO_1_29_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001111"
        )
    port map (
            in0 => \N__17620\,
            in1 => \N__17342\,
            in2 => \N__17336\,
            in3 => \N__17728\,
            lcout => \b2v_inst.state_RNO_1Z0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNO_12_29_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__28332\,
            in1 => \N__21892\,
            in2 => \N__19692\,
            in3 => \N__19526\,
            lcout => \b2v_inst.state_ns_i_0_a2_11_a2_0_3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNO_21_29_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__28333\,
            in1 => \N__17327\,
            in2 => \N__19693\,
            in3 => \N__21893\,
            lcout => \b2v_inst.state_ns_i_0_a2_11_o2_4_0_3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_RX_Byte_7_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001011110000"
        )
    port map (
            in0 => \N__22828\,
            in1 => \N__17321\,
            in2 => \N__26737\,
            in3 => \N__17301\,
            lcout => \SYNTHESIZED_WIRE_10_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34452\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNO_0_10_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100010100000"
        )
    port map (
            in0 => \N__17731\,
            in1 => \N__17524\,
            in2 => \N__17381\,
            in3 => \N__17621\,
            lcout => \b2v_inst.pix_count_anterior5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNO_9_29_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__19525\,
            in1 => \N__17234\,
            in2 => \_gnd_net_\,
            in3 => \N__17228\,
            lcout => \b2v_inst.state_ns_i_0_a2_11_o2_4_0_5_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNO_8_29_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111011111111"
        )
    port map (
            in0 => \N__17730\,
            in1 => \N__27058\,
            in2 => \N__17861\,
            in3 => \N__17221\,
            lcout => \b2v_inst.g3_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNO_10_29_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111000"
        )
    port map (
            in0 => \N__17729\,
            in1 => \N__17510\,
            in2 => \N__17201\,
            in3 => \N__17447\,
            lcout => \b2v_inst.G_40_i_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNIBA4S1_29_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101111111"
        )
    port map (
            in0 => \N__17732\,
            in1 => \N__28136\,
            in2 => \N__17380\,
            in3 => \N__17613\,
            lcout => OPEN,
            ltout => \b2v_inst.N_430_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNIO4NID_10_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111100111011"
        )
    port map (
            in0 => \N__17525\,
            in1 => \N__17882\,
            in2 => \N__17513\,
            in3 => \N__17376\,
            lcout => \b2v_inst.N_430_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.g1_0_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17509\,
            in2 => \_gnd_net_\,
            in3 => \N__17446\,
            lcout => \b2v_inst.g1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_10_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100111010001010"
        )
    port map (
            in0 => \N__25484\,
            in1 => \N__28137\,
            in2 => \N__30434\,
            in3 => \N__17360\,
            lcout => \b2v_inst.stateZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34461\,
            ce => 'H',
            sr => \N__38070\
        );

    \b2v_inst.state_RNIMBKA_10_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28233\,
            in2 => \_gnd_net_\,
            in3 => \N__34582\,
            lcout => \b2v_inst.N_481\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_9_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__28234\,
            in1 => \N__18629\,
            in2 => \N__21303\,
            in3 => \N__23018\,
            lcout => \b2v_inst.stateZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34461\,
            ce => 'H',
            sr => \N__38070\
        );

    \b2v_inst.dir_energia_RNICN7Q1_0_0_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__39349\,
            in1 => \N__39122\,
            in2 => \N__35827\,
            in3 => \N__36448\,
            lcout => \b2v_inst.state_ns_0_i_o2_7_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_energia_RNIBM7Q1_0_1_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__38407\,
            in1 => \N__35570\,
            in2 => \N__38909\,
            in3 => \N__38692\,
            lcout => OPEN,
            ltout => \b2v_inst.state_ns_0_i_o2_6_23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_energia_RNIOG7I4_0_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21931\,
            in2 => \N__17354\,
            in3 => \N__17351\,
            lcout => \b2v_inst.N_512\,
            ltout => \b2v_inst.N_512_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNI3EH15_10_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010101"
        )
    port map (
            in0 => \N__23912\,
            in1 => \N__28338\,
            in2 => \N__17885\,
            in3 => \N__28238\,
            lcout => \b2v_inst.N_430_tz\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_energia_RNO_0_0_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111000001010"
        )
    port map (
            in0 => \N__28239\,
            in1 => \N__34973\,
            in2 => \N__21302\,
            in3 => \N__23913\,
            lcout => \b2v_inst.dir_energia_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_energia_RNIBM7Q1_1_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__38408\,
            in1 => \N__35571\,
            in2 => \N__38910\,
            in3 => \N__38693\,
            lcout => OPEN,
            ltout => \b2v_inst.g0_4_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_fast_RNITQVP4_19_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000001"
        )
    port map (
            in0 => \N__17831\,
            in1 => \N__21935\,
            in2 => \N__17873\,
            in3 => \N__26950\,
            lcout => OPEN,
            ltout => \b2v_inst.g0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNI9QDMD_29_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011110010"
        )
    port map (
            in0 => \N__17870\,
            in1 => \N__17857\,
            in2 => \N__17840\,
            in3 => \N__17837\,
            lcout => \b2v_inst.N_352_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_energia_RNICN7Q1_0_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__39123\,
            in1 => \N__36449\,
            in2 => \N__35812\,
            in3 => \N__39350\,
            lcout => \b2v_inst.g0_4_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.energia_temp_10_LC_9_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17821\,
            lcout => b2v_inst_energia_temp_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34492\,
            ce => \N__26198\,
            sr => \N__38081\
        );

    \b2v_inst.energia_temp_11_LC_9_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17782\,
            lcout => b2v_inst_energia_temp_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34501\,
            ce => \N__26206\,
            sr => \N__38088\
        );

    \b2v_inst.energia_temp_7_LC_9_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17765\,
            lcout => b2v_inst_energia_temp_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34501\,
            ce => \N__26206\,
            sr => \N__38088\
        );

    \b2v_inst.indice_4_LC_10_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22096\,
            in2 => \_gnd_net_\,
            in3 => \N__18361\,
            lcout => \b2v_inst.indiceZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34493\,
            ce => \N__22046\,
            sr => \N__38082\
        );

    \b2v_inst.dir_mem_1_3_LC_10_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001010"
        )
    port map (
            in0 => \N__19060\,
            in1 => \N__18017\,
            in2 => \N__19179\,
            in3 => \N__19247\,
            lcout => \b2v_inst.dir_mem_1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34483\,
            ce => \N__19112\,
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_1_4_LC_10_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110010001100"
        )
    port map (
            in0 => \N__19248\,
            in1 => \N__19036\,
            in2 => \N__19180\,
            in3 => \N__18002\,
            lcout => \b2v_inst.dir_mem_1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34483\,
            ce => \N__19112\,
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_1_6_LC_10_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__19168\,
            in1 => \N__17986\,
            in2 => \N__17966\,
            in3 => \N__19246\,
            lcout => \b2v_inst.dir_mem_1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34483\,
            ce => \N__19112\,
            sr => \_gnd_net_\
        );

    \b2v_inst.un8_dir_mem_2_cry_5_c_RNI14MP3_LC_10_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010000000"
        )
    port map (
            in0 => \N__20734\,
            in1 => \N__20701\,
            in2 => \N__20779\,
            in3 => \N__17948\,
            lcout => \b2v_inst.dir_mem_215lt11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un8_dir_mem_1_cry_6_c_RNICBUJ3_LC_10_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010000000"
        )
    port map (
            in0 => \N__18166\,
            in1 => \N__18139\,
            in2 => \N__17921\,
            in3 => \N__17942\,
            lcout => \b2v_inst.dir_mem_115lt11\,
            ltout => \b2v_inst.dir_mem_115lt11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_1_10_LC_10_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__18968\,
            in1 => \N__17936\,
            in2 => \N__17924\,
            in3 => \N__18949\,
            lcout => \b2v_inst.dir_mem_1Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34472\,
            ce => \N__19104\,
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_1_0_LC_10_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100001"
        )
    port map (
            in0 => \N__18967\,
            in1 => \N__19245\,
            in2 => \N__39316\,
            in3 => \N__18950\,
            lcout => \b2v_inst.dir_mem_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34472\,
            ce => \N__19104\,
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_1_7_LC_10_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011110000"
        )
    port map (
            in0 => \N__19242\,
            in1 => \N__17920\,
            in2 => \N__17900\,
            in3 => \N__19167\,
            lcout => \b2v_inst.dir_mem_1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34472\,
            ce => \N__19104\,
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_1_8_LC_10_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__19165\,
            in1 => \N__18167\,
            in2 => \N__18155\,
            in3 => \N__19243\,
            lcout => \b2v_inst.dir_mem_1Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34472\,
            ce => \N__19104\,
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_1_9_LC_10_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011110000"
        )
    port map (
            in0 => \N__19244\,
            in1 => \N__18140\,
            in2 => \N__18128\,
            in3 => \N__19166\,
            lcout => \b2v_inst.dir_mem_1Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34472\,
            ce => \N__19104\,
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_1_5_LC_10_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__19164\,
            in1 => \N__18113\,
            in2 => \N__18089\,
            in3 => \N__19241\,
            lcout => \b2v_inst.dir_mem_1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34472\,
            ce => \N__19104\,
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_1_LC_10_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19282\,
            lcout => \b2v_inst.dir_memZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34462\,
            ce => \N__22188\,
            sr => \N__38071\
        );

    \b2v_inst.dir_mem_1_RNIGHIR_6_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__25248\,
            in1 => \N__18074\,
            in2 => \N__18065\,
            in3 => \N__25340\,
            lcout => \b2v_inst.addr_ram_iv_i_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNIFAD9_28_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22149\,
            in2 => \_gnd_net_\,
            in3 => \N__31604\,
            lcout => \b2v_inst.N_450_i_1\,
            ltout => \b2v_inst.N_450_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_2_RNI91F21_7_LC_10_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__20756\,
            in1 => \N__18050\,
            in2 => \N__18041\,
            in3 => \N__22431\,
            lcout => \b2v_inst.addr_ram_iv_i_0_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_2_RNIT4KM_10_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__22430\,
            in1 => \N__18038\,
            in2 => \N__20228\,
            in3 => \N__22499\,
            lcout => \b2v_inst.addr_ram_iv_i_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_1_RNIEFIR_5_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__25339\,
            in1 => \N__18026\,
            in2 => \N__18527\,
            in3 => \N__25249\,
            lcout => \b2v_inst.addr_ram_iv_i_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.cantidad_temp_5_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__32586\,
            in1 => \N__34761\,
            in2 => \N__18512\,
            in3 => \N__34625\,
            lcout => b2v_inst_cantidad_temp_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34447\,
            ce => 'H',
            sr => \N__38063\
        );

    \b2v_inst.state_0_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110101010"
        )
    port map (
            in0 => \N__19691\,
            in1 => \N__21314\,
            in2 => \_gnd_net_\,
            in3 => \N__28339\,
            lcout => \b2v_inst.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34447\,
            ce => 'H',
            sr => \N__38063\
        );

    \b2v_inst.state_24_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__27059\,
            in1 => \N__28173\,
            in2 => \_gnd_net_\,
            in3 => \N__28526\,
            lcout => \b2v_inst.stateZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34447\,
            ce => 'H',
            sr => \N__38063\
        );

    \b2v_inst.dir_mem_2_RNI3RE21_4_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__18488\,
            in1 => \N__22531\,
            in2 => \N__19019\,
            in3 => \N__22443\,
            lcout => OPEN,
            ltout => \b2v_inst.addr_ram_iv_i_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_RNIN3333_4_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__18368\,
            in1 => \N__35166\,
            in2 => \N__18476\,
            in3 => \N__36367\,
            lcout => \indice_RNIN3333_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_1_RNICDIR_4_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__18377\,
            in1 => \N__25349\,
            in2 => \N__18218\,
            in3 => \N__25260\,
            lcout => \b2v_inst.addr_ram_iv_i_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_3_4_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001010"
        )
    port map (
            in0 => \N__36368\,
            in1 => \N__18362\,
            in2 => \N__18332\,
            in3 => \N__18269\,
            lcout => \b2v_inst.dir_mem_3Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34437\,
            ce => \N__18203\,
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNO_15_29_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__24659\,
            in1 => \N__33167\,
            in2 => \N__30931\,
            in3 => \N__25828\,
            lcout => \b2v_inst.state_ns_i_0_a2_11_o2_4_0_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNO_0_9_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28337\,
            in2 => \_gnd_net_\,
            in3 => \N__34588\,
            lcout => \b2v_inst.state_ns_0_i_a2_0_0_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNO_16_29_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110010"
        )
    port map (
            in0 => \N__27959\,
            in1 => \N__22444\,
            in2 => \N__26021\,
            in3 => \N__25267\,
            lcout => OPEN,
            ltout => \b2v_inst.state_ns_i_0_a2_11_o2_4_0_6_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNO_6_29_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111111111111"
        )
    port map (
            in0 => \N__26014\,
            in1 => \N__27993\,
            in2 => \N__18620\,
            in3 => \N__18617\,
            lcout => OPEN,
            ltout => \b2v_inst.N_4_i_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNO_2_29_LC_10_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000011"
        )
    port map (
            in0 => \N__28138\,
            in1 => \N__18611\,
            in2 => \N__18602\,
            in3 => \N__18599\,
            lcout => \b2v_inst.state_RNO_2Z0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_energia_RNIBUMB2_8_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__18593\,
            in1 => \N__39138\,
            in2 => \_gnd_net_\,
            in3 => \N__21710\,
            lcout => \b2v_inst.addr_ram_energia_m0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_32_rep1_RNIRV8V_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__25537\,
            in1 => \N__21258\,
            in2 => \N__27909\,
            in3 => \N__20210\,
            lcout => \b2v_inst.N_480\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNO_3_29_LC_10_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__20211\,
            in1 => \N__25538\,
            in2 => \N__21265\,
            in3 => \N__18557\,
            lcout => OPEN,
            ltout => \b2v_inst.state_ns_i_0_a2_11_o2_4_0_7_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_29_LC_10_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__18551\,
            in1 => \N__19388\,
            in2 => \N__18545\,
            in3 => \N__18542\,
            lcout => \b2v_inst.stateZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34453\,
            ce => 'H',
            sr => \N__38074\
        );

    \b2v_inst.dir_energia_0_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000110111011000"
        )
    port map (
            in0 => \N__23872\,
            in1 => \N__18533\,
            in2 => \N__37133\,
            in3 => \N__39359\,
            lcout => \b2v_inst.dir_energiaZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34463\,
            ce => \N__23800\,
            sr => \N__38076\
        );

    \b2v_inst.dir_energia_10_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001110101010"
        )
    port map (
            in0 => \N__23996\,
            in1 => \N__23914\,
            in2 => \N__33686\,
            in3 => \N__23873\,
            lcout => \b2v_inst.dir_energiaZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34463\,
            ce => \N__23800\,
            sr => \N__38076\
        );

    \b2v_inst.dir_energia_2_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101100011111010"
        )
    port map (
            in0 => \N__23870\,
            in1 => \N__33139\,
            in2 => \N__23588\,
            in3 => \N__23969\,
            lcout => \b2v_inst.dir_energiaZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34463\,
            ce => \N__23800\,
            sr => \N__38076\
        );

    \b2v_inst.dir_energia_4_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101111110000"
        )
    port map (
            in0 => \N__33337\,
            in1 => \N__23915\,
            in2 => \N__23555\,
            in3 => \N__23875\,
            lcout => \b2v_inst.dir_energiaZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34463\,
            ce => \N__23800\,
            sr => \N__38076\
        );

    \b2v_inst.dir_energia_1_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111011110100010"
        )
    port map (
            in0 => \N__23869\,
            in1 => \N__23967\,
            in2 => \N__34844\,
            in3 => \N__23603\,
            lcout => \b2v_inst.dir_energiaZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34463\,
            ce => \N__23800\,
            sr => \N__38076\
        );

    \b2v_inst.dir_energia_3_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100111110101010"
        )
    port map (
            in0 => \N__23570\,
            in1 => \N__33256\,
            in2 => \N__23977\,
            in3 => \N__23874\,
            lcout => \b2v_inst.dir_energiaZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34463\,
            ce => \N__23800\,
            sr => \N__38076\
        );

    \b2v_inst.dir_energia_5_LC_10_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111011110100010"
        )
    port map (
            in0 => \N__23871\,
            in1 => \N__23968\,
            in2 => \N__37631\,
            in3 => \N__23534\,
            lcout => \b2v_inst.dir_energiaZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34463\,
            ce => \N__23800\,
            sr => \N__38076\
        );

    \b2v_inst.dir_energia_6_LC_10_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010111001100"
        )
    port map (
            in0 => \N__23948\,
            in1 => \N__24056\,
            in2 => \N__35330\,
            in3 => \N__23867\,
            lcout => \b2v_inst.dir_energiaZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34473\,
            ce => \N__23799\,
            sr => \N__38083\
        );

    \b2v_inst.dir_energia_RNI7QMB2_6_LC_10_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__21709\,
            in1 => \N__18749\,
            in2 => \_gnd_net_\,
            in3 => \N__38412\,
            lcout => OPEN,
            ltout => \b2v_inst.addr_ram_energia_m0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_RNIH7U15_6_LC_10_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__38369\,
            in1 => \N__21636\,
            in2 => \N__18728\,
            in3 => \N__35185\,
            lcout => \SYNTHESIZED_WIRE_12_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_energia_7_LC_10_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101111110001010"
        )
    port map (
            in0 => \N__23865\,
            in1 => \N__35504\,
            in2 => \N__23976\,
            in3 => \N__24041\,
            lcout => \b2v_inst.dir_energiaZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34473\,
            ce => \N__23799\,
            sr => \N__38083\
        );

    \b2v_inst.dir_energia_8_LC_10_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010111001100"
        )
    port map (
            in0 => \N__23949\,
            in1 => \N__24026\,
            in2 => \N__33397\,
            in3 => \N__23868\,
            lcout => \b2v_inst.dir_energiaZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34473\,
            ce => \N__23799\,
            sr => \N__38083\
        );

    \b2v_inst.dir_energia_9_LC_10_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111011110100010"
        )
    port map (
            in0 => \N__23866\,
            in1 => \N__23950\,
            in2 => \N__32873\,
            in3 => \N__24011\,
            lcout => \b2v_inst.dir_energiaZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34473\,
            ce => \N__23799\,
            sr => \N__38083\
        );

    \b2v_inst.dir_energia_RNI9SMB2_7_LC_10_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__18914\,
            in1 => \N__38905\,
            in2 => \_gnd_net_\,
            in3 => \N__21708\,
            lcout => \b2v_inst.addr_ram_energia_m0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_15_LC_10_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19733\,
            lcout => b2v_inst_state_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34484\,
            ce => 'H',
            sr => \N__38089\
        );

    \b2v_inst.energia_temp_12_LC_10_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18874\,
            lcout => b2v_inst_energia_temp_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34494\,
            ce => \N__26207\,
            sr => \N__38094\
        );

    \b2v_inst.indice_5_LC_11_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22086\,
            in2 => \_gnd_net_\,
            in3 => \N__18845\,
            lcout => \b2v_inst.indiceZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34485\,
            ce => \N__22057\,
            sr => \N__38090\
        );

    \b2v_inst.indice_9_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18812\,
            in2 => \_gnd_net_\,
            in3 => \N__22088\,
            lcout => \b2v_inst.indiceZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34485\,
            ce => \N__22057\,
            sr => \N__38090\
        );

    \b2v_inst.indice_7_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__22087\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18785\,
            lcout => \b2v_inst.indiceZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34485\,
            ce => \N__22057\,
            sr => \N__38090\
        );

    \b2v_inst.dir_mem_2_2_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__20679\,
            in1 => \N__19210\,
            in2 => \N__21983\,
            in3 => \N__20638\,
            lcout => \b2v_inst.dir_mem_2Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34474\,
            ce => \N__20602\,
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_2_1_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101111110100"
        )
    port map (
            in0 => \N__20643\,
            in1 => \N__20684\,
            in2 => \N__22001\,
            in3 => \N__38656\,
            lcout => \b2v_inst.dir_mem_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34474\,
            ce => \N__20602\,
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_2_3_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__20680\,
            in1 => \N__19067\,
            in2 => \N__21965\,
            in3 => \N__20639\,
            lcout => \b2v_inst.dir_mem_2Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34474\,
            ce => \N__20602\,
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_2_4_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__20681\,
            in1 => \N__19043\,
            in2 => \N__21950\,
            in3 => \N__20640\,
            lcout => \b2v_inst.dir_mem_2Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34474\,
            ce => \N__20602\,
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_2_5_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__20641\,
            in1 => \N__20682\,
            in2 => \N__22358\,
            in3 => \N__19004\,
            lcout => \b2v_inst.dir_mem_2Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34474\,
            ce => \N__20602\,
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_2_6_LC_11_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__20683\,
            in1 => \N__18986\,
            in2 => \N__22343\,
            in3 => \N__20642\,
            lcout => \b2v_inst.dir_mem_2Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34474\,
            ce => \N__20602\,
            sr => \_gnd_net_\
        );

    \b2v_inst.un8_dir_mem_1_cry_10_c_RNI8DCR_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18966\,
            in2 => \_gnd_net_\,
            in3 => \N__18948\,
            lcout => \b2v_inst.dir_mem_115lto11_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNIULR9_26_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27839\,
            in2 => \_gnd_net_\,
            in3 => \N__20948\,
            lcout => \b2v_inst.N_363_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNISJR9_24_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27838\,
            in2 => \_gnd_net_\,
            in3 => \N__30232\,
            lcout => \b2v_inst.N_463_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_1_RNIKLIR_8_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__18932\,
            in1 => \N__25358\,
            in2 => \N__18926\,
            in3 => \N__25256\,
            lcout => \b2v_inst.addr_ram_iv_i_1_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_RNIBMAH_0_3_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__35910\,
            in1 => \N__36347\,
            in2 => \_gnd_net_\,
            in3 => \N__36572\,
            lcout => \b2v_inst.un9_indice_0_a2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_1_RNI67IR_1_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__25257\,
            in1 => \N__19322\,
            in2 => \N__25366\,
            in3 => \N__19256\,
            lcout => \b2v_inst.addr_ram_iv_i_0_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_2_RNITKE21_1_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__22406\,
            in1 => \N__19310\,
            in2 => \N__19301\,
            in3 => \N__22511\,
            lcout => \b2v_inst.addr_ram_iv_i_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_1_1_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111110001011"
        )
    port map (
            in0 => \N__19286\,
            in1 => \N__19178\,
            in2 => \N__38664\,
            in3 => \N__19249\,
            lcout => \b2v_inst.dir_mem_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34454\,
            ce => \N__19111\,
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_1_2_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110010001100"
        )
    port map (
            in0 => \N__19250\,
            in1 => \N__19211\,
            in2 => \N__19181\,
            in3 => \N__19130\,
            lcout => \b2v_inst.dir_mem_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34454\,
            ce => \N__19111\,
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNI72D9_24_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30217\,
            in2 => \_gnd_net_\,
            in3 => \N__32896\,
            lcout => \b2v_inst.N_489\,
            ltout => \b2v_inst.N_489_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_2_RNI7VE21_6_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__19079\,
            in1 => \N__21809\,
            in2 => \N__19070\,
            in3 => \N__22500\,
            lcout => \b2v_inst.addr_ram_iv_i_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_2_RNIB3F21_8_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__21779\,
            in1 => \N__22501\,
            in2 => \N__20723\,
            in3 => \N__22420\,
            lcout => \b2v_inst.addr_ram_iv_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNI3UC9_22_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20964\,
            in2 => \_gnd_net_\,
            in3 => \N__32024\,
            lcout => \b2v_inst.N_488\,
            ltout => \b2v_inst.N_488_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_1_RNIIJIR_7_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__19508\,
            in1 => \N__19499\,
            in2 => \N__19484\,
            in3 => \N__25364\,
            lcout => OPEN,
            ltout => \b2v_inst.addr_ram_iv_i_0_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_RNI6J333_7_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__19481\,
            in1 => \N__35207\,
            in2 => \N__19475\,
            in3 => \N__38843\,
            lcout => \indice_RNI6J333_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNO_0_29_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__22525\,
            in1 => \N__25255\,
            in2 => \N__22445\,
            in3 => \N__25365\,
            lcout => \b2v_inst.state_RNO_0Z0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_26_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32899\,
            in2 => \_gnd_net_\,
            in3 => \N__23005\,
            lcout => \b2v_inst.stateZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34438\,
            ce => 'H',
            sr => \N__38066\
        );

    \b2v_inst.state_RNIB6D9_26_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20942\,
            in2 => \_gnd_net_\,
            in3 => \N__26441\,
            lcout => \b2v_inst.N_490\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_20_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101000001010"
        )
    port map (
            in0 => \N__31666\,
            in1 => \_gnd_net_\,
            in2 => \N__23015\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst.stateZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34438\,
            ce => 'H',
            sr => \N__38066\
        );

    \b2v_inst.state_22_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__26442\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23004\,
            lcout => \b2v_inst.stateZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34438\,
            ce => 'H',
            sr => \N__38066\
        );

    \b2v_inst.dir_mem_1_RNI45IR_0_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__19376\,
            in1 => \N__25347\,
            in2 => \N__19364\,
            in3 => \N__25259\,
            lcout => \b2v_inst.addr_ram_iv_i_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_2_RNIRIE21_0_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__19532\,
            in1 => \N__22527\,
            in2 => \N__20288\,
            in3 => \N__22438\,
            lcout => \b2v_inst.addr_ram_iv_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_2_RNI1PE21_3_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__22439\,
            in1 => \N__19346\,
            in2 => \N__22532\,
            in3 => \N__19334\,
            lcout => OPEN,
            ltout => \b2v_inst.addr_ram_iv_i_0_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_RNIIU233_3_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__19538\,
            in1 => \N__35172\,
            in2 => \N__19661\,
            in3 => \N__36573\,
            lcout => \indice_RNIIU233_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_1_RNIABIR_3_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__25258\,
            in1 => \N__19565\,
            in2 => \N__25363\,
            in3 => \N__19550\,
            lcout => \b2v_inst.addr_ram_iv_i_0_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_0_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39322\,
            lcout => \b2v_inst.dir_memZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34428\,
            ce => \N__22186\,
            sr => \N__38072\
        );

    \b2v_inst.state_RNIEIRN_4_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__25457\,
            in1 => \N__23450\,
            in2 => \N__23430\,
            in3 => \N__28045\,
            lcout => \b2v_inst.N_618_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_3_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101011110000"
        )
    port map (
            in0 => \N__28046\,
            in1 => \_gnd_net_\,
            in2 => \N__23458\,
            in3 => \N__30422\,
            lcout => b2v_inst_state_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34439\,
            ce => 'H',
            sr => \N__38075\
        );

    \b2v_inst.state_7_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101011110000"
        )
    port map (
            in0 => \N__25458\,
            in1 => \_gnd_net_\,
            in2 => \N__23431\,
            in3 => \N__30421\,
            lcout => b2v_inst_state_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34439\,
            ce => 'H',
            sr => \N__38075\
        );

    \b2v_inst.state_4_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21878\,
            in2 => \_gnd_net_\,
            in3 => \N__22968\,
            lcout => b2v_inst_state_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34439\,
            ce => 'H',
            sr => \N__38075\
        );

    \b2v_inst.state_8_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22995\,
            in3 => \N__34626\,
            lcout => b2v_inst_state_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34439\,
            ce => 'H',
            sr => \N__38075\
        );

    \b2v_inst9.fsm_state_ns_i_i_0_a2_2_2_0_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__23451\,
            in1 => \N__23423\,
            in2 => \N__25672\,
            in3 => \N__24660\,
            lcout => \b2v_inst9.fsm_state_ns_i_i_0_a2_2_2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_13_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30420\,
            in2 => \_gnd_net_\,
            in3 => \N__25829\,
            lcout => b2v_inst_state_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34439\,
            ce => 'H',
            sr => \N__38075\
        );

    \b2v_inst.state_RNIB4B9_16_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21018\,
            in2 => \_gnd_net_\,
            in3 => \N__19728\,
            lcout => \b2v_inst.N_514\,
            ltout => \b2v_inst.N_514_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNICSQN_4_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111100000000"
        )
    port map (
            in0 => \N__37680\,
            in1 => \_gnd_net_\,
            in2 => \N__19757\,
            in3 => \N__33325\,
            lcout => \N_116_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNI72PL_16_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__19729\,
            in1 => \N__26934\,
            in2 => \N__21023\,
            in3 => \N__34694\,
            lcout => \b2v_inst.N_477\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_16_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21022\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst.stateZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34448\,
            ce => 'H',
            sr => \N__38077\
        );

    \b2v_inst.data_a_escribir_RNI3R2E1_4_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__37679\,
            in1 => \N__24806\,
            in2 => \N__33336\,
            in3 => \N__37404\,
            lcout => \N_548_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_fast_19_LC_11_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30874\,
            lcout => \b2v_inst.state_fastZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34448\,
            ce => 'H',
            sr => \N__38077\
        );

    \b2v_inst.state_RNICIL71_0_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__28297\,
            in1 => \N__21864\,
            in2 => \N__19700\,
            in3 => \N__20212\,
            lcout => OPEN,
            ltout => \b2v_inst.N_692_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_32_rep1_RNI0G5H1_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__27910\,
            in1 => \N__25524\,
            in2 => \N__19664\,
            in3 => \N__21254\,
            lcout => \b2v_inst.N_247\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNIH20J1_31_LC_11_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21253\,
            in1 => \N__21827\,
            in2 => \N__25531\,
            in3 => \N__20213\,
            lcout => \b2v_inst.N_494\,
            ltout => \b2v_inst.N_494_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_energia_RNITFMB2_1_LC_11_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__20195\,
            in1 => \_gnd_net_\,
            in2 => \N__20171\,
            in3 => \N__38697\,
            lcout => \b2v_inst.addr_ram_energia_m0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_RNIIBV05_10_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__21634\,
            in1 => \N__19778\,
            in2 => \N__36738\,
            in3 => \N__35189\,
            lcout => \SYNTHESIZED_WIRE_12_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_energia_RNIVHMB2_2_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__21707\,
            in1 => \N__20042\,
            in2 => \_gnd_net_\,
            in3 => \N__36146\,
            lcout => OPEN,
            ltout => \b2v_inst.addr_ram_energia_m0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_RNI5RT15_2_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__21631\,
            in1 => \N__35186\,
            in2 => \N__20021\,
            in3 => \N__36114\,
            lcout => \SYNTHESIZED_WIRE_12_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_energia_RNI5OMB2_5_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__21706\,
            in1 => \N__19916\,
            in2 => \_gnd_net_\,
            in3 => \N__35577\,
            lcout => OPEN,
            ltout => \b2v_inst.addr_ram_energia_m0_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_RNIE4U15_5_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__21633\,
            in1 => \N__35706\,
            in2 => \N__19904\,
            in3 => \N__35188\,
            lcout => \SYNTHESIZED_WIRE_12_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_energia_RNIT4122_10_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__21704\,
            in1 => \N__19799\,
            in2 => \_gnd_net_\,
            in3 => \N__36776\,
            lcout => \b2v_inst.addr_ram_energia_m0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_energia_RNI1KMB2_3_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__19772\,
            in1 => \N__36453\,
            in2 => \_gnd_net_\,
            in3 => \N__21705\,
            lcout => OPEN,
            ltout => \b2v_inst.addr_ram_energia_m0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_RNI8UT15_3_LC_11_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__35187\,
            in1 => \N__21632\,
            in2 => \N__20537\,
            in3 => \N__36580\,
            lcout => \SYNTHESIZED_WIRE_12_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.energia_temp_6_LC_11_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20425\,
            lcout => b2v_inst_energia_temp_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34475\,
            ce => \N__26197\,
            sr => \N__38095\
        );

    \b2v_inst.dir_energia_RNIRDMB2_0_LC_11_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__20396\,
            in1 => \N__39376\,
            in2 => \_gnd_net_\,
            in3 => \N__21719\,
            lcout => \b2v_inst.addr_ram_energia_m0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNI9PQN_1_LC_12_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010101010"
        )
    port map (
            in0 => \N__34838\,
            in1 => \N__37732\,
            in2 => \_gnd_net_\,
            in3 => \N__37503\,
            lcout => \N_120_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNI1TMA4_32_LC_12_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111100000000"
        )
    port map (
            in0 => \N__27997\,
            in1 => \N__27960\,
            in2 => \N__25951\,
            in3 => \N__20582\,
            lcout => \b2v_inst.N_432_1\,
            ltout => \b2v_inst.N_432_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_10_LC_12_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20357\,
            in3 => \N__20354\,
            lcout => \b2v_inst.indiceZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34476\,
            ce => \N__22056\,
            sr => \N__38096\
        );

    \b2v_inst.indice_8_LC_12_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20321\,
            in2 => \_gnd_net_\,
            in3 => \N__22085\,
            lcout => \b2v_inst.indiceZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34476\,
            ce => \N__22056\,
            sr => \N__38096\
        );

    \b2v_inst.dir_mem_2_0_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101010110"
        )
    port map (
            in0 => \N__39227\,
            in1 => \N__20248\,
            in2 => \N__20270\,
            in3 => \N__20645\,
            lcout => \b2v_inst.dir_mem_2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34464\,
            ce => \N__20606\,
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_2_10_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__20646\,
            in1 => \N__20269\,
            in2 => \N__22286\,
            in3 => \N__20249\,
            lcout => \b2v_inst.dir_mem_2Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34464\,
            ce => \N__20606\,
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_2_7_LC_12_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010111000"
        )
    port map (
            in0 => \N__20783\,
            in1 => \N__20685\,
            in2 => \N__22328\,
            in3 => \N__20644\,
            lcout => \b2v_inst.dir_mem_2Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34464\,
            ce => \N__20606\,
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_2_8_LC_12_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110010001100"
        )
    port map (
            in0 => \N__20647\,
            in1 => \N__22313\,
            in2 => \N__20690\,
            in3 => \N__20741\,
            lcout => \b2v_inst.dir_mem_2Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34464\,
            ce => \N__20606\,
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_2_9_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010111000"
        )
    port map (
            in0 => \N__20708\,
            in1 => \N__20689\,
            in2 => \N__22301\,
            in3 => \N__20648\,
            lcout => \b2v_inst.dir_mem_2Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34464\,
            ce => \N__20606\,
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_RNIPLHB_0_LC_12_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38793\,
            in2 => \_gnd_net_\,
            in3 => \N__39226\,
            lcout => \b2v_inst.N_648_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNIHQTC2_11_LC_12_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111100001111"
        )
    port map (
            in0 => \N__20591\,
            in1 => \N__20561\,
            in2 => \N__26031\,
            in3 => \N__23749\,
            lcout => \b2v_inst.N_432_1_tz\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNIP0281_0_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__37510\,
            in1 => \N__34974\,
            in2 => \N__37759\,
            in3 => \N__24404\,
            lcout => \N_556_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_RNIBMAH_3_LC_12_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__39027\,
            in1 => \N__35682\,
            in2 => \_gnd_net_\,
            in3 => \N__36571\,
            lcout => \b2v_inst.indice_4_i_a2_0_7_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNIBRQN_3_LC_12_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010101010"
        )
    port map (
            in0 => \N__33254\,
            in1 => \N__37728\,
            in2 => \_gnd_net_\,
            in3 => \N__37509\,
            lcout => \N_117_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNIQFKA_5_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21882\,
            in2 => \_gnd_net_\,
            in3 => \N__34741\,
            lcout => \b2v_inst.N_577_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_1_RNIMNIR_9_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__20888\,
            in1 => \N__25359\,
            in2 => \N__20876\,
            in3 => \N__25254\,
            lcout => \b2v_inst.addr_ram_iv_i_1_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNINBVD1_1_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__24371\,
            in1 => \N__37753\,
            in2 => \N__34839\,
            in3 => \N__37479\,
            lcout => \N_554_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_2_RNIVME21_2_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__22404\,
            in1 => \N__20843\,
            in2 => \N__20828\,
            in3 => \N__22524\,
            lcout => \b2v_inst.addr_ram_iv_i_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_2_RNID5F21_9_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__21746\,
            in1 => \N__22523\,
            in2 => \N__20816\,
            in3 => \N__22405\,
            lcout => \b2v_inst.addr_ram_iv_i_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_1_RNI89IR_2_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__20804\,
            in1 => \N__25348\,
            in2 => \N__20798\,
            in3 => \N__25253\,
            lcout => \b2v_inst.addr_ram_iv_i_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNO_2_31_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__21890\,
            in1 => \N__20986\,
            in2 => \_gnd_net_\,
            in3 => \N__28331\,
            lcout => \b2v_inst.state_ns_a3_i_0_a2_5_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNIG6QI_21_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__26450\,
            in1 => \N__32897\,
            in2 => \N__31667\,
            in3 => \N__32025\,
            lcout => \b2v_inst.N_829\,
            ltout => \b2v_inst.N_829_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNIHMD31_5_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__21888\,
            in1 => \N__34725\,
            in2 => \N__20786\,
            in3 => \N__34623\,
            lcout => \b2v_inst.un1_data_a_escribir_0_sqmuxa_3_i_i_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_32_rep1_RNIKPV5_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27919\,
            in2 => \_gnd_net_\,
            in3 => \N__21889\,
            lcout => OPEN,
            ltout => \b2v_inst.un1_state_23_i_a2_0_a2_0_a2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNI2KE31_9_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011111"
        )
    port map (
            in0 => \N__20987\,
            in1 => \N__34726\,
            in2 => \N__20975\,
            in3 => \N__34624\,
            lcout => \b2v_inst.N_547_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_21_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111010101010"
        )
    port map (
            in0 => \N__20968\,
            in1 => \N__32026\,
            in2 => \_gnd_net_\,
            in3 => \N__22996\,
            lcout => \b2v_inst.stateZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34429\,
            ce => 'H',
            sr => \N__38067\
        );

    \b2v_inst.state_23_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111110100000"
        )
    port map (
            in0 => \N__32898\,
            in1 => \_gnd_net_\,
            in2 => \N__23014\,
            in3 => \N__30233\,
            lcout => \b2v_inst.stateZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34429\,
            ce => 'H',
            sr => \N__38067\
        );

    \b2v_inst.state_25_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__26451\,
            in1 => \N__20946\,
            in2 => \_gnd_net_\,
            in3 => \N__23000\,
            lcout => \b2v_inst.stateZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34429\,
            ce => 'H',
            sr => \N__38067\
        );

    \b2v_inst.cuenta_RNI6BB31_6_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23153\,
            in1 => \N__20918\,
            in2 => \N__23117\,
            in3 => \N__23297\,
            lcout => \b2v_inst.un2_cuentalto10_i_a2_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.cuenta_RNI2E6K_2_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23185\,
            in1 => \N__23215\,
            in2 => \N__24209\,
            in3 => \N__23248\,
            lcout => \b2v_inst.un2_cuentalto10_i_a2_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_SM_Main_ns_2_0__m16_0_a3_0_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__22619\,
            in1 => \N__21190\,
            in2 => \N__21076\,
            in3 => \N__22786\,
            lcout => OPEN,
            ltout => \b2v_inst1.m16_0_a3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_SM_Main_1_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100011111010"
        )
    port map (
            in0 => \N__22863\,
            in1 => \N__20912\,
            in2 => \N__20891\,
            in3 => \N__22620\,
            lcout => \b2v_inst1.r_SM_MainZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34420\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_Clk_Count_RNO_1_1_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__22737\,
            in1 => \N__22862\,
            in2 => \_gnd_net_\,
            in3 => \N__22785\,
            lcout => OPEN,
            ltout => \b2v_inst1.r_Clk_Count_6_iv_0_a3_1_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_Clk_Count_RNO_0_1_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010110011"
        )
    port map (
            in0 => \N__21191\,
            in1 => \N__22738\,
            in2 => \N__21170\,
            in3 => \N__21166\,
            lcout => OPEN,
            ltout => \b2v_inst1.r_Clk_Count_6_iv_0_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_Clk_Count_1_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011000001100"
        )
    port map (
            in0 => \N__21167\,
            in1 => \N__21067\,
            in2 => \N__21122\,
            in3 => \N__21119\,
            lcout => \b2v_inst1.r_Clk_CountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34420\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNO_0_17_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000100000"
        )
    port map (
            in0 => \N__37405\,
            in1 => \N__21008\,
            in2 => \N__34727\,
            in3 => \N__20996\,
            lcout => OPEN,
            ltout => \b2v_inst.N_653_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_17_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011111000"
        )
    port map (
            in0 => \N__28553\,
            in1 => \N__37406\,
            in2 => \N__21026\,
            in3 => \N__28521\,
            lcout => \b2v_inst.stateZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34430\,
            ce => 'H',
            sr => \N__38078\
        );

    \b2v_inst.state_RNO_1_17_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__23055\,
            in1 => \N__23496\,
            in2 => \_gnd_net_\,
            in3 => \N__23718\,
            lcout => \b2v_inst.state_ns_i_a2_1_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.cuenta_RNIKUJV_0_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001101"
        )
    port map (
            in0 => \N__22936\,
            in1 => \N__23300\,
            in2 => \N__24226\,
            in3 => \N__23170\,
            lcout => OPEN,
            ltout => \b2v_inst.cuenta_RNIKUJVZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.cuenta_RNI5AT71_0_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__23131\,
            in1 => \_gnd_net_\,
            in2 => \N__21002\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \b2v_inst.un20_cuentalto10_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un4_cuenta_cry_1_c_RNICQI02_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__23234\,
            in1 => \N__23200\,
            in2 => \N__20999\,
            in3 => \N__23092\,
            lcout => \b2v_inst.un20_cuentalto10_sx\,
            ltout => \b2v_inst.un20_cuentalto10_sx_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un4_cuenta_cry_7_c_RNIO18R2_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__23056\,
            in1 => \N__23497\,
            in2 => \N__20990\,
            in3 => \N__23719\,
            lcout => \b2v_inst.state18_li_0\,
            ltout => \b2v_inst.state18_li_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_18_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23966\,
            in2 => \N__21476\,
            in3 => \N__34706\,
            lcout => \b2v_inst.stateZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34430\,
            ce => 'H',
            sr => \N__38078\
        );

    \b2v_inst.state_RNI1MHN_31_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__25529\,
            in1 => \N__21250\,
            in2 => \N__25899\,
            in3 => \N__37384\,
            lcout => \N_130_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_30_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25530\,
            lcout => \b2v_inst.stateZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34440\,
            ce => 'H',
            sr => \N__38084\
        );

    \b2v_inst.state_32_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21252\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst.stateZ0Z_32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34440\,
            ce => 'H',
            sr => \N__38084\
        );

    \b2v_inst.state_fast_32_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__21251\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst.state_fastZ0Z_32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34440\,
            ce => 'H',
            sr => \N__38084\
        );

    \b2v_inst.state_5_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101100010001000"
        )
    port map (
            in0 => \N__28313\,
            in1 => \N__21312\,
            in2 => \N__21891\,
            in3 => \N__22992\,
            lcout => \b2v_inst.stateZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34440\,
            ce => 'H',
            sr => \N__38084\
        );

    \b2v_inst.state_6_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101000011011100"
        )
    port map (
            in0 => \N__21313\,
            in1 => \N__25437\,
            in2 => \N__28252\,
            in3 => \N__30426\,
            lcout => \b2v_inst.stateZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34440\,
            ce => 'H',
            sr => \N__38084\
        );

    \b2v_inst.state_32_rep1_RNIKTF9_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__25528\,
            in1 => \N__21249\,
            in2 => \_gnd_net_\,
            in3 => \N__27886\,
            lcout => \b2v_inst.N_828\,
            ltout => \b2v_inst.N_828_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNIRG0E1_2_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101011001100"
        )
    port map (
            in0 => \N__33135\,
            in1 => \N__24893\,
            in2 => \N__21209\,
            in3 => \N__37397\,
            lcout => \N_552_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_energia_RNI13OT_11_LC_12_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__36236\,
            in1 => \N__36780\,
            in2 => \N__23825\,
            in3 => \N__36147\,
            lcout => \b2v_inst.state_ns_0_i_o2_8_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNIVL1E1_3_LC_12_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__37396\,
            in1 => \N__37678\,
            in2 => \N__33255\,
            in3 => \N__24866\,
            lcout => \N_550_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_fast_RNI70OJ_32_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__21899\,
            in1 => \N__28293\,
            in2 => \_gnd_net_\,
            in3 => \N__21863\,
            lcout => \b2v_inst.addr_ram_energia_ss0_0_i_o2_i_o2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_6_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101010101010"
        )
    port map (
            in0 => \N__21821\,
            in1 => \N__22248\,
            in2 => \N__22271\,
            in3 => \N__23764\,
            lcout => \b2v_inst.dir_memZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34455\,
            ce => \N__22196\,
            sr => \N__38097\
        );

    \b2v_inst.dir_mem_8_LC_12_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__23763\,
            in1 => \N__22270\,
            in2 => \N__22250\,
            in3 => \N__21794\,
            lcout => \b2v_inst.dir_memZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34455\,
            ce => \N__22196\,
            sr => \N__38097\
        );

    \b2v_inst.dir_mem_9_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__22266\,
            in1 => \N__23765\,
            in2 => \N__21764\,
            in3 => \N__22249\,
            lcout => \b2v_inst.dir_memZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34455\,
            ce => \N__22196\,
            sr => \N__38097\
        );

    \b2v_inst.dir_energia_RNI3MMB2_4_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__21737\,
            in1 => \N__36247\,
            in2 => \_gnd_net_\,
            in3 => \N__21717\,
            lcout => OPEN,
            ltout => \b2v_inst.addr_ram_energia_m0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_RNIB1U15_4_LC_12_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__21635\,
            in1 => \N__35215\,
            in2 => \N__21599\,
            in3 => \N__36377\,
            lcout => \SYNTHESIZED_WIRE_12_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_RX_Data_R_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21494\,
            lcout => \b2v_inst1.r_RX_Data_RZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34465\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_RX_Data_LC_12_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22277\,
            lcout => \b2v_inst1.r_RX_DataZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34465\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_RNIEPAH_5_LC_13_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__39026\,
            in1 => \N__38355\,
            in2 => \_gnd_net_\,
            in3 => \N__35683\,
            lcout => \b2v_inst.un9_indice_0_a2_2\,
            ltout => \b2v_inst.un9_indice_0_a2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_5_LC_13_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__22237\,
            in1 => \N__22214\,
            in2 => \N__22199\,
            in3 => \N__23748\,
            lcout => \b2v_inst.dir_memZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34466\,
            ce => \N__22195\,
            sr => \N__38104\
        );

    \b2v_inst.indice_0_LC_13_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110111011"
        )
    port map (
            in0 => \N__22095\,
            in1 => \N__39242\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst.indiceZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_13_6_0_\,
            carryout => \b2v_inst.un2_dir_mem_2_cry_0\,
            clk => \N__34456\,
            ce => \N__22058\,
            sr => \N__38098\
        );

    \b2v_inst.un2_dir_mem_2_cry_0_THRU_LUT4_0_LC_13_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38646\,
            in2 => \_gnd_net_\,
            in3 => \N__21986\,
            lcout => \b2v_inst.un2_dir_mem_2_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst.un2_dir_mem_2_cry_0\,
            carryout => \b2v_inst.un2_dir_mem_2_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_2_RNO_0_2_LC_13_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__36113\,
            in3 => \N__21968\,
            lcout => \b2v_inst.dir_mem_2_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \b2v_inst.un2_dir_mem_2_cry_1\,
            carryout => \b2v_inst.un2_dir_mem_2_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_2_RNO_0_3_LC_13_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36569\,
            in2 => \_gnd_net_\,
            in3 => \N__21953\,
            lcout => \b2v_inst.dir_mem_2_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \b2v_inst.un2_dir_mem_2_cry_2\,
            carryout => \b2v_inst.un2_dir_mem_2_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_2_RNO_0_4_LC_13_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__36375\,
            in3 => \N__21938\,
            lcout => \b2v_inst.dir_mem_2_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \b2v_inst.un2_dir_mem_2_cry_3\,
            carryout => \b2v_inst.un2_dir_mem_2_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_2_RNO_0_5_LC_13_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35711\,
            in2 => \N__37307\,
            in3 => \N__22346\,
            lcout => \b2v_inst.dir_mem_2_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \b2v_inst.un2_dir_mem_2_cry_4\,
            carryout => \b2v_inst.un2_dir_mem_2_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_2_RNO_0_6_LC_13_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38370\,
            in2 => \_gnd_net_\,
            in3 => \N__22331\,
            lcout => \b2v_inst.dir_mem_2_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \b2v_inst.un2_dir_mem_2_cry_5\,
            carryout => \b2v_inst.un2_dir_mem_2_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_2_RNO_0_7_LC_13_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37263\,
            in2 => \N__38862\,
            in3 => \N__22316\,
            lcout => \b2v_inst.dir_mem_2_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \b2v_inst.un2_dir_mem_2_cry_6\,
            carryout => \b2v_inst.un2_dir_mem_2_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_2_RNO_0_8_LC_13_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39049\,
            in2 => \_gnd_net_\,
            in3 => \N__22304\,
            lcout => \b2v_inst.dir_mem_2_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \bfn_13_7_0_\,
            carryout => \b2v_inst.un2_dir_mem_2_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_2_RNO_0_9_LC_13_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35937\,
            in2 => \_gnd_net_\,
            in3 => \N__22292\,
            lcout => \b2v_inst.dir_mem_2_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \b2v_inst.un2_dir_mem_2_cry_8\,
            carryout => \b2v_inst.un2_dir_mem_2_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_2_RNO_0_10_LC_13_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36697\,
            in2 => \_gnd_net_\,
            in3 => \N__22289\,
            lcout => \b2v_inst.dir_mem_2_RNO_0Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.cuenta_6_LC_13_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__25955\,
            in1 => \N__24273\,
            in2 => \_gnd_net_\,
            in3 => \N__23135\,
            lcout => \b2v_inst.cuentaZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34441\,
            ce => \N__24185\,
            sr => \N__38085\
        );

    \b2v_inst.cuenta_7_LC_13_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__24274\,
            in1 => \N__25957\,
            in2 => \_gnd_net_\,
            in3 => \N__23096\,
            lcout => \b2v_inst.cuentaZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34441\,
            ce => \N__24185\,
            sr => \N__38085\
        );

    \b2v_inst.cuenta_8_LC_13_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__25956\,
            in1 => \N__24275\,
            in2 => \_gnd_net_\,
            in3 => \N__23060\,
            lcout => \b2v_inst.cuentaZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34441\,
            ce => \N__24185\,
            sr => \N__38085\
        );

    \b2v_inst.cuenta_9_LC_13_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__24276\,
            in1 => \N__25958\,
            in2 => \_gnd_net_\,
            in3 => \N__23501\,
            lcout => \b2v_inst.cuentaZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34441\,
            ce => \N__24185\,
            sr => \N__38085\
        );

    \b2v_inst1.r_SM_Main_ns_2_0__m13_i_a3_1_LC_13_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__22907\,
            in1 => \N__22812\,
            in2 => \_gnd_net_\,
            in3 => \N__22573\,
            lcout => OPEN,
            ltout => \b2v_inst1.N_95_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_SM_Main_0_LC_13_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__22739\,
            in1 => \N__22676\,
            in2 => \N__22661\,
            in3 => \N__22658\,
            lcout => \b2v_inst1.r_SM_MainZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34431\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_2_RNI5TE21_5_LC_13_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__22544\,
            in1 => \N__22526\,
            in2 => \N__22460\,
            in3 => \N__22429\,
            lcout => \b2v_inst.addr_ram_iv_i_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.cuenta_RNIN5ML_10_LC_13_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23512\,
            in1 => \N__23074\,
            in2 => \N__23704\,
            in3 => \N__23273\,
            lcout => \b2v_inst.un2_cuentalto10_i_a2_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst9.data_to_send_esr_RNO_0_5_LC_13_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__24560\,
            in1 => \N__25013\,
            in2 => \N__23036\,
            in3 => \N__30419\,
            lcout => OPEN,
            ltout => \b2v_inst9.data_to_send_10_0_0_0_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst9.data_to_send_esr_5_LC_13_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__25634\,
            in1 => \N__37597\,
            in2 => \N__22370\,
            in3 => \N__24113\,
            lcout => \b2v_inst9.data_to_sendZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34421\,
            ce => \N__24590\,
            sr => \N__38073\
        );

    \b2v_inst9.data_to_send_esr_RNO_0_4_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__24558\,
            in1 => \N__25061\,
            in2 => \N__22367\,
            in3 => \N__30417\,
            lcout => \b2v_inst9.data_to_send_10_0_0_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst9.data_to_send_esr_RNO_0_3_LC_13_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__30418\,
            in1 => \N__25109\,
            in2 => \N__24128\,
            in3 => \N__24559\,
            lcout => OPEN,
            ltout => \b2v_inst9.data_to_send_10_0_0_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst9.data_to_send_esr_3_LC_13_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__33244\,
            in1 => \N__24437\,
            in2 => \N__23039\,
            in3 => \N__25633\,
            lcout => \b2v_inst9.data_to_sendZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34421\,
            ce => \N__24590\,
            sr => \N__38073\
        );

    \b2v_inst9.data_to_send_esr_6_LC_13_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__25635\,
            in1 => \N__35326\,
            in2 => \_gnd_net_\,
            in3 => \N__24353\,
            lcout => \b2v_inst9.data_to_sendZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34421\,
            ce => \N__24590\,
            sr => \N__38073\
        );

    \b2v_inst.cuenta_1_LC_13_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010001000000"
        )
    port map (
            in0 => \N__24254\,
            in1 => \N__22937\,
            in2 => \N__25934\,
            in3 => \N__22994\,
            lcout => \b2v_inst.cuentaZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34411\,
            ce => \N__24181\,
            sr => \N__38079\
        );

    \b2v_inst.state_RNI1P613_32_LC_13_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101000001010"
        )
    port map (
            in0 => \N__23027\,
            in1 => \N__27983\,
            in2 => \N__25933\,
            in3 => \N__27950\,
            lcout => \b2v_inst.N_655\,
            ltout => \b2v_inst.N_655_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.cuenta_0_LC_13_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010111110111"
        )
    port map (
            in0 => \N__23299\,
            in1 => \N__25912\,
            in2 => \N__23021\,
            in3 => \N__22993\,
            lcout => \b2v_inst.cuentaZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34411\,
            ce => \N__24181\,
            sr => \N__38079\
        );

    \b2v_inst.cuenta_RNIR03A_1_LC_13_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23298\,
            in2 => \_gnd_net_\,
            in3 => \N__23268\,
            lcout => \b2v_inst.cuenta_RNIR03AZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.cuenta_2_LC_13_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__25909\,
            in1 => \N__24255\,
            in2 => \_gnd_net_\,
            in3 => \N__23233\,
            lcout => \b2v_inst.cuentaZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34411\,
            ce => \N__24181\,
            sr => \N__38079\
        );

    \b2v_inst.cuenta_3_LC_13_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__24256\,
            in1 => \N__25911\,
            in2 => \_gnd_net_\,
            in3 => \N__23201\,
            lcout => \b2v_inst.cuentaZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34411\,
            ce => \N__24181\,
            sr => \N__38079\
        );

    \b2v_inst.cuenta_4_LC_13_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__25910\,
            in1 => \N__24257\,
            in2 => \_gnd_net_\,
            in3 => \N__23171\,
            lcout => \b2v_inst.cuentaZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34411\,
            ce => \N__24181\,
            sr => \N__38079\
        );

    \b2v_inst.un4_cuenta_cry_1_c_LC_13_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23296\,
            in2 => \N__23272\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_13_12_0_\,
            carryout => \b2v_inst.un4_cuenta_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un4_cuenta_cry_1_c_RNI9V48_LC_13_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23249\,
            in3 => \N__23219\,
            lcout => \b2v_inst.un4_cuenta_cry_1_c_RNI9VZ0Z48\,
            ltout => OPEN,
            carryin => \b2v_inst.un4_cuenta_cry_1\,
            carryout => \b2v_inst.un4_cuenta_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un4_cuenta_cry_2_c_RNIB268_LC_13_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23216\,
            in3 => \N__23189\,
            lcout => \b2v_inst.un4_cuenta_cry_2_c_RNIBZ0Z268\,
            ltout => OPEN,
            carryin => \b2v_inst.un4_cuenta_cry_2\,
            carryout => \b2v_inst.un4_cuenta_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un4_cuenta_cry_3_c_RNID578_LC_13_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23186\,
            in3 => \N__23159\,
            lcout => \b2v_inst.un4_cuenta_cry_3_c_RNIDZ0Z578\,
            ltout => OPEN,
            carryin => \b2v_inst.un4_cuenta_cry_3\,
            carryout => \b2v_inst.un4_cuenta_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un4_cuenta_cry_4_c_RNIF888_LC_13_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24205\,
            in2 => \_gnd_net_\,
            in3 => \N__23156\,
            lcout => \b2v_inst.un4_cuenta_cry_4_c_RNIFZ0Z888\,
            ltout => OPEN,
            carryin => \b2v_inst.un4_cuenta_cry_4\,
            carryout => \b2v_inst.un4_cuenta_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un4_cuenta_cry_5_c_RNIHB98_LC_13_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23152\,
            in2 => \_gnd_net_\,
            in3 => \N__23120\,
            lcout => \b2v_inst.un4_cuenta_cry_5_c_RNIHBZ0Z98\,
            ltout => OPEN,
            carryin => \b2v_inst.un4_cuenta_cry_5\,
            carryout => \b2v_inst.un4_cuenta_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un4_cuenta_cry_6_c_RNIJEA8_LC_13_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23116\,
            in2 => \_gnd_net_\,
            in3 => \N__23081\,
            lcout => \b2v_inst.un4_cuenta_cry_6_c_RNIJEAZ0Z8\,
            ltout => OPEN,
            carryin => \b2v_inst.un4_cuenta_cry_6\,
            carryout => \b2v_inst.un4_cuenta_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un4_cuenta_cry_7_c_RNILHB8_LC_13_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23078\,
            in2 => \_gnd_net_\,
            in3 => \N__23042\,
            lcout => \b2v_inst.un4_cuenta_cry_7_c_RNILHBZ0Z8\,
            ltout => OPEN,
            carryin => \b2v_inst.un4_cuenta_cry_7\,
            carryout => \b2v_inst.un4_cuenta_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un4_cuenta_cry_8_c_RNINKC8_LC_13_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23519\,
            in2 => \_gnd_net_\,
            in3 => \N__23483\,
            lcout => \b2v_inst.un4_cuenta_cry_8_c_RNINKCZ0Z8\,
            ltout => OPEN,
            carryin => \bfn_13_13_0_\,
            carryout => \b2v_inst.un4_cuenta_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un4_cuenta_cry_9_c_RNI01T9_LC_13_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23705\,
            in2 => \_gnd_net_\,
            in3 => \N__23480\,
            lcout => \b2v_inst.un4_cuenta_cry_9_c_RNI01TZ0Z9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNIFA6E1_7_LC_13_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110010101010"
        )
    port map (
            in0 => \N__24701\,
            in1 => \N__35500\,
            in2 => \N__37709\,
            in3 => \N__37449\,
            lcout => \N_458_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst9.data_to_send_esr_RNO_1_0_LC_13_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__24548\,
            in1 => \N__24947\,
            in2 => \N__24475\,
            in3 => \N__34910\,
            lcout => \b2v_inst9.data_to_send_10_0_0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst9.fsm_state_RNISRGO_0_LC_13_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000100"
        )
    port map (
            in0 => \N__26903\,
            in1 => \N__23462\,
            in2 => \N__27206\,
            in3 => \N__28066\,
            lcout => \b2v_inst9.N_740\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst9.fsm_state_RNI44HO_0_LC_13_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010100"
        )
    port map (
            in0 => \N__26902\,
            in1 => \N__23435\,
            in2 => \N__25483\,
            in3 => \N__27203\,
            lcout => \b2v_inst9.N_741\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.energia_temp_0_LC_13_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23405\,
            lcout => b2v_inst_energia_temp_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34442\,
            ce => \N__26180\,
            sr => \N__38099\
        );

    \b2v_inst.energia_temp_1_LC_13_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23371\,
            lcout => b2v_inst_energia_temp_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34442\,
            ce => \N__26180\,
            sr => \N__38099\
        );

    \b2v_inst.energia_temp_13_LC_13_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23333\,
            lcout => b2v_inst_energia_temp_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34442\,
            ce => \N__26180\,
            sr => \N__38099\
        );

    \b2v_inst.energia_temp_2_LC_13_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23681\,
            lcout => b2v_inst_energia_temp_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34442\,
            ce => \N__26180\,
            sr => \N__38099\
        );

    \b2v_inst.energia_temp_3_LC_13_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23654\,
            lcout => b2v_inst_energia_temp_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34442\,
            ce => \N__26180\,
            sr => \N__38099\
        );

    \b2v_inst.data_a_escribir_RNI704E1_5_LC_13_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__37681\,
            in1 => \N__24773\,
            in2 => \N__37626\,
            in3 => \N__37465\,
            lcout => \N_546_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_energia_cry_c_0_LC_13_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39369\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_13_16_0_\,
            carryout => \b2v_inst.dir_energia_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_energia_RNO_0_1_LC_13_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38707\,
            in2 => \_gnd_net_\,
            in3 => \N__23591\,
            lcout => \b2v_inst.dir_energia_s_1\,
            ltout => OPEN,
            carryin => \b2v_inst.dir_energia_cry_0\,
            carryout => \b2v_inst.dir_energia_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_energia_RNO_0_2_LC_13_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36154\,
            in2 => \_gnd_net_\,
            in3 => \N__23573\,
            lcout => \b2v_inst.dir_energia_s_2\,
            ltout => OPEN,
            carryin => \b2v_inst.dir_energia_cry_1\,
            carryout => \b2v_inst.dir_energia_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_energia_RNO_0_3_LC_13_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36463\,
            in2 => \_gnd_net_\,
            in3 => \N__23558\,
            lcout => \b2v_inst.dir_energia_s_3\,
            ltout => OPEN,
            carryin => \b2v_inst.dir_energia_cry_2\,
            carryout => \b2v_inst.dir_energia_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_energia_RNO_0_4_LC_13_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36246\,
            in2 => \_gnd_net_\,
            in3 => \N__23537\,
            lcout => \b2v_inst.dir_energia_s_4\,
            ltout => OPEN,
            carryin => \b2v_inst.dir_energia_cry_3\,
            carryout => \b2v_inst.dir_energia_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_energia_RNO_0_5_LC_13_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35584\,
            in2 => \_gnd_net_\,
            in3 => \N__23522\,
            lcout => \b2v_inst.dir_energia_s_5\,
            ltout => OPEN,
            carryin => \b2v_inst.dir_energia_cry_4\,
            carryout => \b2v_inst.dir_energia_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_energia_RNO_0_6_LC_13_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38422\,
            in2 => \_gnd_net_\,
            in3 => \N__24044\,
            lcout => \b2v_inst.dir_energia_s_6\,
            ltout => OPEN,
            carryin => \b2v_inst.dir_energia_cry_5\,
            carryout => \b2v_inst.dir_energia_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_energia_RNO_0_7_LC_13_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38917\,
            in2 => \_gnd_net_\,
            in3 => \N__24029\,
            lcout => \b2v_inst.dir_energia_s_7\,
            ltout => OPEN,
            carryin => \b2v_inst.dir_energia_cry_6\,
            carryout => \b2v_inst.dir_energia_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_energia_RNO_0_8_LC_13_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39139\,
            in2 => \_gnd_net_\,
            in3 => \N__24014\,
            lcout => \b2v_inst.dir_energia_s_8\,
            ltout => OPEN,
            carryin => \bfn_13_17_0_\,
            carryout => \b2v_inst.dir_energia_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_energia_RNO_0_9_LC_13_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35823\,
            in2 => \_gnd_net_\,
            in3 => \N__23999\,
            lcout => \b2v_inst.dir_energia_s_9\,
            ltout => OPEN,
            carryin => \b2v_inst.dir_energia_cry_8\,
            carryout => \b2v_inst.dir_energia_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_energia_RNO_0_10_LC_13_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36787\,
            in2 => \_gnd_net_\,
            in3 => \N__23981\,
            lcout => \b2v_inst.dir_energia_s_10\,
            ltout => OPEN,
            carryin => \b2v_inst.dir_energia_cry_9\,
            carryout => \b2v_inst.dir_energia_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_energia_11_LC_13_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101001101011100"
        )
    port map (
            in0 => \N__23978\,
            in1 => \N__23818\,
            in2 => \N__23882\,
            in3 => \N__23828\,
            lcout => \b2v_inst.dir_energiaZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34467\,
            ce => \N__23804\,
            sr => \N__38114\
        );

    \b2v_inst.indice_RNI8UI51_10_LC_14_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__23774\,
            in1 => \N__36096\,
            in2 => \N__36726\,
            in3 => \N__38641\,
            lcout => \b2v_inst.un9_indice_0_a2_5_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.cuenta_10_LC_14_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__25953\,
            in1 => \N__24281\,
            in2 => \_gnd_net_\,
            in3 => \N__23726\,
            lcout => \b2v_inst.cuentaZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34443\,
            ce => \N__24180\,
            sr => \N__38100\
        );

    \b2v_inst.cuenta_5_LC_14_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__25954\,
            in1 => \N__24280\,
            in2 => \_gnd_net_\,
            in3 => \N__24230\,
            lcout => \b2v_inst.cuentaZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34432\,
            ce => \N__24179\,
            sr => \N__38091\
        );

    \b2v_inst9.data_to_send_esr_1_LC_14_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__24623\,
            in1 => \N__24311\,
            in2 => \_gnd_net_\,
            in3 => \N__24614\,
            lcout => \b2v_inst9.data_to_sendZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34422\,
            ce => \N__24591\,
            sr => \N__38086\
        );

    \b2v_inst9.data_to_send_esr_4_LC_14_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111101010"
        )
    port map (
            in0 => \N__24119\,
            in1 => \N__25640\,
            in2 => \N__33341\,
            in3 => \N__24137\,
            lcout => \b2v_inst9.data_to_sendZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34422\,
            ce => \N__24591\,
            sr => \N__38086\
        );

    \b2v_inst9.data_to_send_esr_RNO_1_4_LC_14_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__24521\,
            in1 => \N__32630\,
            in2 => \N__24488\,
            in3 => \N__24835\,
            lcout => \b2v_inst9.data_to_send_10_0_0_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst9.data_to_send_esr_RNO_1_5_LC_14_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__24487\,
            in1 => \N__24522\,
            in2 => \N__32600\,
            in3 => \N__24791\,
            lcout => \b2v_inst9.data_to_send_10_0_0_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst9.data_to_send_esr_RNO_2_0_LC_14_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__25632\,
            in1 => \N__24513\,
            in2 => \N__34966\,
            in3 => \N__24425\,
            lcout => \b2v_inst9.data_to_send_10_0_0_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst9.fsm_state_RNI7PQ71_0_LC_14_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__26900\,
            in1 => \N__24104\,
            in2 => \N__27204\,
            in3 => \N__26067\,
            lcout => \b2v_inst9.N_583\,
            ltout => \b2v_inst9.N_583_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst9.fsm_state_RNIQAU12_0_LC_14_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000111"
        )
    port map (
            in0 => \N__30473\,
            in1 => \N__27196\,
            in2 => \N__24092\,
            in3 => \N__26901\,
            lcout => OPEN,
            ltout => \b2v_inst9.un2_n_fsm_state_0_sqmuxa_2_0_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst9.fsm_state_RNI2D372_0_LC_14_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__24089\,
            in1 => \_gnd_net_\,
            in2 => \N__24059\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst9.un2_n_fsm_state_0_sqmuxa_2_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst9.data_to_send_esr_RNO_0_6_LC_14_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__24514\,
            in1 => \N__30376\,
            in2 => \N__24344\,
            in3 => \N__24764\,
            lcout => \b2v_inst9.data_to_send_10_0_0_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst9.data_to_send_esr_RNO_0_7_LC_14_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__30377\,
            in1 => \N__35493\,
            in2 => \N__25639\,
            in3 => \N__24343\,
            lcout => OPEN,
            ltout => \b2v_inst9.data_to_send_10_0_0_0_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst9.data_to_send_esr_7_LC_14_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101011110000"
        )
    port map (
            in0 => \N__24515\,
            in1 => \_gnd_net_\,
            in2 => \N__24347\,
            in3 => \N__24728\,
            lcout => \b2v_inst9.data_to_sendZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34404\,
            ce => \N__24592\,
            sr => \N__38087\
        );

    \b2v_inst9.data_to_send_esr_0_LC_14_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__24332\,
            in1 => \N__24326\,
            in2 => \_gnd_net_\,
            in3 => \N__24287\,
            lcout => \b2v_inst9.data_to_sendZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34404\,
            ce => \N__24592\,
            sr => \N__38087\
        );

    \b2v_inst9.fsm_state_RNIONGO_0_LC_14_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000100"
        )
    port map (
            in0 => \N__26899\,
            in1 => \N__26060\,
            in2 => \N__27205\,
            in3 => \N__25419\,
            lcout => \b2v_inst9.N_738\,
            ltout => \b2v_inst9.N_738_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst9.data_to_send_esr_RNO_2_1_LC_14_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__34825\,
            in1 => \N__25628\,
            in2 => \N__24314\,
            in3 => \N__24389\,
            lcout => \b2v_inst9.data_to_send_10_0_0_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_14_LC_14_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101010101010"
        )
    port map (
            in0 => \N__24662\,
            in1 => \_gnd_net_\,
            in2 => \N__30411\,
            in3 => \N__25816\,
            lcout => b2v_inst_state_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34412\,
            ce => 'H',
            sr => \N__38092\
        );

    \b2v_inst9.fsm_state_RNIP6JC_0_LC_14_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27146\,
            in2 => \_gnd_net_\,
            in3 => \N__26881\,
            lcout => \N_478\,
            ltout => \N_478_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst9.data_to_send_esr_RNO_0_0_LC_14_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__24302\,
            in1 => \N__33380\,
            in2 => \N__24290\,
            in3 => \N__25774\,
            lcout => \b2v_inst9.data_to_send_10_0_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst9.fsm_state_RNI07UL_0_LC_14_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000010"
        )
    port map (
            in0 => \N__24661\,
            in1 => \N__26882\,
            in2 => \N__27182\,
            in3 => \N__25815\,
            lcout => \b2v_inst9.N_832\,
            ltout => \b2v_inst9.N_832_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst9.data_to_send_esr_RNO_0_1_LC_14_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__32853\,
            in1 => \N__24602\,
            in2 => \N__24626\,
            in3 => \N__30371\,
            lcout => \b2v_inst9.data_to_send_10_0_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst9.data_to_send_esr_RNO_1_1_LC_14_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__24549\,
            in1 => \N__26225\,
            in2 => \N__24476\,
            in3 => \N__34874\,
            lcout => \b2v_inst9.data_to_send_10_0_0_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst9.data_to_send_esr_RNO_2_2_LC_14_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__24523\,
            in1 => \N__25624\,
            in2 => \N__33131\,
            in3 => \N__24907\,
            lcout => OPEN,
            ltout => \b2v_inst9.data_to_send_10_0_0_2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst9.data_to_send_esr_2_LC_14_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24530\,
            in2 => \N__24605\,
            in3 => \N__25748\,
            lcout => \b2v_inst9.data_to_sendZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34423\,
            ce => \N__24593\,
            sr => \N__38101\
        );

    \b2v_inst9.data_to_send_esr_RNO_1_2_LC_14_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__24466\,
            in1 => \N__24550\,
            in2 => \N__25145\,
            in3 => \N__32660\,
            lcout => \b2v_inst9.data_to_send_10_0_0_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst9.data_to_send_esr_RNO_1_3_LC_14_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__24524\,
            in1 => \N__34556\,
            in2 => \N__24477\,
            in3 => \N__24880\,
            lcout => \b2v_inst9.data_to_send_10_0_0_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.pix_data_reg_RNIH87G_0_LC_14_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25577\,
            in2 => \N__24421\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst.un14_data_ram_energia_o_axb_0\,
            ltout => OPEN,
            carryin => \bfn_14_14_0_\,
            carryout => \b2v_inst.un14_data_ram_energia_o_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un14_data_ram_energia_o_cry_0_c_RNIEI4M_LC_14_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25571\,
            in2 => \N__24388\,
            in3 => \N__24356\,
            lcout => \b2v_inst.un14_data_ram_energia_o_cry_0_c_RNIEI4MZ0\,
            ltout => OPEN,
            carryin => \b2v_inst.un14_data_ram_energia_o_cry_0\,
            carryout => \b2v_inst.un14_data_ram_energia_o_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un14_data_ram_energia_o_cry_1_c_RNIHM5M_LC_14_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26300\,
            in2 => \N__24908\,
            in3 => \N__24884\,
            lcout => \b2v_inst.un14_data_ram_energia_o_cry_1_c_RNIHM5MZ0\,
            ltout => OPEN,
            carryin => \b2v_inst.un14_data_ram_energia_o_cry_1\,
            carryout => \b2v_inst.un14_data_ram_energia_o_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un14_data_ram_energia_o_cry_2_c_RNIKQ6M_LC_14_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30260\,
            in2 => \N__24881\,
            in3 => \N__24857\,
            lcout => \b2v_inst.un14_data_ram_energia_o_cry_2_c_RNIKQ6MZ0\,
            ltout => OPEN,
            carryin => \b2v_inst.un14_data_ram_energia_o_cry_2\,
            carryout => \b2v_inst.un14_data_ram_energia_o_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un14_data_ram_energia_o_cry_3_c_RNINU7M_LC_14_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24854\,
            in2 => \N__24836\,
            in3 => \N__24794\,
            lcout => \b2v_inst.un14_data_ram_energia_o_cry_3_c_RNINU7MZ0\,
            ltout => OPEN,
            carryin => \b2v_inst.un14_data_ram_energia_o_cry_3\,
            carryout => \b2v_inst.un14_data_ram_energia_o_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un14_data_ram_energia_o_cry_4_c_RNIQ29M_LC_14_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24790\,
            in2 => \N__26294\,
            in3 => \N__24767\,
            lcout => \b2v_inst.un14_data_ram_energia_o_cry_4_c_RNIQ29MZ0\,
            ltout => OPEN,
            carryin => \b2v_inst.un14_data_ram_energia_o_cry_4\,
            carryout => \b2v_inst.un14_data_ram_energia_o_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un14_data_ram_energia_o_cry_5_c_RNIT6AM_LC_14_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26285\,
            in2 => \N__24763\,
            in3 => \N__24731\,
            lcout => \b2v_inst.un14_data_ram_energia_o_cry_5_c_RNIT6AMZ0\,
            ltout => OPEN,
            carryin => \b2v_inst.un14_data_ram_energia_o_cry_5\,
            carryout => \b2v_inst.un14_data_ram_energia_o_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un14_data_ram_energia_o_cry_6_c_RNI0BBM_LC_14_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26279\,
            in2 => \N__24727\,
            in3 => \N__24695\,
            lcout => \b2v_inst.un14_data_ram_energia_o_cry_6_c_RNI0BBMZ0\,
            ltout => OPEN,
            carryin => \b2v_inst.un14_data_ram_energia_o_cry_6\,
            carryout => \b2v_inst.un14_data_ram_energia_o_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un14_data_ram_energia_o_cry_7_c_RNIN84C_LC_14_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24943\,
            in2 => \_gnd_net_\,
            in3 => \N__24680\,
            lcout => \b2v_inst.un14_data_ram_energia_o_cry_7_c_RNIN84CZ0\,
            ltout => OPEN,
            carryin => \bfn_14_15_0_\,
            carryout => \b2v_inst.un14_data_ram_energia_o_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un14_data_ram_energia_o_cry_8_c_RNIPB5C_LC_14_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26221\,
            in2 => \_gnd_net_\,
            in3 => \N__24665\,
            lcout => \b2v_inst.un14_data_ram_energia_o_cry_8_c_RNIPB5CZ0\,
            ltout => OPEN,
            carryin => \b2v_inst.un14_data_ram_energia_o_cry_8\,
            carryout => \b2v_inst.un14_data_ram_energia_o_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un14_data_ram_energia_o_cry_9_c_RNI28GB_LC_14_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25141\,
            in2 => \_gnd_net_\,
            in3 => \N__25112\,
            lcout => \b2v_inst.un14_data_ram_energia_o_cry_9_c_RNI28GBZ0\,
            ltout => OPEN,
            carryin => \b2v_inst.un14_data_ram_energia_o_cry_9\,
            carryout => \b2v_inst.un14_data_ram_energia_o_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un14_data_ram_energia_o_cry_10_c_RNIMOAH_LC_14_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37460\,
            in1 => \N__25105\,
            in2 => \_gnd_net_\,
            in3 => \N__25064\,
            lcout => \SYNTHESIZED_WIRE_13_11\,
            ltout => OPEN,
            carryin => \b2v_inst.un14_data_ram_energia_o_cry_10\,
            carryout => \b2v_inst.un14_data_ram_energia_o_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un14_data_ram_energia_o_cry_11_c_RNIORBH_LC_14_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37459\,
            in1 => \N__25057\,
            in2 => \_gnd_net_\,
            in3 => \N__25016\,
            lcout => \SYNTHESIZED_WIRE_13_12\,
            ltout => OPEN,
            carryin => \b2v_inst.un14_data_ram_energia_o_cry_11\,
            carryout => \b2v_inst.un14_data_ram_energia_o_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un14_data_ram_energia_o_cry_12_c_RNIQUCH_LC_14_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37461\,
            in1 => \N__25009\,
            in2 => \_gnd_net_\,
            in3 => \N__24995\,
            lcout => \SYNTHESIZED_WIRE_13_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.energia_temp_8_LC_14_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24976\,
            lcout => b2v_inst_energia_temp_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34444\,
            ce => \N__26190\,
            sr => \N__38109\
        );

    \b2v_inst.data_a_escribir_RNIRV031_10_LC_14_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__37733\,
            in1 => \N__24932\,
            in2 => \N__33682\,
            in3 => \N__37502\,
            lcout => \N_461_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.reg_ancho_2_5_LC_15_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32124\,
            lcout => \b2v_inst.reg_ancho_2Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34449\,
            ce => \N__32964\,
            sr => \N__38115\
        );

    \b2v_inst.reg_anterior_2_LC_15_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31894\,
            in2 => \_gnd_net_\,
            in3 => \N__32210\,
            lcout => \b2v_inst.reg_anteriorZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34445\,
            ce => \N__31686\,
            sr => \N__38110\
        );

    \b2v_inst.reg_anterior_3_LC_15_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__31895\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32285\,
            lcout => \b2v_inst.reg_anteriorZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34445\,
            ce => \N__31686\,
            sr => \N__38110\
        );

    \b2v_inst.data_a_escribir11_2_c_RNO_LC_15_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__29246\,
            in1 => \N__29988\,
            in2 => \N__27441\,
            in3 => \N__29949\,
            lcout => \b2v_inst.data_a_escribir11_2_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.reg_ancho_2_8_LC_15_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27251\,
            lcout => \b2v_inst.reg_ancho_2Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34433\,
            ce => \N__32930\,
            sr => \N__38105\
        );

    \b2v_inst.data_a_escribir11_4_c_RNO_LC_15_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__27562\,
            in1 => \N__27319\,
            in2 => \N__29909\,
            in3 => \N__27383\,
            lcout => \b2v_inst.data_a_escribir11_4_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.reg_ancho_2_6_LC_15_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31571\,
            lcout => \b2v_inst.reg_ancho_2Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34433\,
            ce => \N__32930\,
            sr => \N__38105\
        );

    \b2v_inst.reg_ancho_2_7_LC_15_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27276\,
            lcout => \b2v_inst.reg_ancho_2Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34433\,
            ce => \N__32930\,
            sr => \N__38105\
        );

    \b2v_inst.data_a_escribir11_0_c_LC_15_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26408\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_8_0_\,
            carryout => \b2v_inst.data_a_escribir11_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir11_1_c_LC_15_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26630\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.data_a_escribir11_0\,
            carryout => \b2v_inst.data_a_escribir11_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir11_2_c_LC_15_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25151\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.data_a_escribir11_1\,
            carryout => \b2v_inst.data_a_escribir11_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir11_3_c_LC_15_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31415\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.data_a_escribir11_2\,
            carryout => \b2v_inst.data_a_escribir11_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir11_4_c_LC_15_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25166\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.data_a_escribir11_3\,
            carryout => \b2v_inst.data_a_escribir11_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir11_5_c_LC_15_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29648\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.data_a_escribir11_4\,
            carryout => \b2v_inst.data_a_escribir11_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir11_6_c_LC_15_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29801\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.data_a_escribir11_5\,
            carryout => \b2v_inst.data_a_escribir11_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir11_7_c_LC_15_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27296\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.data_a_escribir11_6\,
            carryout => \b2v_inst.data_a_escribir11_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir11_8_c_LC_15_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25388\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_9_0_\,
            carryout => \b2v_inst.data_a_escribir11_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir11_9_c_LC_15_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25157\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.data_a_escribir11_8\,
            carryout => \b2v_inst.data_a_escribir11_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir11_10_c_LC_15_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30050\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.data_a_escribir11_9\,
            carryout => \b2v_inst.data_a_escribir12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir12_THRU_LUT4_0_LC_15_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25160\,
            lcout => \b2v_inst.data_a_escribir12_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir11_9_c_RNO_LC_15_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__29105\,
            in1 => \N__30175\,
            in2 => \N__31529\,
            in3 => \N__29157\,
            lcout => \b2v_inst.data_a_escribir11_9_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir11_8_c_RNO_LC_15_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__28588\,
            in1 => \N__28614\,
            in2 => \N__29840\,
            in3 => \N__32309\,
            lcout => \b2v_inst.data_a_escribir11_8_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_3_RNI68I31_10_LC_15_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__25382\,
            in1 => \N__25367\,
            in2 => \N__25286\,
            in3 => \N__25268\,
            lcout => \b2v_inst.addr_ram_iv_i_1_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.eventos_0_LC_15_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1011",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26590\,
            in2 => \_gnd_net_\,
            in3 => \N__25187\,
            lcout => \b2v_inst.eventosZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_15_10_0_\,
            carryout => \b2v_inst.eventos_cry_0\,
            clk => \N__34405\,
            ce => \N__26651\,
            sr => \N__38080\
        );

    \b2v_inst.eventos_1_LC_15_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26569\,
            in2 => \_gnd_net_\,
            in3 => \N__25184\,
            lcout => \b2v_inst.eventosZ0Z_1\,
            ltout => OPEN,
            carryin => \b2v_inst.eventos_cry_0\,
            carryout => \b2v_inst.eventos_cry_1\,
            clk => \N__34405\,
            ce => \N__26651\,
            sr => \N__38080\
        );

    \b2v_inst.eventos_2_LC_15_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31195\,
            in2 => \_gnd_net_\,
            in3 => \N__25181\,
            lcout => \b2v_inst.eventosZ0Z_2\,
            ltout => OPEN,
            carryin => \b2v_inst.eventos_cry_1\,
            carryout => \b2v_inst.eventos_cry_2\,
            clk => \N__34405\,
            ce => \N__26651\,
            sr => \N__38080\
        );

    \b2v_inst.eventos_3_LC_15_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29863\,
            in2 => \_gnd_net_\,
            in3 => \N__25178\,
            lcout => \b2v_inst.eventosZ0Z_3\,
            ltout => OPEN,
            carryin => \b2v_inst.eventos_cry_2\,
            carryout => \b2v_inst.eventos_cry_3\,
            clk => \N__34405\,
            ce => \N__26651\,
            sr => \N__38080\
        );

    \b2v_inst.eventos_4_LC_15_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26617\,
            in2 => \_gnd_net_\,
            in3 => \N__25175\,
            lcout => \b2v_inst.eventosZ0Z_4\,
            ltout => OPEN,
            carryin => \b2v_inst.eventos_cry_3\,
            carryout => \b2v_inst.eventos_cry_4\,
            clk => \N__34405\,
            ce => \N__26651\,
            sr => \N__38080\
        );

    \b2v_inst.eventos_5_LC_15_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27520\,
            in2 => \_gnd_net_\,
            in3 => \N__25172\,
            lcout => \b2v_inst.eventosZ0Z_5\,
            ltout => OPEN,
            carryin => \b2v_inst.eventos_cry_4\,
            carryout => \b2v_inst.eventos_cry_5\,
            clk => \N__34405\,
            ce => \N__26651\,
            sr => \N__38080\
        );

    \b2v_inst.eventos_6_LC_15_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26674\,
            in2 => \_gnd_net_\,
            in3 => \N__25169\,
            lcout => \b2v_inst.eventosZ0Z_6\,
            ltout => OPEN,
            carryin => \b2v_inst.eventos_cry_5\,
            carryout => \b2v_inst.eventos_cry_6\,
            clk => \N__34405\,
            ce => \N__26651\,
            sr => \N__38080\
        );

    \b2v_inst.eventos_7_LC_15_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28480\,
            in2 => \_gnd_net_\,
            in3 => \N__25565\,
            lcout => \b2v_inst.eventosZ0Z_7\,
            ltout => OPEN,
            carryin => \b2v_inst.eventos_cry_6\,
            carryout => \b2v_inst.eventos_cry_7\,
            clk => \N__34405\,
            ce => \N__26651\,
            sr => \N__38080\
        );

    \b2v_inst.eventos_8_LC_15_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30034\,
            in2 => \_gnd_net_\,
            in3 => \N__25562\,
            lcout => \b2v_inst.eventosZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_15_11_0_\,
            carryout => \b2v_inst.eventos_cry_8\,
            clk => \N__34394\,
            ce => \N__26647\,
            sr => \N__38093\
        );

    \b2v_inst.eventos_9_LC_15_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30109\,
            in2 => \_gnd_net_\,
            in3 => \N__25559\,
            lcout => \b2v_inst.eventosZ0Z_9\,
            ltout => OPEN,
            carryin => \b2v_inst.eventos_cry_8\,
            carryout => \b2v_inst.eventos_cry_9\,
            clk => \N__34394\,
            ce => \N__26647\,
            sr => \N__38093\
        );

    \b2v_inst.eventos_10_LC_15_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26552\,
            in2 => \_gnd_net_\,
            in3 => \N__25556\,
            lcout => \b2v_inst.eventosZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34394\,
            ce => \N__26647\,
            sr => \N__38093\
        );

    \b2v_inst.state_RNO_1_31_LC_15_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__25417\,
            in1 => \N__25470\,
            in2 => \N__34746\,
            in3 => \N__28064\,
            lcout => OPEN,
            ltout => \b2v_inst.state_ns_a3_i_0_a2_4_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_31_LC_15_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001111111"
        )
    port map (
            in0 => \N__25784\,
            in1 => \N__25553\,
            in2 => \N__25541\,
            in3 => \N__28016\,
            lcout => \b2v_inst.stateZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34406\,
            ce => 'H',
            sr => \N__38102\
        );

    \b2v_inst.state_RNO_6_31_LC_15_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__25469\,
            in1 => \N__25416\,
            in2 => \N__25731\,
            in3 => \N__25814\,
            lcout => \b2v_inst.state_ns_a3_i_0_a2_1_4_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_1_LC_15_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111110100000"
        )
    port map (
            in0 => \N__25418\,
            in1 => \_gnd_net_\,
            in2 => \N__30412\,
            in3 => \N__26061\,
            lcout => b2v_inst_state_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34406\,
            ce => 'H',
            sr => \N__38102\
        );

    \b2v_inst.state_12_LC_15_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__25722\,
            in1 => \N__30379\,
            in2 => \_gnd_net_\,
            in3 => \N__25691\,
            lcout => b2v_inst_state_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34406\,
            ce => 'H',
            sr => \N__38102\
        );

    \b2v_inst.state_2_LC_15_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__30383\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28065\,
            lcout => b2v_inst_state_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34406\,
            ce => 'H',
            sr => \N__38102\
        );

    \b2v_inst.state_11_LC_15_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__25721\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30378\,
            lcout => \b2v_inst.stateZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34406\,
            ce => 'H',
            sr => \N__38102\
        );

    \b2v_inst.state_RNO_3_31_LC_15_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__25724\,
            in1 => \N__33180\,
            in2 => \N__25935\,
            in3 => \N__25817\,
            lcout => \b2v_inst.state_ns_a3_i_0_a2_6_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst9.fsm_state_RNO_0_1_LC_15_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000110011"
        )
    port map (
            in0 => \N__30472\,
            in1 => \N__27162\,
            in2 => \_gnd_net_\,
            in3 => \N__26884\,
            lcout => OPEN,
            ltout => \b2v_inst9.fsm_state_ns_i_0_i_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst9.fsm_state_1_LC_15_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010000001100"
        )
    port map (
            in0 => \N__26885\,
            in1 => \N__27840\,
            in2 => \N__25778\,
            in3 => \N__27101\,
            lcout => \b2v_inst9.fsm_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34413\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst9.data_to_send_esr_RNO_0_2_LC_15_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__25775\,
            in1 => \N__33648\,
            in2 => \N__25763\,
            in3 => \N__30375\,
            lcout => \b2v_inst9.data_to_send_10_0_0_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst9.fsm_state_RNIS2UL_0_LC_15_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000100"
        )
    port map (
            in0 => \N__26883\,
            in1 => \N__25723\,
            in2 => \N__27188\,
            in3 => \N__25687\,
            lcout => \b2v_inst9.N_739\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.pix_data_reg_0_LC_15_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26690\,
            lcout => \b2v_inst.pix_data_regZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34424\,
            ce => \N__30244\,
            sr => \N__38111\
        );

    \b2v_inst.pix_data_reg_1_LC_15_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26999\,
            lcout => \b2v_inst.pix_data_regZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34424\,
            ce => \N__30244\,
            sr => \N__38111\
        );

    \b2v_inst.pix_data_reg_2_LC_15_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26966\,
            lcout => \b2v_inst.pix_data_regZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34424\,
            ce => \N__30244\,
            sr => \N__38111\
        );

    \b2v_inst.pix_data_reg_5_LC_15_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28802\,
            lcout => \b2v_inst.pix_data_regZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34424\,
            ce => \N__30244\,
            sr => \N__38111\
        );

    \b2v_inst.pix_data_reg_6_LC_15_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28841\,
            lcout => \b2v_inst.pix_data_regZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34424\,
            ce => \N__30244\,
            sr => \N__38111\
        );

    \b2v_inst.pix_data_reg_7_LC_15_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__28853\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst.pix_data_regZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34424\,
            ce => \N__30244\,
            sr => \N__38111\
        );

    \b2v_inst9.fsm_state_0_LC_15_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__26921\,
            in1 => \N__26273\,
            in2 => \N__27845\,
            in3 => \N__27097\,
            lcout => \b2v_inst9.fsm_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34434\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.energia_temp_9_LC_15_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26260\,
            lcout => b2v_inst_energia_temp_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34450\,
            ce => \N__26205\,
            sr => \N__38128\
        );

    \b2v_inst9.txd_reg_LC_15_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110010111011"
        )
    port map (
            in0 => \N__26111\,
            in1 => \N__27192\,
            in2 => \_gnd_net_\,
            in3 => \N__26898\,
            lcout => uart_tx_o_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34457\,
            ce => 'H',
            sr => \N__38135\
        );

    \b2v_inst.reg_ancho_2_0_LC_16_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__27486\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst.reg_ancho_2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34451\,
            ce => \N__32958\,
            sr => \N__38129\
        );

    \b2v_inst.reg_ancho_1_0_LC_16_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26522\,
            in2 => \_gnd_net_\,
            in3 => \N__27479\,
            lcout => \b2v_inst.reg_ancho_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34446\,
            ce => \N__26462\,
            sr => \N__38123\
        );

    \b2v_inst.reg_ancho_1_1_LC_16_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__26524\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31394\,
            lcout => \b2v_inst.reg_ancho_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34446\,
            ce => \N__26462\,
            sr => \N__38123\
        );

    \b2v_inst.reg_ancho_1_10_LC_16_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26523\,
            in2 => \_gnd_net_\,
            in3 => \N__31781\,
            lcout => \b2v_inst.reg_ancho_1Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34446\,
            ce => \N__26462\,
            sr => \N__38123\
        );

    \b2v_inst.reg_ancho_1_2_LC_16_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__26525\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32204\,
            lcout => \b2v_inst.reg_ancho_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34446\,
            ce => \N__26462\,
            sr => \N__38123\
        );

    \b2v_inst.reg_ancho_1_3_LC_16_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26526\,
            in2 => \_gnd_net_\,
            in3 => \N__32282\,
            lcout => \b2v_inst.reg_ancho_1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34446\,
            ce => \N__26462\,
            sr => \N__38123\
        );

    \b2v_inst.reg_ancho_1_4_LC_16_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__26527\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33062\,
            lcout => \b2v_inst.reg_ancho_1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34446\,
            ce => \N__26462\,
            sr => \N__38123\
        );

    \b2v_inst.reg_ancho_1_6_LC_16_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__26528\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31570\,
            lcout => \b2v_inst.reg_ancho_1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34446\,
            ce => \N__26462\,
            sr => \N__38123\
        );

    \b2v_inst.encontrar_maximo_un2_valor_max1_cry_0_c_inv_LC_16_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27430\,
            in2 => \N__26327\,
            in3 => \N__29045\,
            lcout => \b2v_inst.reg_ancho_1_i_0\,
            ltout => OPEN,
            carryin => \bfn_16_6_0_\,
            carryout => \b2v_inst.un2_valor_max1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_un2_valor_max1_cry_1_c_inv_LC_16_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31346\,
            in2 => \N__26318\,
            in3 => \N__28971\,
            lcout => \b2v_inst.reg_ancho_1_i_1\,
            ltout => OPEN,
            carryin => \b2v_inst.un2_valor_max1_cry_0\,
            carryout => \b2v_inst.un2_valor_max1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_un2_valor_max1_cry_2_c_inv_LC_16_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31299\,
            in2 => \N__26309\,
            in3 => \N__31223\,
            lcout => \b2v_inst.reg_ancho_1_i_2\,
            ltout => OPEN,
            carryin => \b2v_inst.un2_valor_max1_cry_1\,
            carryout => \b2v_inst.un2_valor_max1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_un2_valor_max1_cry_3_c_inv_LC_16_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32448\,
            in2 => \N__26399\,
            in3 => \N__31010\,
            lcout => \b2v_inst.reg_ancho_1_i_3\,
            ltout => OPEN,
            carryin => \b2v_inst.un2_valor_max1_cry_2\,
            carryout => \b2v_inst.un2_valor_max1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_un2_valor_max1_cry_4_c_inv_LC_16_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33015\,
            in2 => \N__26390\,
            in3 => \N__29615\,
            lcout => \b2v_inst.reg_ancho_1_i_4\,
            ltout => OPEN,
            carryin => \b2v_inst.un2_valor_max1_cry_3\,
            carryout => \b2v_inst.un2_valor_max1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_un2_valor_max1_cry_5_c_inv_LC_16_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27370\,
            in2 => \N__26381\,
            in3 => \N__29551\,
            lcout => \b2v_inst.reg_ancho_1_i_5\,
            ltout => OPEN,
            carryin => \b2v_inst.un2_valor_max1_cry_4\,
            carryout => \b2v_inst.un2_valor_max1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_un2_valor_max1_cry_6_c_inv_LC_16_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27320\,
            in2 => \N__26372\,
            in3 => \N__29465\,
            lcout => \b2v_inst.reg_ancho_1_i_6\,
            ltout => OPEN,
            carryin => \b2v_inst.un2_valor_max1_cry_5\,
            carryout => \b2v_inst.un2_valor_max1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_un2_valor_max1_cry_7_c_inv_LC_16_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27575\,
            in2 => \N__26363\,
            in3 => \N__29386\,
            lcout => \b2v_inst.reg_ancho_1_i_7\,
            ltout => OPEN,
            carryin => \b2v_inst.un2_valor_max1_cry_6\,
            carryout => \b2v_inst.un2_valor_max1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_un2_valor_max1_cry_8_c_inv_LC_16_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__29948\,
            in1 => \N__29899\,
            in2 => \N__26354\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst.reg_ancho_1_i_8\,
            ltout => OPEN,
            carryin => \bfn_16_7_0_\,
            carryout => \b2v_inst.un2_valor_max1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_un2_valor_max1_cry_9_c_inv_LC_16_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29725\,
            in2 => \N__26345\,
            in3 => \N__29987\,
            lcout => \b2v_inst.reg_ancho_1_i_9\,
            ltout => OPEN,
            carryin => \b2v_inst.un2_valor_max1_cry_8\,
            carryout => \b2v_inst.un2_valor_max1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_un2_valor_max1_cry_10_c_inv_LC_16_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31487\,
            in2 => \N__26336\,
            in3 => \N__29245\,
            lcout => \b2v_inst.reg_ancho_1_i_10\,
            ltout => OPEN,
            carryin => \b2v_inst.un2_valor_max1_cry_9\,
            carryout => \b2v_inst.un2_valor_max1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un2_valor_max1_THRU_LUT4_0_LC_16_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26531\,
            lcout => \b2v_inst.un2_valor_max1_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.reg_ancho_2_9_LC_16_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31994\,
            lcout => \b2v_inst.reg_ancho_2Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34425\,
            ce => \N__32963\,
            sr => \N__38112\
        );

    \b2v_inst.reg_ancho_1_7_LC_16_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__26519\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27283\,
            lcout => \b2v_inst.reg_ancho_1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34414\,
            ce => \N__26458\,
            sr => \N__38106\
        );

    \b2v_inst.reg_ancho_1_8_LC_16_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26520\,
            in2 => \_gnd_net_\,
            in3 => \N__27249\,
            lcout => \b2v_inst.reg_ancho_1Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34414\,
            ce => \N__26458\,
            sr => \N__38106\
        );

    \b2v_inst.reg_ancho_1_9_LC_16_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__31993\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26521\,
            lcout => \b2v_inst.reg_ancho_1Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34414\,
            ce => \N__26458\,
            sr => \N__38106\
        );

    \b2v_inst.reg_ancho_1_5_LC_16_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26518\,
            in2 => \_gnd_net_\,
            in3 => \N__32132\,
            lcout => \b2v_inst.reg_ancho_1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34414\,
            ce => \N__26458\,
            sr => \N__38106\
        );

    \b2v_inst.reg_anterior_0_LC_16_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__27488\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31831\,
            lcout => \b2v_inst.reg_anteriorZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34407\,
            ce => \N__31671\,
            sr => \N__38103\
        );

    \b2v_inst.reg_anterior_8_LC_16_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31833\,
            in2 => \_gnd_net_\,
            in3 => \N__27248\,
            lcout => \b2v_inst.reg_anteriorZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34407\,
            ce => \N__31671\,
            sr => \N__38103\
        );

    \b2v_inst.reg_anterior_7_LC_16_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31832\,
            in2 => \_gnd_net_\,
            in3 => \N__27284\,
            lcout => \b2v_inst.reg_anteriorZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34407\,
            ce => \N__31671\,
            sr => \N__38103\
        );

    \b2v_inst.data_a_escribir11_0_c_RNO_LC_16_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__31241\,
            in1 => \N__28982\,
            in2 => \N__31042\,
            in3 => \N__29060\,
            lcout => \b2v_inst.data_a_escribir11_0_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_2_0_LC_16_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111101011111"
        )
    port map (
            in0 => \N__29061\,
            in1 => \N__27449\,
            in2 => \N__30910\,
            in3 => \N__32540\,
            lcout => OPEN,
            ltout => \b2v_inst.data_a_escribir_RNO_2Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_1_0_LC_16_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100001111"
        )
    port map (
            in0 => \N__26591\,
            in1 => \N__30860\,
            in2 => \N__26579\,
            in3 => \N__31110\,
            lcout => OPEN,
            ltout => \b2v_inst.un1_reg_anterior_0_i_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_0_LC_16_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001101101011010"
        )
    port map (
            in0 => \N__31112\,
            in1 => \N__27539\,
            in2 => \N__26576\,
            in3 => \N__30625\,
            lcout => b2v_inst_data_a_escribir_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34395\,
            ce => \N__30553\,
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_2_1_LC_16_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111101011111"
        )
    port map (
            in0 => \N__28983\,
            in1 => \N__31350\,
            in2 => \N__30911\,
            in3 => \N__32541\,
            lcout => OPEN,
            ltout => \b2v_inst.data_a_escribir_RNO_2Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_1_1_LC_16_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100001111"
        )
    port map (
            in0 => \N__26573\,
            in1 => \N__30861\,
            in2 => \N__26558\,
            in3 => \N__31111\,
            lcout => OPEN,
            ltout => \b2v_inst.un1_reg_anterior_0_i_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_1_LC_16_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001101101011010"
        )
    port map (
            in0 => \N__31113\,
            in1 => \N__27533\,
            in2 => \N__26555\,
            in3 => \N__30626\,
            lcout => b2v_inst_data_a_escribir_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34395\,
            ce => \N__30553\,
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_2_10_LC_16_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__29258\,
            in1 => \N__31490\,
            in2 => \_gnd_net_\,
            in3 => \N__32537\,
            lcout => \b2v_inst.N_269\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_3_10_LC_16_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26551\,
            in2 => \N__30982\,
            in3 => \N__31114\,
            lcout => OPEN,
            ltout => \b2v_inst.un1_reg_anterior_iv_0_0_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_1_10_LC_16_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110001"
        )
    port map (
            in0 => \N__31116\,
            in1 => \N__26540\,
            in2 => \N__26534\,
            in3 => \N__30607\,
            lcout => \b2v_inst.un1_reg_anterior_iv_0_1_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_3_6_LC_16_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111100001111"
        )
    port map (
            in0 => \N__26678\,
            in1 => \_gnd_net_\,
            in2 => \N__30981\,
            in3 => \N__31115\,
            lcout => OPEN,
            ltout => \b2v_inst.un1_reg_anterior_iv_0_0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_1_6_LC_16_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110001"
        )
    port map (
            in0 => \N__31117\,
            in1 => \N__26657\,
            in2 => \N__26660\,
            in3 => \N__30606\,
            lcout => \b2v_inst.un1_reg_anterior_iv_0_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_2_6_LC_16_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32536\,
            in1 => \N__27350\,
            in2 => \_gnd_net_\,
            in3 => \N__29486\,
            lcout => \b2v_inst.N_272\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNILIBG_20_LC_16_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__31118\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30946\,
            lcout => \b2v_inst.data_a_escribir_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_3_LC_16_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001111001110"
        )
    port map (
            in0 => \N__30608\,
            in1 => \N__31119\,
            in2 => \N__29120\,
            in3 => \N__29852\,
            lcout => b2v_inst_data_a_escribir_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34391\,
            ce => \N__30556\,
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir11_1_c_RNO_LC_16_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__29552\,
            in1 => \N__29474\,
            in2 => \N__29395\,
            in3 => \N__29633\,
            lcout => \b2v_inst.data_a_escribir11_1_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_3_4_LC_16_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111011101"
        )
    port map (
            in0 => \N__30945\,
            in1 => \N__31164\,
            in2 => \_gnd_net_\,
            in3 => \N__26618\,
            lcout => OPEN,
            ltout => \b2v_inst.un1_reg_anterior_iv_0_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_1_4_LC_16_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110001"
        )
    port map (
            in0 => \N__31165\,
            in1 => \N__26597\,
            in2 => \N__26603\,
            in3 => \N__30612\,
            lcout => OPEN,
            ltout => \b2v_inst.un1_reg_anterior_iv_0_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_4_LC_16_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100001101"
        )
    port map (
            in0 => \N__30614\,
            in1 => \N__31167\,
            in2 => \N__26600\,
            in3 => \N__26819\,
            lcout => b2v_inst_data_a_escribir_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34396\,
            ce => \N__30552\,
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_2_4_LC_16_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__33020\,
            in1 => \N__29634\,
            in2 => \_gnd_net_\,
            in3 => \N__32539\,
            lcout => \b2v_inst.N_274\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_2_7_LC_16_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111100111111"
        )
    port map (
            in0 => \N__27586\,
            in1 => \N__29390\,
            in2 => \N__30980\,
            in3 => \N__32538\,
            lcout => \b2v_inst.data_a_escribir_RNO_2Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_0_4_LC_16_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30176\,
            in1 => \N__31442\,
            in2 => \_gnd_net_\,
            in3 => \N__32408\,
            lcout => \b2v_inst.N_268\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_10_LC_16_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111101"
        )
    port map (
            in0 => \N__30613\,
            in1 => \N__31166\,
            in2 => \N__32324\,
            in3 => \N__26813\,
            lcout => b2v_inst_data_a_escribir_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34396\,
            ce => \N__30552\,
            sr => \_gnd_net_\
        );

    \b2v_inst4.reg_data_3_LC_16_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26807\,
            lcout => \SYNTHESIZED_WIRE_5_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34408\,
            ce => \N__28783\,
            sr => \N__38113\
        );

    \b2v_inst4.reg_data_4_LC_16_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__26780\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \SYNTHESIZED_WIRE_5_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34408\,
            ce => \N__28783\,
            sr => \N__38113\
        );

    \b2v_inst4.reg_data_6_LC_16_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26762\,
            lcout => \SYNTHESIZED_WIRE_5_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34408\,
            ce => \N__28783\,
            sr => \N__38113\
        );

    \b2v_inst4.reg_data_7_LC_16_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26744\,
            lcout => \SYNTHESIZED_WIRE_5_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34408\,
            ce => \N__28783\,
            sr => \N__38113\
        );

    \b2v_inst4.reg_data_0_LC_16_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26720\,
            lcout => \SYNTHESIZED_WIRE_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34408\,
            ce => \N__28783\,
            sr => \N__38113\
        );

    \b2v_inst.un12_pix_count_intlto7_N_2L1_LC_16_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__26965\,
            in1 => \N__26998\,
            in2 => \N__30277\,
            in3 => \N__26689\,
            lcout => OPEN,
            ltout => \b2v_inst.un12_pix_count_intlto7_N_2LZ0Z1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un12_pix_count_intlto7_LC_16_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011100000000"
        )
    port map (
            in0 => \N__27073\,
            in1 => \N__28840\,
            in2 => \N__27062\,
            in3 => \N__28823\,
            lcout => \b2v_inst.un13_pix_count_int_li_0\,
            ltout => \b2v_inst.un13_pix_count_int_li_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNI3K574_29_LC_16_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27032\,
            in3 => \N__28208\,
            lcout => \b2v_inst.N_654_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst4.reg_data_1_LC_16_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27029\,
            lcout => \SYNTHESIZED_WIRE_5_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34415\,
            ce => \N__28779\,
            sr => \N__38116\
        );

    \b2v_inst4.reg_data_2_LC_16_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26987\,
            lcout => \SYNTHESIZED_WIRE_5_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34415\,
            ce => \N__28779\,
            sr => \N__38116\
        );

    \b2v_inst.state_fast_RNITDD01_19_LC_16_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__34745\,
            in1 => \N__37498\,
            in2 => \N__26954\,
            in3 => \N__33187\,
            lcout => \b2v_inst.N_484\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst9.fsm_state_RNO_0_0_LC_16_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111000000"
        )
    port map (
            in0 => \N__30471\,
            in1 => \N__27191\,
            in2 => \N__26915\,
            in3 => \N__26897\,
            lcout => \b2v_inst9.fsm_state_srsts_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst9.bit_counter_RNIM4971_3_LC_16_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__28693\,
            in1 => \N__28632\,
            in2 => \N__28676\,
            in3 => \N__28707\,
            lcout => \b2v_inst9.N_522\,
            ltout => \b2v_inst9.N_522_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst9.fsm_state_RNIND1P1_0_LC_16_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101111111"
        )
    port map (
            in0 => \N__27844\,
            in1 => \N__27189\,
            in2 => \N__26906\,
            in3 => \N__26874\,
            lcout => \b2v_inst9.fsm_state_RNIND1P1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst9.bit_counter_RNIBIKJ_1_LC_16_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28671\,
            in2 => \_gnd_net_\,
            in3 => \N__28692\,
            lcout => OPEN,
            ltout => \b2v_inst9.N_84_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst9.bit_counter_RNIJOID1_3_LC_16_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__27190\,
            in1 => \N__28633\,
            in2 => \N__27104\,
            in3 => \N__28708\,
            lcout => \b2v_inst9.N_582\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final4_2_cry_0_c_LC_17_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29023\,
            in2 => \N__27434\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_17_5_0_\,
            carryout => \b2v_inst.valor_max_final4_2_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final4_2_cry_1_c_LC_17_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31351\,
            in2 => \N__28951\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.valor_max_final4_2_cry_0\,
            carryout => \b2v_inst.valor_max_final4_2_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final4_2_cry_2_c_LC_17_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31300\,
            in2 => \N__28916\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.valor_max_final4_2_cry_1\,
            carryout => \b2v_inst.valor_max_final4_2_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final4_2_cry_3_c_LC_17_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28882\,
            in2 => \N__32459\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.valor_max_final4_2_cry_2\,
            carryout => \b2v_inst.valor_max_final4_2_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final4_2_cry_4_c_LC_17_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33019\,
            in2 => \N__29591\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.valor_max_final4_2_cry_3\,
            carryout => \b2v_inst.valor_max_final4_2_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final4_2_cry_5_c_LC_17_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29512\,
            in2 => \N__27394\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.valor_max_final4_2_cry_4\,
            carryout => \b2v_inst.valor_max_final4_2_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final4_2_cry_6_c_LC_17_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29426\,
            in2 => \N__27348\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.valor_max_final4_2_cry_5\,
            carryout => \b2v_inst.valor_max_final4_2_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final4_2_cry_7_c_LC_17_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29351\,
            in2 => \N__27590\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.valor_max_final4_2_cry_6\,
            carryout => \b2v_inst.valor_max_final4_2_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final4_2_cry_8_c_LC_17_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29320\,
            in2 => \N__29926\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_17_6_0_\,
            carryout => \b2v_inst.valor_max_final4_2_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final4_2_cry_9_c_LC_17_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29726\,
            in2 => \N__29291\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.valor_max_final4_2_cry_8\,
            carryout => \b2v_inst.valor_max_final4_2_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final4_2_cry_10_c_LC_17_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31489\,
            in2 => \N__29213\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.valor_max_final4_2_cry_9\,
            carryout => \b2v_inst.valor_max_final42\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final4_2_cry_10_c_RNI9G0Q_LC_17_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101101011011"
        )
    port map (
            in0 => \N__32349\,
            in1 => \N__29177\,
            in2 => \N__32542\,
            in3 => \N__27299\,
            lcout => \b2v_inst.m54_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir11_7_c_RNO_LC_17_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__30723\,
            in1 => \N__30691\,
            in2 => \N__30136\,
            in3 => \N__29443\,
            lcout => \b2v_inst.data_a_escribir11_7_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.reg_ancho_3_6_LC_17_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__31905\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31563\,
            lcout => \b2v_inst.reg_ancho_3Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34416\,
            ce => \N__32060\,
            sr => \N__38117\
        );

    \b2v_inst.reg_ancho_3_7_LC_17_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27270\,
            in2 => \_gnd_net_\,
            in3 => \N__31906\,
            lcout => \b2v_inst.reg_ancho_3Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34416\,
            ce => \N__32060\,
            sr => \N__38117\
        );

    \b2v_inst.reg_ancho_3_8_LC_17_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__31907\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27250\,
            lcout => \b2v_inst.reg_ancho_3Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34416\,
            ce => \N__32060\,
            sr => \N__38117\
        );

    \b2v_inst.reg_ancho_3_9_LC_17_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__31989\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31908\,
            lcout => \b2v_inst.reg_ancho_3Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34416\,
            ce => \N__32060\,
            sr => \N__38117\
        );

    \b2v_inst.reg_ancho_3_1_LC_17_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__31904\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31396\,
            lcout => \b2v_inst.reg_ancho_3Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34416\,
            ce => \N__32060\,
            sr => \N__38117\
        );

    \b2v_inst.reg_ancho_3_0_LC_17_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31903\,
            in2 => \_gnd_net_\,
            in3 => \N__27487\,
            lcout => \b2v_inst.reg_ancho_3Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34416\,
            ce => \N__32060\,
            sr => \N__38117\
        );

    \b2v_inst.encontrar_maximo_valor_max_final4_3_cry_0_c_LC_17_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27505\,
            in2 => \N__27448\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_17_8_0_\,
            carryout => \b2v_inst.valor_max_final4_3_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final4_3_cry_1_c_LC_17_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27745\,
            in2 => \N__31352\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.valor_max_final4_3_cry_0\,
            carryout => \b2v_inst.valor_max_final4_3_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final4_3_cry_2_c_LC_17_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27727\,
            in2 => \N__31304\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.valor_max_final4_3_cry_1\,
            carryout => \b2v_inst.valor_max_final4_3_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final4_3_cry_3_c_LC_17_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27709\,
            in2 => \N__32458\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.valor_max_final4_3_cry_2\,
            carryout => \b2v_inst.valor_max_final4_3_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final4_3_cry_4_c_LC_17_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33014\,
            in2 => \N__27692\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.valor_max_final4_3_cry_3\,
            carryout => \b2v_inst.valor_max_final4_3_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final4_3_cry_5_c_LC_17_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27393\,
            in2 => \N__27671\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.valor_max_final4_3_cry_4\,
            carryout => \b2v_inst.valor_max_final4_3_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final4_3_cry_6_c_LC_17_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27649\,
            in2 => \N__27349\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.valor_max_final4_3_cry_5\,
            carryout => \b2v_inst.valor_max_final4_3_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final4_3_cry_7_c_LC_17_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27585\,
            in2 => \N__27632\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.valor_max_final4_3_cry_6\,
            carryout => \b2v_inst.valor_max_final4_3_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final4_3_cry_8_c_LC_17_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29927\,
            in2 => \N__27611\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_17_9_0_\,
            carryout => \b2v_inst.valor_max_final4_3_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final4_3_cry_9_c_LC_17_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29737\,
            in2 => \N__28406\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.valor_max_final4_3_cry_8\,
            carryout => \b2v_inst.valor_max_final4_3_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final4_3_cry_10_c_LC_17_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31483\,
            in2 => \N__28385\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.valor_max_final4_3_cry_9\,
            carryout => \b2v_inst.valor_max_final43\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.valor_max_final43_THRU_LUT4_0_LC_17_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27542\,
            lcout => \b2v_inst.valor_max_final43_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_0_0_LC_17_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111101111111"
        )
    port map (
            in0 => \N__28615\,
            in1 => \N__32405\,
            in2 => \N__30987\,
            in3 => \N__29674\,
            lcout => \b2v_inst.data_a_escribir_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_0_1_LC_17_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111100111111"
        )
    port map (
            in0 => \N__28589\,
            in1 => \N__29701\,
            in2 => \N__30988\,
            in3 => \N__32406\,
            lcout => \b2v_inst.data_a_escribir_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_3_5_LC_17_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100110011"
        )
    port map (
            in0 => \N__27527\,
            in1 => \N__30961\,
            in2 => \_gnd_net_\,
            in3 => \N__31129\,
            lcout => \b2v_inst.un1_reg_anterior_iv_0_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final4_1_cry_0_c_inv_LC_17_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29066\,
            in2 => \N__27506\,
            in3 => \N__28610\,
            lcout => \b2v_inst.reg_anterior_i_0\,
            ltout => OPEN,
            carryin => \bfn_17_10_0_\,
            carryout => \b2v_inst.valor_max_final4_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final4_1_cry_1_c_inv_LC_17_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__28574\,
            in1 => \N__28994\,
            in2 => \N__27746\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst.reg_anterior_i_1\,
            ltout => OPEN,
            carryin => \b2v_inst.valor_max_final4_1_cry_0\,
            carryout => \b2v_inst.valor_max_final4_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final4_1_cry_2_c_inv_LC_17_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31256\,
            in2 => \N__27728\,
            in3 => \N__29837\,
            lcout => \b2v_inst.reg_anterior_i_2\,
            ltout => OPEN,
            carryin => \b2v_inst.valor_max_final4_1_cry_1\,
            carryout => \b2v_inst.valor_max_final4_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final4_1_cry_3_c_inv_LC_17_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__29158\,
            in1 => \N__31041\,
            in2 => \N__27710\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst.reg_anterior_i_3\,
            ltout => OPEN,
            carryin => \b2v_inst.valor_max_final4_1_cry_2\,
            carryout => \b2v_inst.valor_max_final4_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final4_1_cry_4_c_inv_LC_17_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29636\,
            in2 => \N__27691\,
            in3 => \N__30171\,
            lcout => \b2v_inst.reg_anterior_i_4\,
            ltout => OPEN,
            carryin => \b2v_inst.valor_max_final4_1_cry_3\,
            carryout => \b2v_inst.valor_max_final4_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final4_1_cry_5_c_inv_LC_17_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29559\,
            in2 => \N__27670\,
            in3 => \N__29101\,
            lcout => \b2v_inst.reg_anterior_i_5\,
            ltout => OPEN,
            carryin => \b2v_inst.valor_max_final4_1_cry_4\,
            carryout => \b2v_inst.valor_max_final4_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final4_1_cry_6_c_inv_LC_17_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__31525\,
            in1 => \N__29485\,
            in2 => \N__27650\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst.reg_anterior_i_6\,
            ltout => OPEN,
            carryin => \b2v_inst.valor_max_final4_1_cry_5\,
            carryout => \b2v_inst.valor_max_final4_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final4_1_cry_7_c_inv_LC_17_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29396\,
            in2 => \N__27631\,
            in3 => \N__30657\,
            lcout => \b2v_inst.reg_anterior_i_7\,
            ltout => OPEN,
            carryin => \b2v_inst.valor_max_final4_1_cry_6\,
            carryout => \b2v_inst.valor_max_final4_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final4_1_cry_8_c_inv_LC_17_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29966\,
            in2 => \N__27610\,
            in3 => \N__30761\,
            lcout => \b2v_inst.reg_anterior_i_8\,
            ltout => OPEN,
            carryin => \bfn_17_11_0_\,
            carryout => \b2v_inst.valor_max_final4_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final4_1_cry_9_c_inv_LC_17_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__31950\,
            in1 => \N__30003\,
            in2 => \N__28405\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst.reg_anterior_i_9\,
            ltout => OPEN,
            carryin => \b2v_inst.valor_max_final4_1_cry_8\,
            carryout => \b2v_inst.valor_max_final4_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final4_1_cry_10_c_inv_LC_17_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29257\,
            in2 => \N__28384\,
            in3 => \N__31719\,
            lcout => \b2v_inst.reg_anterior_i_10\,
            ltout => OPEN,
            carryin => \b2v_inst.valor_max_final4_1_cry_9\,
            carryout => \b2v_inst.valor_max_final41\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final4_3_cry_10_c_RNIUCPE1_LC_17_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011010011110100"
        )
    port map (
            in0 => \N__28364\,
            in1 => \N__32398\,
            in2 => \N__28355\,
            in3 => \N__28343\,
            lcout => \b2v_inst.N_711\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.reg_anterior_1_LC_17_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31858\,
            in2 => \_gnd_net_\,
            in3 => \N__31400\,
            lcout => \b2v_inst.reg_anteriorZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34380\,
            ce => \N__31672\,
            sr => \N__38107\
        );

    \b2v_inst.state_RNO_4_31_LC_17_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__28340\,
            in1 => \N__28206\,
            in2 => \N__27920\,
            in3 => \N__28253\,
            lcout => \b2v_inst.N_694\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNO_5_31_LC_17_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__28207\,
            in1 => \N__28076\,
            in2 => \N__28067\,
            in3 => \N__27918\,
            lcout => OPEN,
            ltout => \b2v_inst.N_695_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNO_0_31_LC_17_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__27962\,
            in1 => \N__28025\,
            in2 => \N__28019\,
            in3 => \N__28004\,
            lcout => \b2v_inst.state_ns_a3_i_0_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_32_rep1_RNIUROT1_LC_17_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111110000"
        )
    port map (
            in0 => \N__28003\,
            in1 => \N__27961\,
            in2 => \N__30983\,
            in3 => \N__27917\,
            lcout => OPEN,
            ltout => \b2v_inst.un1_reset_inv_0_0_tz_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_32_rep1_RNIP5K4F_LC_17_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010101000"
        )
    port map (
            in0 => \N__27833\,
            in1 => \N__28546\,
            in2 => \N__28529\,
            in3 => \N__28525\,
            lcout => \b2v_inst.un1_reset_inv_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_1_7_LC_17_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101001111111"
        )
    port map (
            in0 => \N__31176\,
            in1 => \N__30956\,
            in2 => \N__28490\,
            in3 => \N__28469\,
            lcout => \b2v_inst.un1_reg_anterior_0_i_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst9.un1_cycle_counter_2_cry_0_c_LC_17_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30416\,
            in2 => \N__30308\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_17_13_0_\,
            carryout => \b2v_inst9.un1_cycle_counter_2_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst9.un1_cycle_counter_2_cry_0_THRU_LUT4_0_LC_17_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__28427\,
            in3 => \N__28463\,
            lcout => \b2v_inst9.un1_cycle_counter_2_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst9.un1_cycle_counter_2_cry_0\,
            carryout => \b2v_inst9.un1_cycle_counter_2_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst9.un1_cycle_counter_2_cry_1_THRU_LUT4_0_LC_17_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30493\,
            in2 => \_gnd_net_\,
            in3 => \N__28460\,
            lcout => \b2v_inst9.un1_cycle_counter_2_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst9.un1_cycle_counter_2_cry_1\,
            carryout => \b2v_inst9.un1_cycle_counter_2_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst9.cycle_counter_3_LC_17_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__28453\,
            in1 => \N__38151\,
            in2 => \_gnd_net_\,
            in3 => \N__28457\,
            lcout => \b2v_inst9.cycle_counterZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34397\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst9.cycle_counter_RNIQAGD_0_3_LC_17_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__30304\,
            in1 => \N__28452\,
            in2 => \N__28426\,
            in3 => \N__30492\,
            lcout => \b2v_inst9.N_175_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst9.cycle_counter_RNIQAGD_3_LC_17_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__30491\,
            in1 => \N__28418\,
            in2 => \N__28454\,
            in3 => \N__30303\,
            lcout => \b2v_inst9.cycle_counter_RNIQAGDZ0Z_3\,
            ltout => \b2v_inst9.cycle_counter_RNIQAGDZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst9.cycle_counter_1_LC_17_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000000100000"
        )
    port map (
            in0 => \N__28425\,
            in1 => \N__38150\,
            in2 => \N__28436\,
            in3 => \N__28433\,
            lcout => \b2v_inst9.cycle_counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34397\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un12_pix_count_intlto7_N_3L3_LC_17_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101010101"
        )
    port map (
            in0 => \N__28852\,
            in1 => \N__28839\,
            in2 => \_gnd_net_\,
            in3 => \N__28795\,
            lcout => \b2v_inst.un12_pix_count_intlto7_N_3LZ0Z3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst4.reg_data_5_LC_17_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28817\,
            lcout => \SYNTHESIZED_WIRE_5_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34417\,
            ce => \N__28784\,
            sr => \N__38130\
        );

    \b2v_inst9.bit_counter_0_LC_17_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28654\,
            in1 => \N__28709\,
            in2 => \N__28727\,
            in3 => \N__28726\,
            lcout => \b2v_inst9.bit_counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_17_16_0_\,
            carryout => \b2v_inst9.un1_bit_counter_3_cry_0\,
            clk => \N__34426\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst9.bit_counter_1_LC_17_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28652\,
            in1 => \N__28694\,
            in2 => \_gnd_net_\,
            in3 => \N__28679\,
            lcout => \b2v_inst9.bit_counterZ1Z_1\,
            ltout => OPEN,
            carryin => \b2v_inst9.un1_bit_counter_3_cry_0\,
            carryout => \b2v_inst9.un1_bit_counter_3_cry_1\,
            clk => \N__34426\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst9.bit_counter_2_LC_17_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28655\,
            in1 => \N__28675\,
            in2 => \_gnd_net_\,
            in3 => \N__28658\,
            lcout => \b2v_inst9.bit_counterZ0Z_2\,
            ltout => OPEN,
            carryin => \b2v_inst9.un1_bit_counter_3_cry_1\,
            carryout => \b2v_inst9.un1_bit_counter_3_cry_2\,
            clk => \N__34426\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst9.bit_counter_3_LC_17_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28653\,
            in1 => \N__28634\,
            in2 => \_gnd_net_\,
            in3 => \N__28637\,
            lcout => \b2v_inst9.bit_counterZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34426\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.reg_anterior_5_LC_18_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31919\,
            in2 => \_gnd_net_\,
            in3 => \N__32117\,
            lcout => \b2v_inst.reg_anteriorZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34427\,
            ce => \N__31687\,
            sr => \N__38136\
        );

    \b2v_inst.encontrar_maximo_un2_valor_max2_cry_0_c_LC_18_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28619\,
            in2 => \N__29024\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_18_6_0_\,
            carryout => \b2v_inst.un2_valor_max2_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_un2_valor_max2_cry_1_c_LC_18_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28584\,
            in2 => \N__28952\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.un2_valor_max2_cry_0\,
            carryout => \b2v_inst.un2_valor_max2_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_un2_valor_max2_cry_2_c_LC_18_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29839\,
            in2 => \N__28915\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.un2_valor_max2_cry_1\,
            carryout => \b2v_inst.un2_valor_max2_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_un2_valor_max2_cry_3_c_LC_18_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29153\,
            in2 => \N__28883\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.un2_valor_max2_cry_2\,
            carryout => \b2v_inst.un2_valor_max2_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_un2_valor_max2_cry_4_c_LC_18_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30158\,
            in2 => \N__29590\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.un2_valor_max2_cry_3\,
            carryout => \b2v_inst.un2_valor_max2_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_un2_valor_max2_cry_5_c_LC_18_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29090\,
            in2 => \N__29513\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.un2_valor_max2_cry_4\,
            carryout => \b2v_inst.un2_valor_max2_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_un2_valor_max2_cry_6_c_LC_18_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31514\,
            in2 => \N__29425\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.un2_valor_max2_cry_5\,
            carryout => \b2v_inst.un2_valor_max2_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_un2_valor_max2_cry_7_c_LC_18_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30669\,
            in2 => \N__29350\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.un2_valor_max2_cry_6\,
            carryout => \b2v_inst.un2_valor_max2_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_un2_valor_max2_cry_8_c_LC_18_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30770\,
            in2 => \N__29321\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_18_7_0_\,
            carryout => \b2v_inst.un2_valor_max2_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_un2_valor_max2_cry_9_c_LC_18_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31955\,
            in2 => \N__29290\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.un2_valor_max2_cry_8\,
            carryout => \b2v_inst.un2_valor_max2_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_un2_valor_max2_cry_10_c_LC_18_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31726\,
            in2 => \N__29212\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.un2_valor_max2_cry_9\,
            carryout => \b2v_inst.un2_valor_max2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un2_valor_max2_THRU_LUT4_0_LC_18_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29165\,
            lcout => \b2v_inst.un2_valor_max2_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_0_3_LC_18_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111101011111"
        )
    port map (
            in0 => \N__32231\,
            in1 => \N__29162\,
            in2 => \N__30992\,
            in3 => \N__32392\,
            lcout => \b2v_inst.data_a_escribir_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_0_6_LC_18_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32393\,
            in1 => \N__31518\,
            in2 => \_gnd_net_\,
            in3 => \N__29444\,
            lcout => \b2v_inst.valor_max2_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_0_5_LC_18_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32391\,
            in1 => \N__29097\,
            in2 => \_gnd_net_\,
            in3 => \N__32083\,
            lcout => \b2v_inst.N_267\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final4_0_cry_0_c_inv_LC_18_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__29664\,
            in1 => \N__29065\,
            in2 => \N__29022\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst.reg_ancho_3_i_0\,
            ltout => OPEN,
            carryin => \bfn_18_8_0_\,
            carryout => \b2v_inst.valor_max_final4_0_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final4_0_cry_1_c_inv_LC_18_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28990\,
            in2 => \N__28944\,
            in3 => \N__29691\,
            lcout => \b2v_inst.reg_ancho_3_i_1\,
            ltout => OPEN,
            carryin => \b2v_inst.valor_max_final4_0_cry_0\,
            carryout => \b2v_inst.valor_max_final4_0_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final4_0_cry_2_c_inv_LC_18_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31245\,
            in2 => \N__28911\,
            in3 => \N__32153\,
            lcout => \b2v_inst.reg_ancho_3_i_2\,
            ltout => OPEN,
            carryin => \b2v_inst.valor_max_final4_0_cry_1\,
            carryout => \b2v_inst.valor_max_final4_0_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final4_0_cry_3_c_inv_LC_18_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__32230\,
            in1 => \N__31037\,
            in2 => \N__28881\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst.reg_ancho_3_i_3\,
            ltout => OPEN,
            carryin => \b2v_inst.valor_max_final4_0_cry_2\,
            carryout => \b2v_inst.valor_max_final4_0_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final4_0_cry_4_c_inv_LC_18_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29635\,
            in2 => \N__29589\,
            in3 => \N__31426\,
            lcout => \b2v_inst.reg_ancho_3_i_4\,
            ltout => OPEN,
            carryin => \b2v_inst.valor_max_final4_0_cry_3\,
            carryout => \b2v_inst.valor_max_final4_0_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final4_0_cry_5_c_inv_LC_18_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29505\,
            in2 => \N__29561\,
            in3 => \N__32082\,
            lcout => \b2v_inst.reg_ancho_3_i_5\,
            ltout => OPEN,
            carryin => \b2v_inst.valor_max_final4_0_cry_4\,
            carryout => \b2v_inst.valor_max_final4_0_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final4_0_cry_6_c_inv_LC_18_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29484\,
            in2 => \N__29424\,
            in3 => \N__29442\,
            lcout => \b2v_inst.reg_ancho_3_i_6\,
            ltout => OPEN,
            carryin => \b2v_inst.valor_max_final4_0_cry_5\,
            carryout => \b2v_inst.valor_max_final4_0_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final4_0_cry_7_c_inv_LC_18_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29391\,
            in2 => \N__29349\,
            in3 => \N__30690\,
            lcout => \b2v_inst.reg_ancho_3_i_7\,
            ltout => OPEN,
            carryin => \b2v_inst.valor_max_final4_0_cry_6\,
            carryout => \b2v_inst.valor_max_final4_0_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final4_0_cry_8_c_inv_LC_18_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__30724\,
            in1 => \N__29964\,
            in2 => \N__29319\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst.reg_ancho_3_i_8\,
            ltout => OPEN,
            carryin => \bfn_18_9_0_\,
            carryout => \b2v_inst.valor_max_final4_0_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final4_0_cry_9_c_inv_LC_18_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30004\,
            in2 => \N__29286\,
            in3 => \N__30132\,
            lcout => \b2v_inst.reg_ancho_3_i_9\,
            ltout => OPEN,
            carryin => \b2v_inst.valor_max_final4_0_cry_8\,
            carryout => \b2v_inst.valor_max_final4_0_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final4_0_cry_10_c_inv_LC_18_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29256\,
            in2 => \N__29208\,
            in3 => \N__32301\,
            lcout => \b2v_inst.reg_ancho_3_i_10\,
            ltout => OPEN,
            carryin => \b2v_inst.valor_max_final4_0_cry_9\,
            carryout => \b2v_inst.valor_max_final40\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.valor_max_final40_THRU_LUT4_0_LC_18_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29180\,
            lcout => \b2v_inst.valor_max_final40_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_0_9_LC_18_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__32546\,
            in1 => \_gnd_net_\,
            in2 => \N__29741\,
            in3 => \N__30005\,
            lcout => \b2v_inst.N_543\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_0_8_LC_18_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__29965\,
            in1 => \N__29925\,
            in2 => \_gnd_net_\,
            in3 => \N__32545\,
            lcout => \b2v_inst.N_542\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_1_3_LC_18_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110001111111"
        )
    port map (
            in0 => \N__30971\,
            in1 => \N__31180\,
            in2 => \N__29873\,
            in3 => \N__32465\,
            lcout => \b2v_inst.un1_reg_anterior_0_i_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_0_2_LC_18_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111100111111"
        )
    port map (
            in0 => \N__29838\,
            in1 => \N__32152\,
            in2 => \N__30989\,
            in3 => \N__32397\,
            lcout => \b2v_inst.data_a_escribir_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir11_6_c_RNO_LC_18_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__31438\,
            in1 => \N__32229\,
            in2 => \N__32084\,
            in3 => \N__32151\,
            lcout => \b2v_inst.data_a_escribir11_6_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_1_5_LC_18_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110001"
        )
    port map (
            in0 => \N__31177\,
            in1 => \N__29789\,
            in2 => \N__29774\,
            in3 => \N__30627\,
            lcout => OPEN,
            ltout => \b2v_inst.un1_reg_anterior_iv_0_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_5_LC_18_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100001101"
        )
    port map (
            in0 => \N__30629\,
            in1 => \N__29765\,
            in2 => \N__29753\,
            in3 => \N__31179\,
            lcout => b2v_inst_data_a_escribir_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34381\,
            ce => \N__30555\,
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_2_LC_18_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001111001110"
        )
    port map (
            in0 => \N__30628\,
            in1 => \N__31178\,
            in2 => \N__29750\,
            in3 => \N__31049\,
            lcout => b2v_inst_data_a_escribir_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34381\,
            ce => \N__30555\,
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir11_5_c_RNO_LC_18_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__29736\,
            in1 => \N__29702\,
            in2 => \N__31488\,
            in3 => \N__29675\,
            lcout => \b2v_inst.data_a_escribir11_5_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_2_9_LC_18_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__31954\,
            in1 => \N__30137\,
            in2 => \_gnd_net_\,
            in3 => \N__32407\,
            lcout => \b2v_inst.N_545\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_3_9_LC_18_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100110011"
        )
    port map (
            in0 => \N__30110\,
            in1 => \N__30957\,
            in2 => \_gnd_net_\,
            in3 => \N__31168\,
            lcout => OPEN,
            ltout => \b2v_inst.un1_reg_anterior_iv_0_0_0_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_1_9_LC_18_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111110000"
        )
    port map (
            in0 => \N__31169\,
            in1 => \N__30095\,
            in2 => \N__30089\,
            in3 => \N__30609\,
            lcout => OPEN,
            ltout => \b2v_inst.un1_reg_anterior_iv_0_0_1_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_9_LC_18_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100001110"
        )
    port map (
            in0 => \N__30611\,
            in1 => \N__30086\,
            in2 => \N__30077\,
            in3 => \N__31171\,
            lcout => b2v_inst_data_a_escribir_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34378\,
            ce => \N__30557\,
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_6_LC_18_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111101"
        )
    port map (
            in0 => \N__30610\,
            in1 => \N__31170\,
            in2 => \N__30074\,
            in3 => \N__30059\,
            lcout => b2v_inst_data_a_escribir_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34378\,
            ce => \N__30557\,
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir11_10_c_RNO_LC_18_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__31946\,
            in1 => \N__30768\,
            in2 => \N__31730\,
            in3 => \N__30670\,
            lcout => \b2v_inst.data_a_escribir11_10_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_3_8_LC_18_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100110011"
        )
    port map (
            in0 => \N__30038\,
            in1 => \N__30990\,
            in2 => \_gnd_net_\,
            in3 => \N__31172\,
            lcout => OPEN,
            ltout => \b2v_inst.un1_reg_anterior_iv_0_0_0_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_1_8_LC_18_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111110000"
        )
    port map (
            in0 => \N__31173\,
            in1 => \N__30704\,
            in2 => \N__30020\,
            in3 => \N__30622\,
            lcout => OPEN,
            ltout => \b2v_inst.un1_reg_anterior_iv_0_0_1_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_8_LC_18_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100001110"
        )
    port map (
            in0 => \N__30623\,
            in1 => \N__30017\,
            in2 => \N__30008\,
            in3 => \N__31175\,
            lcout => b2v_inst_data_a_escribir_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34382\,
            ce => \N__30554\,
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_2_8_LC_18_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30769\,
            in1 => \N__30728\,
            in2 => \_gnd_net_\,
            in3 => \N__32395\,
            lcout => \b2v_inst.N_544\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_0_7_LC_18_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101111111111"
        )
    port map (
            in0 => \N__32396\,
            in1 => \N__30698\,
            in2 => \N__30674\,
            in3 => \N__30991\,
            lcout => OPEN,
            ltout => \b2v_inst.data_a_escribir_RNO_0Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_7_LC_18_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010011101100110"
        )
    port map (
            in0 => \N__31174\,
            in1 => \N__30638\,
            in2 => \N__30632\,
            in3 => \N__30624\,
            lcout => b2v_inst_data_a_escribir_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34382\,
            ce => \N__30554\,
            sr => \_gnd_net_\
        );

    \b2v_inst9.cycle_counter_2_LC_18_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001000100000"
        )
    port map (
            in0 => \N__30467\,
            in1 => \N__38155\,
            in2 => \N__30497\,
            in3 => \N__30503\,
            lcout => \b2v_inst9.cycle_counterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34392\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst9.cycle_counter_0_LC_18_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010000001000"
        )
    port map (
            in0 => \N__30302\,
            in1 => \N__30466\,
            in2 => \N__38156\,
            in3 => \N__30433\,
            lcout => \b2v_inst9.cycle_counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34392\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.pix_data_reg_3_LC_18_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30281\,
            lcout => \b2v_inst.pix_data_regZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34398\,
            ce => \N__30248\,
            sr => \N__38131\
        );

    \b2v_inst.cantidad_temp_2_LC_18_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__34765\,
            in1 => \N__32656\,
            in2 => \N__30191\,
            in3 => \N__34642\,
            lcout => b2v_inst_cantidad_temp_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34409\,
            ce => 'H',
            sr => \N__38137\
        );

    \b2v_inst.reg_anterior_4_LC_19_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31917\,
            in2 => \_gnd_net_\,
            in3 => \N__33050\,
            lcout => \b2v_inst.reg_anteriorZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34410\,
            ce => \N__31673\,
            sr => \N__38138\
        );

    \b2v_inst.reg_anterior_6_LC_19_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__31918\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31562\,
            lcout => \b2v_inst.reg_anteriorZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34410\,
            ce => \N__31673\,
            sr => \N__38138\
        );

    \b2v_inst.reg_ancho_2_10_LC_19_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31780\,
            lcout => \b2v_inst.reg_ancho_2Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34399\,
            ce => \N__32959\,
            sr => \N__38132\
        );

    \b2v_inst.reg_ancho_3_4_LC_19_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31902\,
            in2 => \_gnd_net_\,
            in3 => \N__33061\,
            lcout => \b2v_inst.reg_ancho_3Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34393\,
            ce => \N__32059\,
            sr => \N__38124\
        );

    \b2v_inst.data_a_escribir11_3_c_RNO_LC_19_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__32434\,
            in1 => \N__31282\,
            in2 => \N__33010\,
            in3 => \N__31330\,
            lcout => \b2v_inst.data_a_escribir11_3_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.reg_ancho_2_1_LC_19_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31395\,
            lcout => \b2v_inst.reg_ancho_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34383\,
            ce => \N__32965\,
            sr => \N__38118\
        );

    \b2v_inst.reg_ancho_2_2_LC_19_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32209\,
            lcout => \b2v_inst.reg_ancho_2Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34383\,
            ce => \N__32965\,
            sr => \N__38118\
        );

    \b2v_inst.data_a_escribir_RNO_2_2_LC_19_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111100111111"
        )
    port map (
            in0 => \N__31283\,
            in1 => \N__31255\,
            in2 => \N__30979\,
            in3 => \N__32544\,
            lcout => OPEN,
            ltout => \b2v_inst.data_a_escribir_RNO_2Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_1_2_LC_19_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100001111"
        )
    port map (
            in0 => \N__31202\,
            in1 => \N__30941\,
            in2 => \N__31184\,
            in3 => \N__31181\,
            lcout => \b2v_inst.un1_reg_anterior_0_i_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_2_3_LC_19_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111100111111"
        )
    port map (
            in0 => \N__32438\,
            in1 => \N__31043\,
            in2 => \N__30978\,
            in3 => \N__32543\,
            lcout => \b2v_inst.data_a_escribir_RNO_2Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.reg_ancho_2_3_LC_19_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32283\,
            lcout => \b2v_inst.reg_ancho_2Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34383\,
            ce => \N__32965\,
            sr => \N__38118\
        );

    \b2v_inst.data_a_escribir_RNO_0_10_LC_19_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__31718\,
            in1 => \N__32305\,
            in2 => \_gnd_net_\,
            in3 => \N__32394\,
            lcout => \b2v_inst.N_264\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.reg_ancho_3_10_LC_19_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31898\,
            in2 => \_gnd_net_\,
            in3 => \N__31776\,
            lcout => \b2v_inst.reg_ancho_3Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34379\,
            ce => \N__32052\,
            sr => \N__38108\
        );

    \b2v_inst.reg_ancho_3_3_LC_19_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__31900\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32284\,
            lcout => \b2v_inst.reg_ancho_3Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34379\,
            ce => \N__32052\,
            sr => \N__38108\
        );

    \b2v_inst.reg_ancho_3_2_LC_19_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31899\,
            in2 => \_gnd_net_\,
            in3 => \N__32205\,
            lcout => \b2v_inst.reg_ancho_3Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34379\,
            ce => \N__32052\,
            sr => \N__38108\
        );

    \b2v_inst.reg_ancho_3_5_LC_19_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__31901\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32131\,
            lcout => \b2v_inst.reg_ancho_3Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34379\,
            ce => \N__32052\,
            sr => \N__38108\
        );

    \b2v_inst.reg_anterior_9_LC_19_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__31897\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31985\,
            lcout => \b2v_inst.reg_anteriorZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34373\,
            ce => \N__31688\,
            sr => \N__38119\
        );

    \b2v_inst.reg_anterior_10_LC_19_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31896\,
            in2 => \_gnd_net_\,
            in3 => \N__31772\,
            lcout => \b2v_inst.reg_anteriorZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34373\,
            ce => \N__31688\,
            sr => \N__38119\
        );

    \b2v_inst.cantidad_temp_0_LC_19_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__34908\,
            in1 => \N__34627\,
            in2 => \N__32705\,
            in3 => \N__34762\,
            lcout => b2v_inst_cantidad_temp_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34384\,
            ce => 'H',
            sr => \N__38133\
        );

    \b2v_inst.cantidad_temp_1_LC_19_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__34628\,
            in1 => \N__34870\,
            in2 => \N__32690\,
            in3 => \N__34764\,
            lcout => b2v_inst_cantidad_temp_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34384\,
            ce => 'H',
            sr => \N__38133\
        );

    \b2v_inst.cantidad_temp_4_LC_19_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__32623\,
            in1 => \N__34629\,
            in2 => \N__32678\,
            in3 => \N__34763\,
            lcout => b2v_inst_cantidad_temp_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34384\,
            ce => 'H',
            sr => \N__38133\
        );

    \b2v_inst.un16_data_ram_cantidad_o_cry_1_c_LC_19_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34865\,
            in2 => \N__34909\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_19_14_0_\,
            carryout => \b2v_inst.un16_data_ram_cantidad_o_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un16_data_ram_cantidad_o_cry_1_c_RNI77CO_LC_19_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32652\,
            in2 => \_gnd_net_\,
            in3 => \N__32636\,
            lcout => \b2v_inst.un16_data_ram_cantidad_o_cry_1_c_RNI77COZ0\,
            ltout => OPEN,
            carryin => \b2v_inst.un16_data_ram_cantidad_o_cry_1\,
            carryout => \b2v_inst.un16_data_ram_cantidad_o_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un16_data_ram_cantidad_o_cry_2_c_RNI9ADO_LC_19_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34545\,
            in2 => \_gnd_net_\,
            in3 => \N__32633\,
            lcout => \b2v_inst.un16_data_ram_cantidad_o_cry_2_c_RNI9ADOZ0\,
            ltout => OPEN,
            carryin => \b2v_inst.un16_data_ram_cantidad_o_cry_2\,
            carryout => \b2v_inst.un16_data_ram_cantidad_o_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un16_data_ram_cantidad_o_cry_3_c_RNIBDEO_LC_19_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32619\,
            in2 => \_gnd_net_\,
            in3 => \N__32603\,
            lcout => \b2v_inst.un16_data_ram_cantidad_o_cry_3_c_RNIBDEOZ0\,
            ltout => OPEN,
            carryin => \b2v_inst.un16_data_ram_cantidad_o_cry_3\,
            carryout => \b2v_inst.un16_data_ram_cantidad_o_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un16_data_ram_cantidad_o_cry_4_c_RNIDGFO_LC_19_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32599\,
            in2 => \_gnd_net_\,
            in3 => \N__32567\,
            lcout => \b2v_inst.un16_data_ram_cantidad_o_cry_4_c_RNIDGFOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNIH17G1_2_LC_19_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__37792\,
            in1 => \N__32564\,
            in2 => \N__33140\,
            in3 => \N__37547\,
            lcout => \N_553_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNIN99G1_4_LC_19_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__37808\,
            in1 => \N__33347\,
            in2 => \N__33329\,
            in3 => \N__37530\,
            lcout => \N_549_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNIK58G1_3_LC_19_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__37807\,
            in1 => \N__33263\,
            in2 => \N__33257\,
            in3 => \N__37531\,
            lcout => \N_551_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNIHBT91_10_LC_19_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35196\,
            in2 => \_gnd_net_\,
            in3 => \N__33188\,
            lcout => \b2v_inst.N_645\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNI8OQN_0_LC_20_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010101010"
        )
    port map (
            in0 => \N__34976\,
            in1 => \N__37841\,
            in2 => \_gnd_net_\,
            in3 => \N__37561\,
            lcout => \N_121_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNIAQQN_2_LC_20_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010101010"
        )
    port map (
            in0 => \N__33124\,
            in1 => \N__37836\,
            in2 => \_gnd_net_\,
            in3 => \N__37562\,
            lcout => \N_118_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.reg_ancho_2_4_LC_20_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33054\,
            lcout => \b2v_inst.reg_ancho_2Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34385\,
            ce => \N__32966\,
            sr => \N__38134\
        );

    \b2v_inst.data_a_escribir_RNIH1RN_9_LC_20_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010101010"
        )
    port map (
            in0 => \N__32859\,
            in1 => \N__37823\,
            in2 => \_gnd_net_\,
            in3 => \N__37497\,
            lcout => \N_111_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_RNI1E333_6_LC_20_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__32819\,
            in1 => \N__38377\,
            in2 => \N__32801\,
            in3 => \N__35240\,
            lcout => \N_298\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_RNIS8333_5_LC_20_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__35243\,
            in1 => \N__34046\,
            in2 => \N__34031\,
            in3 => \N__35726\,
            lcout => \indice_RNIS8333_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_RNIBO333_8_LC_20_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__35241\,
            in1 => \N__33929\,
            in2 => \N__33911\,
            in3 => \N__39081\,
            lcout => \indice_RNIBO333_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_RNIGT333_9_LC_20_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__33812\,
            in1 => \N__35953\,
            in2 => \N__33797\,
            in3 => \N__35242\,
            lcout => \indice_RNIGT333_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNIDTQN_5_LC_20_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101000101010"
        )
    port map (
            in0 => \N__37598\,
            in1 => \N__37819\,
            in2 => \N__37560\,
            in3 => \_gnd_net_\,
            lcout => \N_115_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNIPNGN_10_LC_20_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37550\,
            in2 => \N__37835\,
            in3 => \N__33669\,
            lcout => \N_110_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_RNI3F233_0_LC_20_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__33620\,
            in1 => \N__35238\,
            in2 => \N__33605\,
            in3 => \N__39318\,
            lcout => \indice_RNI3F233_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_RNIO3V73_10_LC_20_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__35239\,
            in1 => \N__33512\,
            in2 => \N__33494\,
            in3 => \N__36751\,
            lcout => \N_37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNIG0RN_8_LC_20_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111100000000"
        )
    port map (
            in0 => \N__37544\,
            in1 => \_gnd_net_\,
            in2 => \N__37840\,
            in3 => \N__33381\,
            lcout => \N_112_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNIFVQN_7_LC_20_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010101010"
        )
    port map (
            in0 => \N__35484\,
            in1 => \N__37831\,
            in2 => \_gnd_net_\,
            in3 => \N__37543\,
            lcout => \N_113_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_RNI8K233_1_LC_20_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__35450\,
            in1 => \N__35209\,
            in2 => \N__35432\,
            in3 => \N__38660\,
            lcout => \indice_RNI8K233_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNIEUQN_6_LC_20_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010101010"
        )
    port map (
            in0 => \N__35315\,
            in1 => \N__37809\,
            in2 => \_gnd_net_\,
            in3 => \N__37545\,
            lcout => \N_114_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_RNIDP233_2_LC_20_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__35258\,
            in1 => \N__35208\,
            in2 => \N__35075\,
            in3 => \N__36122\,
            lcout => \indice_RNIDP233_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNIIIS11_0_LC_20_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100001011101"
        )
    port map (
            in0 => \N__37546\,
            in1 => \N__34975\,
            in2 => \N__37830\,
            in3 => \N__34907\,
            lcout => \N_557_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.cantidad_temp_RNILL3K_1_LC_20_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34903\,
            in2 => \_gnd_net_\,
            in3 => \N__34866\,
            lcout => OPEN,
            ltout => \b2v_inst.cantidad_temp_RNILL3KZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNIUEUB1_1_LC_20_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__34840\,
            in1 => \N__37549\,
            in2 => \N__34775\,
            in3 => \N__37793\,
            lcout => \N_555_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.cantidad_temp_3_LC_20_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__34549\,
            in1 => \N__34766\,
            in2 => \N__34652\,
            in3 => \N__34643\,
            lcout => b2v_inst_cantidad_temp_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34386\,
            ce => 'H',
            sr => \N__38139\
        );

    \b2v_inst.data_a_escribir_RNIQDAG1_5_LC_20_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__37813\,
            in1 => \N__37637\,
            in2 => \N__37627\,
            in3 => \N__37548\,
            lcout => \N_547_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_20_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_energia_RNIFL4P2_10_LC_20_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001010000"
        )
    port map (
            in0 => \N__38458\,
            in1 => \N__36788\,
            in2 => \N__36752\,
            in3 => \N__38242\,
            lcout => \N_445_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_energia_RNIJFLU2_3_LC_20_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__36581\,
            in1 => \N__38460\,
            in2 => \N__36467\,
            in3 => \N__38246\,
            lcout => \N_357_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_energia_RNILHLU2_4_LC_20_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001000100"
        )
    port map (
            in0 => \N__38461\,
            in1 => \N__36376\,
            in2 => \N__36257\,
            in3 => \N__38244\,
            lcout => \N_356_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_energia_RNIHDLU2_2_LC_20_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101000000"
        )
    port map (
            in0 => \N__38459\,
            in1 => \N__38243\,
            in2 => \N__36164\,
            in3 => \N__36121\,
            lcout => \N_358_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_energia_RNIVRLU2_9_LC_20_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001000100"
        )
    port map (
            in0 => \N__38463\,
            in1 => \N__35933\,
            in2 => \N__35831\,
            in3 => \N__38245\,
            lcout => \N_444_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_energia_RNINJLU2_5_LC_20_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__35722\,
            in1 => \N__38462\,
            in2 => \N__35594\,
            in3 => \N__38247\,
            lcout => \N_355_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_energia_RNID9LU2_0_LC_20_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101000000"
        )
    port map (
            in0 => \N__38464\,
            in1 => \N__38260\,
            in2 => \N__39383\,
            in3 => \N__39323\,
            lcout => \N_360_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_energia_RNITPLU2_8_LC_20_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001010000"
        )
    port map (
            in0 => \N__38468\,
            in1 => \N__39146\,
            in2 => \N__39100\,
            in3 => \N__38264\,
            lcout => \N_443_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_energia_RNIRNLU2_7_LC_20_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__38263\,
            in1 => \N__38467\,
            in2 => \N__38927\,
            in3 => \N__38866\,
            lcout => \N_353_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_energia_RNIFBLU2_1_LC_20_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101000000"
        )
    port map (
            in0 => \N__38465\,
            in1 => \N__38261\,
            in2 => \N__38714\,
            in3 => \N__38666\,
            lcout => \N_359_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_energia_RNIPLLU2_6_LC_20_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001010000"
        )
    port map (
            in0 => \N__38466\,
            in1 => \N__38429\,
            in2 => \N__38381\,
            in3 => \N__38262\,
            lcout => \N_354_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
