-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Oct 3 2024 21:30:25

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "anda_plis" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of anda_plis
entity anda_plis is
port (
    uart_tx_o : out std_logic;
    uart_rx_i : in std_logic;
    reset : in std_logic;
    clk : in std_logic);
end anda_plis;

-- Architecture of anda_plis
-- View name is \INTERFACE\
architecture \INTERFACE\ of anda_plis is

signal \N__24159\ : std_logic;
signal \N__24158\ : std_logic;
signal \N__24157\ : std_logic;
signal \N__24150\ : std_logic;
signal \N__24149\ : std_logic;
signal \N__24148\ : std_logic;
signal \N__24141\ : std_logic;
signal \N__24140\ : std_logic;
signal \N__24139\ : std_logic;
signal \N__24132\ : std_logic;
signal \N__24131\ : std_logic;
signal \N__24130\ : std_logic;
signal \N__24113\ : std_logic;
signal \N__24110\ : std_logic;
signal \N__24107\ : std_logic;
signal \N__24104\ : std_logic;
signal \N__24101\ : std_logic;
signal \N__24098\ : std_logic;
signal \N__24095\ : std_logic;
signal \N__24094\ : std_logic;
signal \N__24093\ : std_logic;
signal \N__24092\ : std_logic;
signal \N__24089\ : std_logic;
signal \N__24086\ : std_logic;
signal \N__24083\ : std_logic;
signal \N__24082\ : std_logic;
signal \N__24081\ : std_logic;
signal \N__24078\ : std_logic;
signal \N__24073\ : std_logic;
signal \N__24070\ : std_logic;
signal \N__24067\ : std_logic;
signal \N__24064\ : std_logic;
signal \N__24063\ : std_logic;
signal \N__24060\ : std_logic;
signal \N__24057\ : std_logic;
signal \N__24054\ : std_logic;
signal \N__24051\ : std_logic;
signal \N__24048\ : std_logic;
signal \N__24045\ : std_logic;
signal \N__24042\ : std_logic;
signal \N__24037\ : std_logic;
signal \N__24032\ : std_logic;
signal \N__24029\ : std_logic;
signal \N__24020\ : std_logic;
signal \N__24019\ : std_logic;
signal \N__24018\ : std_logic;
signal \N__24017\ : std_logic;
signal \N__24016\ : std_logic;
signal \N__24015\ : std_logic;
signal \N__24014\ : std_logic;
signal \N__24011\ : std_logic;
signal \N__24006\ : std_logic;
signal \N__24005\ : std_logic;
signal \N__24004\ : std_logic;
signal \N__24003\ : std_logic;
signal \N__23998\ : std_logic;
signal \N__23993\ : std_logic;
signal \N__23992\ : std_logic;
signal \N__23991\ : std_logic;
signal \N__23990\ : std_logic;
signal \N__23989\ : std_logic;
signal \N__23988\ : std_logic;
signal \N__23987\ : std_logic;
signal \N__23986\ : std_logic;
signal \N__23985\ : std_logic;
signal \N__23984\ : std_logic;
signal \N__23981\ : std_logic;
signal \N__23978\ : std_logic;
signal \N__23973\ : std_logic;
signal \N__23970\ : std_logic;
signal \N__23965\ : std_logic;
signal \N__23960\ : std_logic;
signal \N__23957\ : std_logic;
signal \N__23950\ : std_logic;
signal \N__23947\ : std_logic;
signal \N__23942\ : std_logic;
signal \N__23921\ : std_logic;
signal \N__23920\ : std_logic;
signal \N__23919\ : std_logic;
signal \N__23918\ : std_logic;
signal \N__23917\ : std_logic;
signal \N__23916\ : std_logic;
signal \N__23915\ : std_logic;
signal \N__23914\ : std_logic;
signal \N__23913\ : std_logic;
signal \N__23912\ : std_logic;
signal \N__23911\ : std_logic;
signal \N__23910\ : std_logic;
signal \N__23905\ : std_logic;
signal \N__23904\ : std_logic;
signal \N__23903\ : std_logic;
signal \N__23902\ : std_logic;
signal \N__23901\ : std_logic;
signal \N__23900\ : std_logic;
signal \N__23897\ : std_logic;
signal \N__23894\ : std_logic;
signal \N__23891\ : std_logic;
signal \N__23886\ : std_logic;
signal \N__23883\ : std_logic;
signal \N__23878\ : std_logic;
signal \N__23873\ : std_logic;
signal \N__23870\ : std_logic;
signal \N__23863\ : std_logic;
signal \N__23858\ : std_logic;
signal \N__23837\ : std_logic;
signal \N__23836\ : std_logic;
signal \N__23835\ : std_logic;
signal \N__23834\ : std_logic;
signal \N__23833\ : std_logic;
signal \N__23832\ : std_logic;
signal \N__23831\ : std_logic;
signal \N__23830\ : std_logic;
signal \N__23829\ : std_logic;
signal \N__23824\ : std_logic;
signal \N__23823\ : std_logic;
signal \N__23822\ : std_logic;
signal \N__23821\ : std_logic;
signal \N__23820\ : std_logic;
signal \N__23815\ : std_logic;
signal \N__23810\ : std_logic;
signal \N__23809\ : std_logic;
signal \N__23804\ : std_logic;
signal \N__23801\ : std_logic;
signal \N__23798\ : std_logic;
signal \N__23793\ : std_logic;
signal \N__23790\ : std_logic;
signal \N__23787\ : std_logic;
signal \N__23782\ : std_logic;
signal \N__23779\ : std_logic;
signal \N__23762\ : std_logic;
signal \N__23759\ : std_logic;
signal \N__23756\ : std_logic;
signal \N__23755\ : std_logic;
signal \N__23754\ : std_logic;
signal \N__23753\ : std_logic;
signal \N__23750\ : std_logic;
signal \N__23749\ : std_logic;
signal \N__23748\ : std_logic;
signal \N__23743\ : std_logic;
signal \N__23742\ : std_logic;
signal \N__23741\ : std_logic;
signal \N__23740\ : std_logic;
signal \N__23739\ : std_logic;
signal \N__23738\ : std_logic;
signal \N__23735\ : std_logic;
signal \N__23730\ : std_logic;
signal \N__23729\ : std_logic;
signal \N__23728\ : std_logic;
signal \N__23727\ : std_logic;
signal \N__23724\ : std_logic;
signal \N__23721\ : std_logic;
signal \N__23718\ : std_logic;
signal \N__23715\ : std_logic;
signal \N__23712\ : std_logic;
signal \N__23709\ : std_logic;
signal \N__23708\ : std_logic;
signal \N__23707\ : std_logic;
signal \N__23706\ : std_logic;
signal \N__23705\ : std_logic;
signal \N__23704\ : std_logic;
signal \N__23703\ : std_logic;
signal \N__23700\ : std_logic;
signal \N__23695\ : std_logic;
signal \N__23690\ : std_logic;
signal \N__23685\ : std_logic;
signal \N__23682\ : std_logic;
signal \N__23679\ : std_logic;
signal \N__23672\ : std_logic;
signal \N__23667\ : std_logic;
signal \N__23664\ : std_logic;
signal \N__23661\ : std_logic;
signal \N__23656\ : std_logic;
signal \N__23647\ : std_logic;
signal \N__23630\ : std_logic;
signal \N__23629\ : std_logic;
signal \N__23626\ : std_logic;
signal \N__23625\ : std_logic;
signal \N__23624\ : std_logic;
signal \N__23623\ : std_logic;
signal \N__23622\ : std_logic;
signal \N__23621\ : std_logic;
signal \N__23620\ : std_logic;
signal \N__23619\ : std_logic;
signal \N__23618\ : std_logic;
signal \N__23617\ : std_logic;
signal \N__23614\ : std_logic;
signal \N__23613\ : std_logic;
signal \N__23612\ : std_logic;
signal \N__23609\ : std_logic;
signal \N__23608\ : std_logic;
signal \N__23607\ : std_logic;
signal \N__23604\ : std_logic;
signal \N__23603\ : std_logic;
signal \N__23600\ : std_logic;
signal \N__23599\ : std_logic;
signal \N__23598\ : std_logic;
signal \N__23595\ : std_logic;
signal \N__23594\ : std_logic;
signal \N__23593\ : std_logic;
signal \N__23592\ : std_logic;
signal \N__23591\ : std_logic;
signal \N__23590\ : std_logic;
signal \N__23589\ : std_logic;
signal \N__23588\ : std_logic;
signal \N__23583\ : std_logic;
signal \N__23574\ : std_logic;
signal \N__23571\ : std_logic;
signal \N__23566\ : std_logic;
signal \N__23563\ : std_logic;
signal \N__23558\ : std_logic;
signal \N__23553\ : std_logic;
signal \N__23550\ : std_logic;
signal \N__23545\ : std_logic;
signal \N__23540\ : std_logic;
signal \N__23533\ : std_logic;
signal \N__23526\ : std_logic;
signal \N__23519\ : std_logic;
signal \N__23498\ : std_logic;
signal \N__23497\ : std_logic;
signal \N__23496\ : std_logic;
signal \N__23495\ : std_logic;
signal \N__23494\ : std_logic;
signal \N__23491\ : std_logic;
signal \N__23490\ : std_logic;
signal \N__23489\ : std_logic;
signal \N__23488\ : std_logic;
signal \N__23485\ : std_logic;
signal \N__23484\ : std_logic;
signal \N__23483\ : std_logic;
signal \N__23482\ : std_logic;
signal \N__23479\ : std_logic;
signal \N__23476\ : std_logic;
signal \N__23475\ : std_logic;
signal \N__23474\ : std_logic;
signal \N__23471\ : std_logic;
signal \N__23468\ : std_logic;
signal \N__23465\ : std_logic;
signal \N__23462\ : std_logic;
signal \N__23459\ : std_logic;
signal \N__23456\ : std_logic;
signal \N__23455\ : std_logic;
signal \N__23452\ : std_logic;
signal \N__23449\ : std_logic;
signal \N__23446\ : std_logic;
signal \N__23445\ : std_logic;
signal \N__23442\ : std_logic;
signal \N__23439\ : std_logic;
signal \N__23436\ : std_logic;
signal \N__23433\ : std_logic;
signal \N__23430\ : std_logic;
signal \N__23427\ : std_logic;
signal \N__23420\ : std_logic;
signal \N__23417\ : std_logic;
signal \N__23412\ : std_logic;
signal \N__23409\ : std_logic;
signal \N__23406\ : std_logic;
signal \N__23403\ : std_logic;
signal \N__23398\ : std_logic;
signal \N__23395\ : std_logic;
signal \N__23392\ : std_logic;
signal \N__23379\ : std_logic;
signal \N__23366\ : std_logic;
signal \N__23365\ : std_logic;
signal \N__23362\ : std_logic;
signal \N__23359\ : std_logic;
signal \N__23354\ : std_logic;
signal \N__23351\ : std_logic;
signal \N__23348\ : std_logic;
signal \N__23347\ : std_logic;
signal \N__23346\ : std_logic;
signal \N__23345\ : std_logic;
signal \N__23344\ : std_logic;
signal \N__23343\ : std_logic;
signal \N__23342\ : std_logic;
signal \N__23341\ : std_logic;
signal \N__23336\ : std_logic;
signal \N__23333\ : std_logic;
signal \N__23330\ : std_logic;
signal \N__23327\ : std_logic;
signal \N__23324\ : std_logic;
signal \N__23321\ : std_logic;
signal \N__23320\ : std_logic;
signal \N__23317\ : std_logic;
signal \N__23316\ : std_logic;
signal \N__23315\ : std_logic;
signal \N__23314\ : std_logic;
signal \N__23313\ : std_logic;
signal \N__23310\ : std_logic;
signal \N__23305\ : std_logic;
signal \N__23302\ : std_logic;
signal \N__23301\ : std_logic;
signal \N__23296\ : std_logic;
signal \N__23295\ : std_logic;
signal \N__23294\ : std_logic;
signal \N__23291\ : std_logic;
signal \N__23286\ : std_logic;
signal \N__23285\ : std_logic;
signal \N__23282\ : std_logic;
signal \N__23279\ : std_logic;
signal \N__23276\ : std_logic;
signal \N__23271\ : std_logic;
signal \N__23268\ : std_logic;
signal \N__23265\ : std_logic;
signal \N__23262\ : std_logic;
signal \N__23255\ : std_logic;
signal \N__23252\ : std_logic;
signal \N__23249\ : std_logic;
signal \N__23238\ : std_logic;
signal \N__23225\ : std_logic;
signal \N__23222\ : std_logic;
signal \N__23219\ : std_logic;
signal \N__23218\ : std_logic;
signal \N__23217\ : std_logic;
signal \N__23216\ : std_logic;
signal \N__23215\ : std_logic;
signal \N__23212\ : std_logic;
signal \N__23211\ : std_logic;
signal \N__23210\ : std_logic;
signal \N__23207\ : std_logic;
signal \N__23206\ : std_logic;
signal \N__23203\ : std_logic;
signal \N__23202\ : std_logic;
signal \N__23201\ : std_logic;
signal \N__23200\ : std_logic;
signal \N__23199\ : std_logic;
signal \N__23196\ : std_logic;
signal \N__23195\ : std_logic;
signal \N__23192\ : std_logic;
signal \N__23185\ : std_logic;
signal \N__23182\ : std_logic;
signal \N__23177\ : std_logic;
signal \N__23176\ : std_logic;
signal \N__23175\ : std_logic;
signal \N__23174\ : std_logic;
signal \N__23173\ : std_logic;
signal \N__23168\ : std_logic;
signal \N__23167\ : std_logic;
signal \N__23166\ : std_logic;
signal \N__23163\ : std_logic;
signal \N__23158\ : std_logic;
signal \N__23153\ : std_logic;
signal \N__23152\ : std_logic;
signal \N__23149\ : std_logic;
signal \N__23144\ : std_logic;
signal \N__23135\ : std_logic;
signal \N__23134\ : std_logic;
signal \N__23131\ : std_logic;
signal \N__23126\ : std_logic;
signal \N__23119\ : std_logic;
signal \N__23116\ : std_logic;
signal \N__23113\ : std_logic;
signal \N__23110\ : std_logic;
signal \N__23107\ : std_logic;
signal \N__23104\ : std_logic;
signal \N__23097\ : std_logic;
signal \N__23084\ : std_logic;
signal \N__23083\ : std_logic;
signal \N__23082\ : std_logic;
signal \N__23081\ : std_logic;
signal \N__23078\ : std_logic;
signal \N__23077\ : std_logic;
signal \N__23076\ : std_logic;
signal \N__23071\ : std_logic;
signal \N__23068\ : std_logic;
signal \N__23065\ : std_logic;
signal \N__23064\ : std_logic;
signal \N__23063\ : std_logic;
signal \N__23060\ : std_logic;
signal \N__23059\ : std_logic;
signal \N__23058\ : std_logic;
signal \N__23055\ : std_logic;
signal \N__23054\ : std_logic;
signal \N__23051\ : std_logic;
signal \N__23048\ : std_logic;
signal \N__23045\ : std_logic;
signal \N__23038\ : std_logic;
signal \N__23037\ : std_logic;
signal \N__23036\ : std_logic;
signal \N__23029\ : std_logic;
signal \N__23028\ : std_logic;
signal \N__23027\ : std_logic;
signal \N__23024\ : std_logic;
signal \N__23023\ : std_logic;
signal \N__23022\ : std_logic;
signal \N__23021\ : std_logic;
signal \N__23012\ : std_logic;
signal \N__23007\ : std_logic;
signal \N__23004\ : std_logic;
signal \N__22997\ : std_logic;
signal \N__22996\ : std_logic;
signal \N__22991\ : std_logic;
signal \N__22988\ : std_logic;
signal \N__22985\ : std_logic;
signal \N__22982\ : std_logic;
signal \N__22977\ : std_logic;
signal \N__22974\ : std_logic;
signal \N__22969\ : std_logic;
signal \N__22966\ : std_logic;
signal \N__22961\ : std_logic;
signal \N__22952\ : std_logic;
signal \N__22951\ : std_logic;
signal \N__22950\ : std_logic;
signal \N__22949\ : std_logic;
signal \N__22948\ : std_logic;
signal \N__22947\ : std_logic;
signal \N__22946\ : std_logic;
signal \N__22945\ : std_logic;
signal \N__22928\ : std_logic;
signal \N__22925\ : std_logic;
signal \N__22922\ : std_logic;
signal \N__22921\ : std_logic;
signal \N__22920\ : std_logic;
signal \N__22919\ : std_logic;
signal \N__22918\ : std_logic;
signal \N__22917\ : std_logic;
signal \N__22916\ : std_logic;
signal \N__22915\ : std_logic;
signal \N__22914\ : std_logic;
signal \N__22913\ : std_logic;
signal \N__22912\ : std_logic;
signal \N__22911\ : std_logic;
signal \N__22910\ : std_logic;
signal \N__22909\ : std_logic;
signal \N__22908\ : std_logic;
signal \N__22907\ : std_logic;
signal \N__22906\ : std_logic;
signal \N__22905\ : std_logic;
signal \N__22904\ : std_logic;
signal \N__22903\ : std_logic;
signal \N__22902\ : std_logic;
signal \N__22901\ : std_logic;
signal \N__22900\ : std_logic;
signal \N__22899\ : std_logic;
signal \N__22898\ : std_logic;
signal \N__22897\ : std_logic;
signal \N__22896\ : std_logic;
signal \N__22895\ : std_logic;
signal \N__22894\ : std_logic;
signal \N__22893\ : std_logic;
signal \N__22892\ : std_logic;
signal \N__22891\ : std_logic;
signal \N__22890\ : std_logic;
signal \N__22889\ : std_logic;
signal \N__22888\ : std_logic;
signal \N__22887\ : std_logic;
signal \N__22886\ : std_logic;
signal \N__22885\ : std_logic;
signal \N__22884\ : std_logic;
signal \N__22883\ : std_logic;
signal \N__22882\ : std_logic;
signal \N__22881\ : std_logic;
signal \N__22880\ : std_logic;
signal \N__22879\ : std_logic;
signal \N__22878\ : std_logic;
signal \N__22877\ : std_logic;
signal \N__22876\ : std_logic;
signal \N__22875\ : std_logic;
signal \N__22778\ : std_logic;
signal \N__22775\ : std_logic;
signal \N__22772\ : std_logic;
signal \N__22769\ : std_logic;
signal \N__22766\ : std_logic;
signal \N__22763\ : std_logic;
signal \N__22760\ : std_logic;
signal \N__22757\ : std_logic;
signal \N__22754\ : std_logic;
signal \N__22751\ : std_logic;
signal \N__22750\ : std_logic;
signal \N__22749\ : std_logic;
signal \N__22748\ : std_logic;
signal \N__22747\ : std_logic;
signal \N__22746\ : std_logic;
signal \N__22743\ : std_logic;
signal \N__22740\ : std_logic;
signal \N__22737\ : std_logic;
signal \N__22734\ : std_logic;
signal \N__22733\ : std_logic;
signal \N__22730\ : std_logic;
signal \N__22727\ : std_logic;
signal \N__22724\ : std_logic;
signal \N__22715\ : std_logic;
signal \N__22710\ : std_logic;
signal \N__22709\ : std_logic;
signal \N__22708\ : std_logic;
signal \N__22705\ : std_logic;
signal \N__22700\ : std_logic;
signal \N__22699\ : std_logic;
signal \N__22698\ : std_logic;
signal \N__22695\ : std_logic;
signal \N__22694\ : std_logic;
signal \N__22691\ : std_logic;
signal \N__22690\ : std_logic;
signal \N__22689\ : std_logic;
signal \N__22686\ : std_logic;
signal \N__22683\ : std_logic;
signal \N__22680\ : std_logic;
signal \N__22679\ : std_logic;
signal \N__22676\ : std_logic;
signal \N__22673\ : std_logic;
signal \N__22670\ : std_logic;
signal \N__22667\ : std_logic;
signal \N__22664\ : std_logic;
signal \N__22661\ : std_logic;
signal \N__22658\ : std_logic;
signal \N__22655\ : std_logic;
signal \N__22650\ : std_logic;
signal \N__22647\ : std_logic;
signal \N__22642\ : std_logic;
signal \N__22637\ : std_logic;
signal \N__22634\ : std_logic;
signal \N__22631\ : std_logic;
signal \N__22624\ : std_logic;
signal \N__22621\ : std_logic;
signal \N__22618\ : std_logic;
signal \N__22607\ : std_logic;
signal \N__22606\ : std_logic;
signal \N__22605\ : std_logic;
signal \N__22602\ : std_logic;
signal \N__22599\ : std_logic;
signal \N__22598\ : std_logic;
signal \N__22597\ : std_logic;
signal \N__22596\ : std_logic;
signal \N__22595\ : std_logic;
signal \N__22594\ : std_logic;
signal \N__22593\ : std_logic;
signal \N__22590\ : std_logic;
signal \N__22589\ : std_logic;
signal \N__22588\ : std_logic;
signal \N__22587\ : std_logic;
signal \N__22582\ : std_logic;
signal \N__22579\ : std_logic;
signal \N__22578\ : std_logic;
signal \N__22577\ : std_logic;
signal \N__22574\ : std_logic;
signal \N__22573\ : std_logic;
signal \N__22572\ : std_logic;
signal \N__22571\ : std_logic;
signal \N__22570\ : std_logic;
signal \N__22569\ : std_logic;
signal \N__22566\ : std_logic;
signal \N__22565\ : std_logic;
signal \N__22564\ : std_logic;
signal \N__22563\ : std_logic;
signal \N__22562\ : std_logic;
signal \N__22561\ : std_logic;
signal \N__22558\ : std_logic;
signal \N__22555\ : std_logic;
signal \N__22554\ : std_logic;
signal \N__22551\ : std_logic;
signal \N__22550\ : std_logic;
signal \N__22547\ : std_logic;
signal \N__22544\ : std_logic;
signal \N__22541\ : std_logic;
signal \N__22538\ : std_logic;
signal \N__22533\ : std_logic;
signal \N__22530\ : std_logic;
signal \N__22527\ : std_logic;
signal \N__22524\ : std_logic;
signal \N__22521\ : std_logic;
signal \N__22518\ : std_logic;
signal \N__22517\ : std_logic;
signal \N__22516\ : std_logic;
signal \N__22515\ : std_logic;
signal \N__22514\ : std_logic;
signal \N__22511\ : std_logic;
signal \N__22510\ : std_logic;
signal \N__22509\ : std_logic;
signal \N__22506\ : std_logic;
signal \N__22503\ : std_logic;
signal \N__22502\ : std_logic;
signal \N__22501\ : std_logic;
signal \N__22500\ : std_logic;
signal \N__22497\ : std_logic;
signal \N__22496\ : std_logic;
signal \N__22493\ : std_logic;
signal \N__22490\ : std_logic;
signal \N__22487\ : std_logic;
signal \N__22484\ : std_logic;
signal \N__22483\ : std_logic;
signal \N__22482\ : std_logic;
signal \N__22481\ : std_logic;
signal \N__22480\ : std_logic;
signal \N__22477\ : std_logic;
signal \N__22472\ : std_logic;
signal \N__22469\ : std_logic;
signal \N__22468\ : std_logic;
signal \N__22465\ : std_logic;
signal \N__22462\ : std_logic;
signal \N__22461\ : std_logic;
signal \N__22456\ : std_logic;
signal \N__22455\ : std_logic;
signal \N__22454\ : std_logic;
signal \N__22453\ : std_logic;
signal \N__22448\ : std_logic;
signal \N__22447\ : std_logic;
signal \N__22444\ : std_logic;
signal \N__22439\ : std_logic;
signal \N__22432\ : std_logic;
signal \N__22429\ : std_logic;
signal \N__22426\ : std_logic;
signal \N__22423\ : std_logic;
signal \N__22420\ : std_logic;
signal \N__22419\ : std_logic;
signal \N__22416\ : std_logic;
signal \N__22413\ : std_logic;
signal \N__22412\ : std_logic;
signal \N__22411\ : std_logic;
signal \N__22410\ : std_logic;
signal \N__22407\ : std_logic;
signal \N__22406\ : std_logic;
signal \N__22405\ : std_logic;
signal \N__22402\ : std_logic;
signal \N__22399\ : std_logic;
signal \N__22396\ : std_logic;
signal \N__22393\ : std_logic;
signal \N__22392\ : std_logic;
signal \N__22389\ : std_logic;
signal \N__22388\ : std_logic;
signal \N__22385\ : std_logic;
signal \N__22382\ : std_logic;
signal \N__22381\ : std_logic;
signal \N__22380\ : std_logic;
signal \N__22377\ : std_logic;
signal \N__22374\ : std_logic;
signal \N__22371\ : std_logic;
signal \N__22368\ : std_logic;
signal \N__22365\ : std_logic;
signal \N__22362\ : std_logic;
signal \N__22359\ : std_logic;
signal \N__22356\ : std_logic;
signal \N__22355\ : std_logic;
signal \N__22354\ : std_logic;
signal \N__22353\ : std_logic;
signal \N__22352\ : std_logic;
signal \N__22351\ : std_logic;
signal \N__22348\ : std_logic;
signal \N__22343\ : std_logic;
signal \N__22340\ : std_logic;
signal \N__22335\ : std_logic;
signal \N__22332\ : std_logic;
signal \N__22329\ : std_logic;
signal \N__22326\ : std_logic;
signal \N__22323\ : std_logic;
signal \N__22320\ : std_logic;
signal \N__22319\ : std_logic;
signal \N__22318\ : std_logic;
signal \N__22315\ : std_logic;
signal \N__22312\ : std_logic;
signal \N__22297\ : std_logic;
signal \N__22294\ : std_logic;
signal \N__22291\ : std_logic;
signal \N__22288\ : std_logic;
signal \N__22285\ : std_logic;
signal \N__22282\ : std_logic;
signal \N__22281\ : std_logic;
signal \N__22280\ : std_logic;
signal \N__22277\ : std_logic;
signal \N__22274\ : std_logic;
signal \N__22271\ : std_logic;
signal \N__22268\ : std_logic;
signal \N__22267\ : std_logic;
signal \N__22264\ : std_logic;
signal \N__22263\ : std_logic;
signal \N__22256\ : std_logic;
signal \N__22253\ : std_logic;
signal \N__22252\ : std_logic;
signal \N__22251\ : std_logic;
signal \N__22248\ : std_logic;
signal \N__22245\ : std_logic;
signal \N__22244\ : std_logic;
signal \N__22243\ : std_logic;
signal \N__22242\ : std_logic;
signal \N__22237\ : std_logic;
signal \N__22234\ : std_logic;
signal \N__22231\ : std_logic;
signal \N__22230\ : std_logic;
signal \N__22219\ : std_logic;
signal \N__22216\ : std_logic;
signal \N__22213\ : std_logic;
signal \N__22210\ : std_logic;
signal \N__22207\ : std_logic;
signal \N__22204\ : std_logic;
signal \N__22201\ : std_logic;
signal \N__22198\ : std_logic;
signal \N__22195\ : std_logic;
signal \N__22188\ : std_logic;
signal \N__22187\ : std_logic;
signal \N__22182\ : std_logic;
signal \N__22177\ : std_logic;
signal \N__22174\ : std_logic;
signal \N__22171\ : std_logic;
signal \N__22168\ : std_logic;
signal \N__22165\ : std_logic;
signal \N__22162\ : std_logic;
signal \N__22155\ : std_logic;
signal \N__22150\ : std_logic;
signal \N__22145\ : std_logic;
signal \N__22142\ : std_logic;
signal \N__22139\ : std_logic;
signal \N__22136\ : std_logic;
signal \N__22129\ : std_logic;
signal \N__22126\ : std_logic;
signal \N__22123\ : std_logic;
signal \N__22120\ : std_logic;
signal \N__22115\ : std_logic;
signal \N__22114\ : std_logic;
signal \N__22111\ : std_logic;
signal \N__22108\ : std_logic;
signal \N__22103\ : std_logic;
signal \N__22102\ : std_logic;
signal \N__22099\ : std_logic;
signal \N__22096\ : std_logic;
signal \N__22093\ : std_logic;
signal \N__22090\ : std_logic;
signal \N__22085\ : std_logic;
signal \N__22084\ : std_logic;
signal \N__22083\ : std_logic;
signal \N__22082\ : std_logic;
signal \N__22081\ : std_logic;
signal \N__22078\ : std_logic;
signal \N__22075\ : std_logic;
signal \N__22072\ : std_logic;
signal \N__22069\ : std_logic;
signal \N__22064\ : std_logic;
signal \N__22053\ : std_logic;
signal \N__22050\ : std_logic;
signal \N__22047\ : std_logic;
signal \N__22044\ : std_logic;
signal \N__22035\ : std_logic;
signal \N__22030\ : std_logic;
signal \N__22021\ : std_logic;
signal \N__22014\ : std_logic;
signal \N__22009\ : std_logic;
signal \N__22006\ : std_logic;
signal \N__22003\ : std_logic;
signal \N__21998\ : std_logic;
signal \N__21995\ : std_logic;
signal \N__21992\ : std_logic;
signal \N__21989\ : std_logic;
signal \N__21986\ : std_logic;
signal \N__21983\ : std_logic;
signal \N__21978\ : std_logic;
signal \N__21975\ : std_logic;
signal \N__21972\ : std_logic;
signal \N__21971\ : std_logic;
signal \N__21968\ : std_logic;
signal \N__21965\ : std_logic;
signal \N__21964\ : std_logic;
signal \N__21961\ : std_logic;
signal \N__21948\ : std_logic;
signal \N__21947\ : std_logic;
signal \N__21946\ : std_logic;
signal \N__21945\ : std_logic;
signal \N__21940\ : std_logic;
signal \N__21937\ : std_logic;
signal \N__21932\ : std_logic;
signal \N__21923\ : std_logic;
signal \N__21916\ : std_logic;
signal \N__21905\ : std_logic;
signal \N__21902\ : std_logic;
signal \N__21899\ : std_logic;
signal \N__21894\ : std_logic;
signal \N__21891\ : std_logic;
signal \N__21890\ : std_logic;
signal \N__21885\ : std_logic;
signal \N__21884\ : std_logic;
signal \N__21881\ : std_logic;
signal \N__21878\ : std_logic;
signal \N__21875\ : std_logic;
signal \N__21874\ : std_logic;
signal \N__21871\ : std_logic;
signal \N__21866\ : std_logic;
signal \N__21861\ : std_logic;
signal \N__21850\ : std_logic;
signal \N__21847\ : std_logic;
signal \N__21844\ : std_logic;
signal \N__21841\ : std_logic;
signal \N__21838\ : std_logic;
signal \N__21833\ : std_logic;
signal \N__21830\ : std_logic;
signal \N__21827\ : std_logic;
signal \N__21824\ : std_logic;
signal \N__21821\ : std_logic;
signal \N__21818\ : std_logic;
signal \N__21811\ : std_logic;
signal \N__21804\ : std_logic;
signal \N__21801\ : std_logic;
signal \N__21798\ : std_logic;
signal \N__21793\ : std_logic;
signal \N__21788\ : std_logic;
signal \N__21785\ : std_logic;
signal \N__21782\ : std_logic;
signal \N__21779\ : std_logic;
signal \N__21776\ : std_logic;
signal \N__21767\ : std_logic;
signal \N__21766\ : std_logic;
signal \N__21763\ : std_logic;
signal \N__21760\ : std_logic;
signal \N__21757\ : std_logic;
signal \N__21752\ : std_logic;
signal \N__21749\ : std_logic;
signal \N__21748\ : std_logic;
signal \N__21747\ : std_logic;
signal \N__21742\ : std_logic;
signal \N__21739\ : std_logic;
signal \N__21734\ : std_logic;
signal \N__21733\ : std_logic;
signal \N__21732\ : std_logic;
signal \N__21729\ : std_logic;
signal \N__21726\ : std_logic;
signal \N__21725\ : std_logic;
signal \N__21724\ : std_logic;
signal \N__21723\ : std_logic;
signal \N__21720\ : std_logic;
signal \N__21715\ : std_logic;
signal \N__21712\ : std_logic;
signal \N__21709\ : std_logic;
signal \N__21706\ : std_logic;
signal \N__21695\ : std_logic;
signal \N__21694\ : std_logic;
signal \N__21693\ : std_logic;
signal \N__21692\ : std_logic;
signal \N__21691\ : std_logic;
signal \N__21690\ : std_logic;
signal \N__21689\ : std_logic;
signal \N__21686\ : std_logic;
signal \N__21681\ : std_logic;
signal \N__21678\ : std_logic;
signal \N__21675\ : std_logic;
signal \N__21670\ : std_logic;
signal \N__21667\ : std_logic;
signal \N__21666\ : std_logic;
signal \N__21663\ : std_logic;
signal \N__21662\ : std_logic;
signal \N__21661\ : std_logic;
signal \N__21660\ : std_logic;
signal \N__21659\ : std_logic;
signal \N__21658\ : std_logic;
signal \N__21657\ : std_logic;
signal \N__21656\ : std_logic;
signal \N__21653\ : std_logic;
signal \N__21650\ : std_logic;
signal \N__21647\ : std_logic;
signal \N__21644\ : std_logic;
signal \N__21643\ : std_logic;
signal \N__21640\ : std_logic;
signal \N__21639\ : std_logic;
signal \N__21636\ : std_logic;
signal \N__21633\ : std_logic;
signal \N__21626\ : std_logic;
signal \N__21623\ : std_logic;
signal \N__21620\ : std_logic;
signal \N__21617\ : std_logic;
signal \N__21612\ : std_logic;
signal \N__21607\ : std_logic;
signal \N__21600\ : std_logic;
signal \N__21581\ : std_logic;
signal \N__21578\ : std_logic;
signal \N__21575\ : std_logic;
signal \N__21572\ : std_logic;
signal \N__21569\ : std_logic;
signal \N__21566\ : std_logic;
signal \N__21563\ : std_logic;
signal \N__21562\ : std_logic;
signal \N__21561\ : std_logic;
signal \N__21560\ : std_logic;
signal \N__21559\ : std_logic;
signal \N__21556\ : std_logic;
signal \N__21553\ : std_logic;
signal \N__21552\ : std_logic;
signal \N__21549\ : std_logic;
signal \N__21544\ : std_logic;
signal \N__21543\ : std_logic;
signal \N__21542\ : std_logic;
signal \N__21539\ : std_logic;
signal \N__21534\ : std_logic;
signal \N__21533\ : std_logic;
signal \N__21532\ : std_logic;
signal \N__21531\ : std_logic;
signal \N__21530\ : std_logic;
signal \N__21529\ : std_logic;
signal \N__21528\ : std_logic;
signal \N__21527\ : std_logic;
signal \N__21522\ : std_logic;
signal \N__21517\ : std_logic;
signal \N__21512\ : std_logic;
signal \N__21507\ : std_logic;
signal \N__21500\ : std_logic;
signal \N__21495\ : std_logic;
signal \N__21482\ : std_logic;
signal \N__21479\ : std_logic;
signal \N__21478\ : std_logic;
signal \N__21477\ : std_logic;
signal \N__21476\ : std_logic;
signal \N__21473\ : std_logic;
signal \N__21468\ : std_logic;
signal \N__21467\ : std_logic;
signal \N__21464\ : std_logic;
signal \N__21463\ : std_logic;
signal \N__21462\ : std_logic;
signal \N__21457\ : std_logic;
signal \N__21456\ : std_logic;
signal \N__21455\ : std_logic;
signal \N__21454\ : std_logic;
signal \N__21453\ : std_logic;
signal \N__21450\ : std_logic;
signal \N__21445\ : std_logic;
signal \N__21444\ : std_logic;
signal \N__21443\ : std_logic;
signal \N__21440\ : std_logic;
signal \N__21439\ : std_logic;
signal \N__21436\ : std_logic;
signal \N__21431\ : std_logic;
signal \N__21426\ : std_logic;
signal \N__21421\ : std_logic;
signal \N__21416\ : std_logic;
signal \N__21411\ : std_logic;
signal \N__21404\ : std_logic;
signal \N__21395\ : std_logic;
signal \N__21392\ : std_logic;
signal \N__21389\ : std_logic;
signal \N__21386\ : std_logic;
signal \N__21383\ : std_logic;
signal \N__21380\ : std_logic;
signal \N__21377\ : std_logic;
signal \N__21374\ : std_logic;
signal \N__21371\ : std_logic;
signal \N__21368\ : std_logic;
signal \N__21365\ : std_logic;
signal \N__21362\ : std_logic;
signal \N__21359\ : std_logic;
signal \N__21356\ : std_logic;
signal \N__21355\ : std_logic;
signal \N__21354\ : std_logic;
signal \N__21353\ : std_logic;
signal \N__21352\ : std_logic;
signal \N__21351\ : std_logic;
signal \N__21348\ : std_logic;
signal \N__21345\ : std_logic;
signal \N__21342\ : std_logic;
signal \N__21339\ : std_logic;
signal \N__21336\ : std_logic;
signal \N__21333\ : std_logic;
signal \N__21330\ : std_logic;
signal \N__21327\ : std_logic;
signal \N__21324\ : std_logic;
signal \N__21311\ : std_logic;
signal \N__21310\ : std_logic;
signal \N__21305\ : std_logic;
signal \N__21302\ : std_logic;
signal \N__21299\ : std_logic;
signal \N__21296\ : std_logic;
signal \N__21293\ : std_logic;
signal \N__21290\ : std_logic;
signal \N__21287\ : std_logic;
signal \N__21284\ : std_logic;
signal \N__21281\ : std_logic;
signal \N__21278\ : std_logic;
signal \N__21275\ : std_logic;
signal \N__21272\ : std_logic;
signal \N__21269\ : std_logic;
signal \N__21266\ : std_logic;
signal \N__21265\ : std_logic;
signal \N__21262\ : std_logic;
signal \N__21261\ : std_logic;
signal \N__21258\ : std_logic;
signal \N__21255\ : std_logic;
signal \N__21252\ : std_logic;
signal \N__21251\ : std_logic;
signal \N__21248\ : std_logic;
signal \N__21243\ : std_logic;
signal \N__21240\ : std_logic;
signal \N__21233\ : std_logic;
signal \N__21232\ : std_logic;
signal \N__21229\ : std_logic;
signal \N__21226\ : std_logic;
signal \N__21225\ : std_logic;
signal \N__21224\ : std_logic;
signal \N__21223\ : std_logic;
signal \N__21222\ : std_logic;
signal \N__21221\ : std_logic;
signal \N__21220\ : std_logic;
signal \N__21215\ : std_logic;
signal \N__21210\ : std_logic;
signal \N__21207\ : std_logic;
signal \N__21206\ : std_logic;
signal \N__21205\ : std_logic;
signal \N__21204\ : std_logic;
signal \N__21197\ : std_logic;
signal \N__21190\ : std_logic;
signal \N__21183\ : std_logic;
signal \N__21176\ : std_logic;
signal \N__21175\ : std_logic;
signal \N__21174\ : std_logic;
signal \N__21173\ : std_logic;
signal \N__21172\ : std_logic;
signal \N__21165\ : std_logic;
signal \N__21162\ : std_logic;
signal \N__21159\ : std_logic;
signal \N__21158\ : std_logic;
signal \N__21157\ : std_logic;
signal \N__21156\ : std_logic;
signal \N__21155\ : std_logic;
signal \N__21152\ : std_logic;
signal \N__21147\ : std_logic;
signal \N__21146\ : std_logic;
signal \N__21145\ : std_logic;
signal \N__21142\ : std_logic;
signal \N__21135\ : std_logic;
signal \N__21134\ : std_logic;
signal \N__21133\ : std_logic;
signal \N__21128\ : std_logic;
signal \N__21125\ : std_logic;
signal \N__21122\ : std_logic;
signal \N__21119\ : std_logic;
signal \N__21116\ : std_logic;
signal \N__21111\ : std_logic;
signal \N__21106\ : std_logic;
signal \N__21095\ : std_logic;
signal \N__21094\ : std_logic;
signal \N__21093\ : std_logic;
signal \N__21092\ : std_logic;
signal \N__21091\ : std_logic;
signal \N__21090\ : std_logic;
signal \N__21087\ : std_logic;
signal \N__21086\ : std_logic;
signal \N__21085\ : std_logic;
signal \N__21084\ : std_logic;
signal \N__21083\ : std_logic;
signal \N__21080\ : std_logic;
signal \N__21077\ : std_logic;
signal \N__21072\ : std_logic;
signal \N__21069\ : std_logic;
signal \N__21066\ : std_logic;
signal \N__21063\ : std_logic;
signal \N__21060\ : std_logic;
signal \N__21059\ : std_logic;
signal \N__21058\ : std_logic;
signal \N__21053\ : std_logic;
signal \N__21046\ : std_logic;
signal \N__21039\ : std_logic;
signal \N__21038\ : std_logic;
signal \N__21035\ : std_logic;
signal \N__21032\ : std_logic;
signal \N__21029\ : std_logic;
signal \N__21024\ : std_logic;
signal \N__21021\ : std_logic;
signal \N__21018\ : std_logic;
signal \N__21005\ : std_logic;
signal \N__21004\ : std_logic;
signal \N__21003\ : std_logic;
signal \N__21002\ : std_logic;
signal \N__20997\ : std_logic;
signal \N__20994\ : std_logic;
signal \N__20991\ : std_logic;
signal \N__20990\ : std_logic;
signal \N__20987\ : std_logic;
signal \N__20984\ : std_logic;
signal \N__20981\ : std_logic;
signal \N__20978\ : std_logic;
signal \N__20975\ : std_logic;
signal \N__20972\ : std_logic;
signal \N__20969\ : std_logic;
signal \N__20966\ : std_logic;
signal \N__20957\ : std_logic;
signal \N__20954\ : std_logic;
signal \N__20953\ : std_logic;
signal \N__20950\ : std_logic;
signal \N__20947\ : std_logic;
signal \N__20944\ : std_logic;
signal \N__20941\ : std_logic;
signal \N__20936\ : std_logic;
signal \N__20935\ : std_logic;
signal \N__20934\ : std_logic;
signal \N__20933\ : std_logic;
signal \N__20932\ : std_logic;
signal \N__20929\ : std_logic;
signal \N__20928\ : std_logic;
signal \N__20927\ : std_logic;
signal \N__20924\ : std_logic;
signal \N__20921\ : std_logic;
signal \N__20918\ : std_logic;
signal \N__20915\ : std_logic;
signal \N__20914\ : std_logic;
signal \N__20913\ : std_logic;
signal \N__20912\ : std_logic;
signal \N__20909\ : std_logic;
signal \N__20906\ : std_logic;
signal \N__20903\ : std_logic;
signal \N__20900\ : std_logic;
signal \N__20899\ : std_logic;
signal \N__20898\ : std_logic;
signal \N__20897\ : std_logic;
signal \N__20890\ : std_logic;
signal \N__20883\ : std_logic;
signal \N__20878\ : std_logic;
signal \N__20873\ : std_logic;
signal \N__20872\ : std_logic;
signal \N__20869\ : std_logic;
signal \N__20868\ : std_logic;
signal \N__20867\ : std_logic;
signal \N__20862\ : std_logic;
signal \N__20857\ : std_logic;
signal \N__20852\ : std_logic;
signal \N__20847\ : std_logic;
signal \N__20842\ : std_logic;
signal \N__20831\ : std_logic;
signal \N__20828\ : std_logic;
signal \N__20827\ : std_logic;
signal \N__20826\ : std_logic;
signal \N__20825\ : std_logic;
signal \N__20824\ : std_logic;
signal \N__20823\ : std_logic;
signal \N__20822\ : std_logic;
signal \N__20815\ : std_logic;
signal \N__20812\ : std_logic;
signal \N__20809\ : std_logic;
signal \N__20804\ : std_logic;
signal \N__20801\ : std_logic;
signal \N__20798\ : std_logic;
signal \N__20797\ : std_logic;
signal \N__20792\ : std_logic;
signal \N__20789\ : std_logic;
signal \N__20786\ : std_logic;
signal \N__20783\ : std_logic;
signal \N__20780\ : std_logic;
signal \N__20777\ : std_logic;
signal \N__20768\ : std_logic;
signal \N__20765\ : std_logic;
signal \N__20764\ : std_logic;
signal \N__20763\ : std_logic;
signal \N__20760\ : std_logic;
signal \N__20757\ : std_logic;
signal \N__20756\ : std_logic;
signal \N__20755\ : std_logic;
signal \N__20754\ : std_logic;
signal \N__20751\ : std_logic;
signal \N__20748\ : std_logic;
signal \N__20745\ : std_logic;
signal \N__20742\ : std_logic;
signal \N__20737\ : std_logic;
signal \N__20734\ : std_logic;
signal \N__20723\ : std_logic;
signal \N__20722\ : std_logic;
signal \N__20719\ : std_logic;
signal \N__20716\ : std_logic;
signal \N__20713\ : std_logic;
signal \N__20712\ : std_logic;
signal \N__20711\ : std_logic;
signal \N__20710\ : std_logic;
signal \N__20707\ : std_logic;
signal \N__20704\ : std_logic;
signal \N__20699\ : std_logic;
signal \N__20696\ : std_logic;
signal \N__20687\ : std_logic;
signal \N__20686\ : std_logic;
signal \N__20685\ : std_logic;
signal \N__20682\ : std_logic;
signal \N__20677\ : std_logic;
signal \N__20674\ : std_logic;
signal \N__20671\ : std_logic;
signal \N__20666\ : std_logic;
signal \N__20665\ : std_logic;
signal \N__20664\ : std_logic;
signal \N__20661\ : std_logic;
signal \N__20658\ : std_logic;
signal \N__20653\ : std_logic;
signal \N__20650\ : std_logic;
signal \N__20647\ : std_logic;
signal \N__20642\ : std_logic;
signal \N__20639\ : std_logic;
signal \N__20638\ : std_logic;
signal \N__20637\ : std_logic;
signal \N__20636\ : std_logic;
signal \N__20635\ : std_logic;
signal \N__20634\ : std_logic;
signal \N__20633\ : std_logic;
signal \N__20632\ : std_logic;
signal \N__20631\ : std_logic;
signal \N__20630\ : std_logic;
signal \N__20627\ : std_logic;
signal \N__20624\ : std_logic;
signal \N__20621\ : std_logic;
signal \N__20618\ : std_logic;
signal \N__20617\ : std_logic;
signal \N__20614\ : std_logic;
signal \N__20611\ : std_logic;
signal \N__20610\ : std_logic;
signal \N__20605\ : std_logic;
signal \N__20604\ : std_logic;
signal \N__20603\ : std_logic;
signal \N__20600\ : std_logic;
signal \N__20597\ : std_logic;
signal \N__20588\ : std_logic;
signal \N__20585\ : std_logic;
signal \N__20580\ : std_logic;
signal \N__20579\ : std_logic;
signal \N__20578\ : std_logic;
signal \N__20577\ : std_logic;
signal \N__20576\ : std_logic;
signal \N__20573\ : std_logic;
signal \N__20570\ : std_logic;
signal \N__20565\ : std_logic;
signal \N__20562\ : std_logic;
signal \N__20561\ : std_logic;
signal \N__20558\ : std_logic;
signal \N__20557\ : std_logic;
signal \N__20550\ : std_logic;
signal \N__20547\ : std_logic;
signal \N__20540\ : std_logic;
signal \N__20531\ : std_logic;
signal \N__20528\ : std_logic;
signal \N__20525\ : std_logic;
signal \N__20522\ : std_logic;
signal \N__20519\ : std_logic;
signal \N__20504\ : std_logic;
signal \N__20503\ : std_logic;
signal \N__20502\ : std_logic;
signal \N__20501\ : std_logic;
signal \N__20500\ : std_logic;
signal \N__20495\ : std_logic;
signal \N__20494\ : std_logic;
signal \N__20493\ : std_logic;
signal \N__20492\ : std_logic;
signal \N__20489\ : std_logic;
signal \N__20486\ : std_logic;
signal \N__20485\ : std_logic;
signal \N__20484\ : std_logic;
signal \N__20483\ : std_logic;
signal \N__20482\ : std_logic;
signal \N__20479\ : std_logic;
signal \N__20478\ : std_logic;
signal \N__20477\ : std_logic;
signal \N__20476\ : std_logic;
signal \N__20473\ : std_logic;
signal \N__20468\ : std_logic;
signal \N__20465\ : std_logic;
signal \N__20462\ : std_logic;
signal \N__20459\ : std_logic;
signal \N__20454\ : std_logic;
signal \N__20453\ : std_logic;
signal \N__20448\ : std_logic;
signal \N__20445\ : std_logic;
signal \N__20442\ : std_logic;
signal \N__20441\ : std_logic;
signal \N__20436\ : std_logic;
signal \N__20425\ : std_logic;
signal \N__20422\ : std_logic;
signal \N__20419\ : std_logic;
signal \N__20416\ : std_logic;
signal \N__20411\ : std_logic;
signal \N__20408\ : std_logic;
signal \N__20407\ : std_logic;
signal \N__20406\ : std_logic;
signal \N__20405\ : std_logic;
signal \N__20404\ : std_logic;
signal \N__20403\ : std_logic;
signal \N__20402\ : std_logic;
signal \N__20399\ : std_logic;
signal \N__20394\ : std_logic;
signal \N__20391\ : std_logic;
signal \N__20384\ : std_logic;
signal \N__20375\ : std_logic;
signal \N__20370\ : std_logic;
signal \N__20367\ : std_logic;
signal \N__20354\ : std_logic;
signal \N__20351\ : std_logic;
signal \N__20348\ : std_logic;
signal \N__20345\ : std_logic;
signal \N__20342\ : std_logic;
signal \N__20339\ : std_logic;
signal \N__20336\ : std_logic;
signal \N__20333\ : std_logic;
signal \N__20332\ : std_logic;
signal \N__20331\ : std_logic;
signal \N__20330\ : std_logic;
signal \N__20329\ : std_logic;
signal \N__20328\ : std_logic;
signal \N__20327\ : std_logic;
signal \N__20326\ : std_logic;
signal \N__20325\ : std_logic;
signal \N__20324\ : std_logic;
signal \N__20323\ : std_logic;
signal \N__20320\ : std_logic;
signal \N__20317\ : std_logic;
signal \N__20312\ : std_logic;
signal \N__20309\ : std_logic;
signal \N__20304\ : std_logic;
signal \N__20299\ : std_logic;
signal \N__20298\ : std_logic;
signal \N__20297\ : std_logic;
signal \N__20296\ : std_logic;
signal \N__20295\ : std_logic;
signal \N__20294\ : std_logic;
signal \N__20291\ : std_logic;
signal \N__20286\ : std_logic;
signal \N__20281\ : std_logic;
signal \N__20278\ : std_logic;
signal \N__20277\ : std_logic;
signal \N__20276\ : std_logic;
signal \N__20271\ : std_logic;
signal \N__20266\ : std_logic;
signal \N__20257\ : std_logic;
signal \N__20254\ : std_logic;
signal \N__20249\ : std_logic;
signal \N__20246\ : std_logic;
signal \N__20243\ : std_logic;
signal \N__20242\ : std_logic;
signal \N__20239\ : std_logic;
signal \N__20234\ : std_logic;
signal \N__20227\ : std_logic;
signal \N__20222\ : std_logic;
signal \N__20213\ : std_logic;
signal \N__20210\ : std_logic;
signal \N__20207\ : std_logic;
signal \N__20204\ : std_logic;
signal \N__20201\ : std_logic;
signal \N__20198\ : std_logic;
signal \N__20195\ : std_logic;
signal \N__20192\ : std_logic;
signal \N__20189\ : std_logic;
signal \N__20186\ : std_logic;
signal \N__20183\ : std_logic;
signal \N__20180\ : std_logic;
signal \N__20179\ : std_logic;
signal \N__20176\ : std_logic;
signal \N__20173\ : std_logic;
signal \N__20168\ : std_logic;
signal \N__20165\ : std_logic;
signal \N__20162\ : std_logic;
signal \N__20159\ : std_logic;
signal \N__20156\ : std_logic;
signal \N__20153\ : std_logic;
signal \N__20150\ : std_logic;
signal \N__20147\ : std_logic;
signal \N__20146\ : std_logic;
signal \N__20143\ : std_logic;
signal \N__20142\ : std_logic;
signal \N__20141\ : std_logic;
signal \N__20140\ : std_logic;
signal \N__20139\ : std_logic;
signal \N__20136\ : std_logic;
signal \N__20133\ : std_logic;
signal \N__20128\ : std_logic;
signal \N__20125\ : std_logic;
signal \N__20124\ : std_logic;
signal \N__20123\ : std_logic;
signal \N__20118\ : std_logic;
signal \N__20117\ : std_logic;
signal \N__20116\ : std_logic;
signal \N__20115\ : std_logic;
signal \N__20114\ : std_logic;
signal \N__20113\ : std_logic;
signal \N__20110\ : std_logic;
signal \N__20107\ : std_logic;
signal \N__20106\ : std_logic;
signal \N__20103\ : std_logic;
signal \N__20098\ : std_logic;
signal \N__20097\ : std_logic;
signal \N__20096\ : std_logic;
signal \N__20095\ : std_logic;
signal \N__20094\ : std_logic;
signal \N__20093\ : std_logic;
signal \N__20090\ : std_logic;
signal \N__20085\ : std_logic;
signal \N__20082\ : std_logic;
signal \N__20077\ : std_logic;
signal \N__20072\ : std_logic;
signal \N__20069\ : std_logic;
signal \N__20064\ : std_logic;
signal \N__20059\ : std_logic;
signal \N__20054\ : std_logic;
signal \N__20051\ : std_logic;
signal \N__20048\ : std_logic;
signal \N__20027\ : std_logic;
signal \N__20024\ : std_logic;
signal \N__20021\ : std_logic;
signal \N__20020\ : std_logic;
signal \N__20019\ : std_logic;
signal \N__20016\ : std_logic;
signal \N__20013\ : std_logic;
signal \N__20010\ : std_logic;
signal \N__20007\ : std_logic;
signal \N__20000\ : std_logic;
signal \N__19997\ : std_logic;
signal \N__19994\ : std_logic;
signal \N__19991\ : std_logic;
signal \N__19988\ : std_logic;
signal \N__19985\ : std_logic;
signal \N__19982\ : std_logic;
signal \N__19979\ : std_logic;
signal \N__19976\ : std_logic;
signal \N__19973\ : std_logic;
signal \N__19970\ : std_logic;
signal \N__19967\ : std_logic;
signal \N__19964\ : std_logic;
signal \N__19963\ : std_logic;
signal \N__19962\ : std_logic;
signal \N__19961\ : std_logic;
signal \N__19952\ : std_logic;
signal \N__19949\ : std_logic;
signal \N__19946\ : std_logic;
signal \N__19943\ : std_logic;
signal \N__19940\ : std_logic;
signal \N__19937\ : std_logic;
signal \N__19934\ : std_logic;
signal \N__19933\ : std_logic;
signal \N__19930\ : std_logic;
signal \N__19927\ : std_logic;
signal \N__19926\ : std_logic;
signal \N__19921\ : std_logic;
signal \N__19920\ : std_logic;
signal \N__19917\ : std_logic;
signal \N__19914\ : std_logic;
signal \N__19911\ : std_logic;
signal \N__19908\ : std_logic;
signal \N__19905\ : std_logic;
signal \N__19900\ : std_logic;
signal \N__19895\ : std_logic;
signal \N__19894\ : std_logic;
signal \N__19891\ : std_logic;
signal \N__19890\ : std_logic;
signal \N__19889\ : std_logic;
signal \N__19886\ : std_logic;
signal \N__19883\ : std_logic;
signal \N__19880\ : std_logic;
signal \N__19877\ : std_logic;
signal \N__19876\ : std_logic;
signal \N__19875\ : std_logic;
signal \N__19874\ : std_logic;
signal \N__19873\ : std_logic;
signal \N__19870\ : std_logic;
signal \N__19869\ : std_logic;
signal \N__19866\ : std_logic;
signal \N__19863\ : std_logic;
signal \N__19862\ : std_logic;
signal \N__19857\ : std_logic;
signal \N__19852\ : std_logic;
signal \N__19849\ : std_logic;
signal \N__19846\ : std_logic;
signal \N__19843\ : std_logic;
signal \N__19838\ : std_logic;
signal \N__19835\ : std_logic;
signal \N__19830\ : std_logic;
signal \N__19817\ : std_logic;
signal \N__19816\ : std_logic;
signal \N__19815\ : std_logic;
signal \N__19812\ : std_logic;
signal \N__19809\ : std_logic;
signal \N__19808\ : std_logic;
signal \N__19807\ : std_logic;
signal \N__19806\ : std_logic;
signal \N__19805\ : std_logic;
signal \N__19804\ : std_logic;
signal \N__19801\ : std_logic;
signal \N__19798\ : std_logic;
signal \N__19795\ : std_logic;
signal \N__19792\ : std_logic;
signal \N__19789\ : std_logic;
signal \N__19786\ : std_logic;
signal \N__19781\ : std_logic;
signal \N__19778\ : std_logic;
signal \N__19773\ : std_logic;
signal \N__19760\ : std_logic;
signal \N__19759\ : std_logic;
signal \N__19758\ : std_logic;
signal \N__19757\ : std_logic;
signal \N__19756\ : std_logic;
signal \N__19755\ : std_logic;
signal \N__19754\ : std_logic;
signal \N__19751\ : std_logic;
signal \N__19744\ : std_logic;
signal \N__19741\ : std_logic;
signal \N__19740\ : std_logic;
signal \N__19735\ : std_logic;
signal \N__19728\ : std_logic;
signal \N__19727\ : std_logic;
signal \N__19726\ : std_logic;
signal \N__19725\ : std_logic;
signal \N__19724\ : std_logic;
signal \N__19723\ : std_logic;
signal \N__19722\ : std_logic;
signal \N__19721\ : std_logic;
signal \N__19718\ : std_logic;
signal \N__19713\ : std_logic;
signal \N__19708\ : std_logic;
signal \N__19703\ : std_logic;
signal \N__19696\ : std_logic;
signal \N__19685\ : std_logic;
signal \N__19682\ : std_logic;
signal \N__19679\ : std_logic;
signal \N__19676\ : std_logic;
signal \N__19673\ : std_logic;
signal \N__19672\ : std_logic;
signal \N__19671\ : std_logic;
signal \N__19668\ : std_logic;
signal \N__19667\ : std_logic;
signal \N__19666\ : std_logic;
signal \N__19665\ : std_logic;
signal \N__19660\ : std_logic;
signal \N__19657\ : std_logic;
signal \N__19656\ : std_logic;
signal \N__19655\ : std_logic;
signal \N__19652\ : std_logic;
signal \N__19649\ : std_logic;
signal \N__19646\ : std_logic;
signal \N__19643\ : std_logic;
signal \N__19640\ : std_logic;
signal \N__19637\ : std_logic;
signal \N__19634\ : std_logic;
signal \N__19631\ : std_logic;
signal \N__19616\ : std_logic;
signal \N__19615\ : std_logic;
signal \N__19614\ : std_logic;
signal \N__19613\ : std_logic;
signal \N__19610\ : std_logic;
signal \N__19607\ : std_logic;
signal \N__19604\ : std_logic;
signal \N__19603\ : std_logic;
signal \N__19598\ : std_logic;
signal \N__19595\ : std_logic;
signal \N__19592\ : std_logic;
signal \N__19589\ : std_logic;
signal \N__19588\ : std_logic;
signal \N__19587\ : std_logic;
signal \N__19584\ : std_logic;
signal \N__19581\ : std_logic;
signal \N__19576\ : std_logic;
signal \N__19573\ : std_logic;
signal \N__19570\ : std_logic;
signal \N__19563\ : std_logic;
signal \N__19556\ : std_logic;
signal \N__19553\ : std_logic;
signal \N__19550\ : std_logic;
signal \N__19549\ : std_logic;
signal \N__19548\ : std_logic;
signal \N__19541\ : std_logic;
signal \N__19538\ : std_logic;
signal \N__19537\ : std_logic;
signal \N__19536\ : std_logic;
signal \N__19533\ : std_logic;
signal \N__19530\ : std_logic;
signal \N__19523\ : std_logic;
signal \N__19520\ : std_logic;
signal \N__19519\ : std_logic;
signal \N__19518\ : std_logic;
signal \N__19517\ : std_logic;
signal \N__19516\ : std_logic;
signal \N__19515\ : std_logic;
signal \N__19514\ : std_logic;
signal \N__19511\ : std_logic;
signal \N__19508\ : std_logic;
signal \N__19505\ : std_logic;
signal \N__19504\ : std_logic;
signal \N__19501\ : std_logic;
signal \N__19498\ : std_logic;
signal \N__19495\ : std_logic;
signal \N__19492\ : std_logic;
signal \N__19489\ : std_logic;
signal \N__19486\ : std_logic;
signal \N__19483\ : std_logic;
signal \N__19478\ : std_logic;
signal \N__19473\ : std_logic;
signal \N__19472\ : std_logic;
signal \N__19469\ : std_logic;
signal \N__19468\ : std_logic;
signal \N__19467\ : std_logic;
signal \N__19466\ : std_logic;
signal \N__19463\ : std_logic;
signal \N__19460\ : std_logic;
signal \N__19455\ : std_logic;
signal \N__19452\ : std_logic;
signal \N__19449\ : std_logic;
signal \N__19446\ : std_logic;
signal \N__19439\ : std_logic;
signal \N__19432\ : std_logic;
signal \N__19429\ : std_logic;
signal \N__19418\ : std_logic;
signal \N__19417\ : std_logic;
signal \N__19416\ : std_logic;
signal \N__19415\ : std_logic;
signal \N__19412\ : std_logic;
signal \N__19411\ : std_logic;
signal \N__19408\ : std_logic;
signal \N__19405\ : std_logic;
signal \N__19402\ : std_logic;
signal \N__19399\ : std_logic;
signal \N__19396\ : std_logic;
signal \N__19385\ : std_logic;
signal \N__19382\ : std_logic;
signal \N__19379\ : std_logic;
signal \N__19376\ : std_logic;
signal \N__19373\ : std_logic;
signal \N__19372\ : std_logic;
signal \N__19369\ : std_logic;
signal \N__19366\ : std_logic;
signal \N__19363\ : std_logic;
signal \N__19362\ : std_logic;
signal \N__19361\ : std_logic;
signal \N__19358\ : std_logic;
signal \N__19357\ : std_logic;
signal \N__19354\ : std_logic;
signal \N__19351\ : std_logic;
signal \N__19348\ : std_logic;
signal \N__19345\ : std_logic;
signal \N__19342\ : std_logic;
signal \N__19331\ : std_logic;
signal \N__19328\ : std_logic;
signal \N__19325\ : std_logic;
signal \N__19322\ : std_logic;
signal \N__19321\ : std_logic;
signal \N__19320\ : std_logic;
signal \N__19319\ : std_logic;
signal \N__19316\ : std_logic;
signal \N__19315\ : std_logic;
signal \N__19312\ : std_logic;
signal \N__19309\ : std_logic;
signal \N__19306\ : std_logic;
signal \N__19303\ : std_logic;
signal \N__19302\ : std_logic;
signal \N__19301\ : std_logic;
signal \N__19296\ : std_logic;
signal \N__19293\ : std_logic;
signal \N__19290\ : std_logic;
signal \N__19287\ : std_logic;
signal \N__19282\ : std_logic;
signal \N__19277\ : std_logic;
signal \N__19274\ : std_logic;
signal \N__19265\ : std_logic;
signal \N__19264\ : std_logic;
signal \N__19261\ : std_logic;
signal \N__19260\ : std_logic;
signal \N__19257\ : std_logic;
signal \N__19256\ : std_logic;
signal \N__19255\ : std_logic;
signal \N__19252\ : std_logic;
signal \N__19249\ : std_logic;
signal \N__19246\ : std_logic;
signal \N__19243\ : std_logic;
signal \N__19240\ : std_logic;
signal \N__19237\ : std_logic;
signal \N__19234\ : std_logic;
signal \N__19229\ : std_logic;
signal \N__19220\ : std_logic;
signal \N__19217\ : std_logic;
signal \N__19214\ : std_logic;
signal \N__19213\ : std_logic;
signal \N__19212\ : std_logic;
signal \N__19209\ : std_logic;
signal \N__19206\ : std_logic;
signal \N__19205\ : std_logic;
signal \N__19202\ : std_logic;
signal \N__19201\ : std_logic;
signal \N__19200\ : std_logic;
signal \N__19199\ : std_logic;
signal \N__19198\ : std_logic;
signal \N__19195\ : std_logic;
signal \N__19192\ : std_logic;
signal \N__19189\ : std_logic;
signal \N__19186\ : std_logic;
signal \N__19181\ : std_logic;
signal \N__19176\ : std_logic;
signal \N__19169\ : std_logic;
signal \N__19160\ : std_logic;
signal \N__19159\ : std_logic;
signal \N__19156\ : std_logic;
signal \N__19153\ : std_logic;
signal \N__19150\ : std_logic;
signal \N__19149\ : std_logic;
signal \N__19146\ : std_logic;
signal \N__19143\ : std_logic;
signal \N__19140\ : std_logic;
signal \N__19137\ : std_logic;
signal \N__19130\ : std_logic;
signal \N__19127\ : std_logic;
signal \N__19126\ : std_logic;
signal \N__19123\ : std_logic;
signal \N__19120\ : std_logic;
signal \N__19119\ : std_logic;
signal \N__19116\ : std_logic;
signal \N__19113\ : std_logic;
signal \N__19112\ : std_logic;
signal \N__19109\ : std_logic;
signal \N__19106\ : std_logic;
signal \N__19103\ : std_logic;
signal \N__19098\ : std_logic;
signal \N__19091\ : std_logic;
signal \N__19088\ : std_logic;
signal \N__19085\ : std_logic;
signal \N__19082\ : std_logic;
signal \N__19081\ : std_logic;
signal \N__19080\ : std_logic;
signal \N__19077\ : std_logic;
signal \N__19076\ : std_logic;
signal \N__19075\ : std_logic;
signal \N__19072\ : std_logic;
signal \N__19071\ : std_logic;
signal \N__19070\ : std_logic;
signal \N__19067\ : std_logic;
signal \N__19066\ : std_logic;
signal \N__19063\ : std_logic;
signal \N__19062\ : std_logic;
signal \N__19059\ : std_logic;
signal \N__19056\ : std_logic;
signal \N__19053\ : std_logic;
signal \N__19052\ : std_logic;
signal \N__19049\ : std_logic;
signal \N__19048\ : std_logic;
signal \N__19045\ : std_logic;
signal \N__19042\ : std_logic;
signal \N__19039\ : std_logic;
signal \N__19036\ : std_logic;
signal \N__19033\ : std_logic;
signal \N__19026\ : std_logic;
signal \N__19023\ : std_logic;
signal \N__19020\ : std_logic;
signal \N__19017\ : std_logic;
signal \N__18998\ : std_logic;
signal \N__18997\ : std_logic;
signal \N__18994\ : std_logic;
signal \N__18991\ : std_logic;
signal \N__18990\ : std_logic;
signal \N__18987\ : std_logic;
signal \N__18986\ : std_logic;
signal \N__18985\ : std_logic;
signal \N__18984\ : std_logic;
signal \N__18983\ : std_logic;
signal \N__18982\ : std_logic;
signal \N__18981\ : std_logic;
signal \N__18978\ : std_logic;
signal \N__18975\ : std_logic;
signal \N__18972\ : std_logic;
signal \N__18969\ : std_logic;
signal \N__18962\ : std_logic;
signal \N__18957\ : std_logic;
signal \N__18952\ : std_logic;
signal \N__18941\ : std_logic;
signal \N__18940\ : std_logic;
signal \N__18939\ : std_logic;
signal \N__18938\ : std_logic;
signal \N__18937\ : std_logic;
signal \N__18934\ : std_logic;
signal \N__18933\ : std_logic;
signal \N__18932\ : std_logic;
signal \N__18931\ : std_logic;
signal \N__18928\ : std_logic;
signal \N__18927\ : std_logic;
signal \N__18924\ : std_logic;
signal \N__18923\ : std_logic;
signal \N__18922\ : std_logic;
signal \N__18919\ : std_logic;
signal \N__18918\ : std_logic;
signal \N__18917\ : std_logic;
signal \N__18916\ : std_logic;
signal \N__18915\ : std_logic;
signal \N__18914\ : std_logic;
signal \N__18911\ : std_logic;
signal \N__18908\ : std_logic;
signal \N__18905\ : std_logic;
signal \N__18900\ : std_logic;
signal \N__18897\ : std_logic;
signal \N__18892\ : std_logic;
signal \N__18887\ : std_logic;
signal \N__18884\ : std_logic;
signal \N__18881\ : std_logic;
signal \N__18876\ : std_logic;
signal \N__18873\ : std_logic;
signal \N__18870\ : std_logic;
signal \N__18867\ : std_logic;
signal \N__18864\ : std_logic;
signal \N__18863\ : std_logic;
signal \N__18860\ : std_logic;
signal \N__18857\ : std_logic;
signal \N__18854\ : std_logic;
signal \N__18849\ : std_logic;
signal \N__18842\ : std_logic;
signal \N__18841\ : std_logic;
signal \N__18836\ : std_logic;
signal \N__18831\ : std_logic;
signal \N__18828\ : std_logic;
signal \N__18825\ : std_logic;
signal \N__18822\ : std_logic;
signal \N__18817\ : std_logic;
signal \N__18814\ : std_logic;
signal \N__18811\ : std_logic;
signal \N__18808\ : std_logic;
signal \N__18803\ : std_logic;
signal \N__18800\ : std_logic;
signal \N__18787\ : std_logic;
signal \N__18782\ : std_logic;
signal \N__18779\ : std_logic;
signal \N__18776\ : std_logic;
signal \N__18775\ : std_logic;
signal \N__18774\ : std_logic;
signal \N__18773\ : std_logic;
signal \N__18772\ : std_logic;
signal \N__18771\ : std_logic;
signal \N__18770\ : std_logic;
signal \N__18769\ : std_logic;
signal \N__18768\ : std_logic;
signal \N__18767\ : std_logic;
signal \N__18766\ : std_logic;
signal \N__18765\ : std_logic;
signal \N__18764\ : std_logic;
signal \N__18763\ : std_logic;
signal \N__18762\ : std_logic;
signal \N__18759\ : std_logic;
signal \N__18756\ : std_logic;
signal \N__18753\ : std_logic;
signal \N__18750\ : std_logic;
signal \N__18749\ : std_logic;
signal \N__18746\ : std_logic;
signal \N__18745\ : std_logic;
signal \N__18742\ : std_logic;
signal \N__18735\ : std_logic;
signal \N__18730\ : std_logic;
signal \N__18727\ : std_logic;
signal \N__18724\ : std_logic;
signal \N__18719\ : std_logic;
signal \N__18716\ : std_logic;
signal \N__18713\ : std_logic;
signal \N__18710\ : std_logic;
signal \N__18709\ : std_logic;
signal \N__18708\ : std_logic;
signal \N__18707\ : std_logic;
signal \N__18704\ : std_logic;
signal \N__18703\ : std_logic;
signal \N__18700\ : std_logic;
signal \N__18699\ : std_logic;
signal \N__18696\ : std_logic;
signal \N__18693\ : std_logic;
signal \N__18686\ : std_logic;
signal \N__18683\ : std_logic;
signal \N__18678\ : std_logic;
signal \N__18675\ : std_logic;
signal \N__18670\ : std_logic;
signal \N__18667\ : std_logic;
signal \N__18662\ : std_logic;
signal \N__18659\ : std_logic;
signal \N__18656\ : std_logic;
signal \N__18653\ : std_logic;
signal \N__18650\ : std_logic;
signal \N__18639\ : std_logic;
signal \N__18620\ : std_logic;
signal \N__18617\ : std_logic;
signal \N__18614\ : std_logic;
signal \N__18613\ : std_logic;
signal \N__18610\ : std_logic;
signal \N__18607\ : std_logic;
signal \N__18606\ : std_logic;
signal \N__18605\ : std_logic;
signal \N__18604\ : std_logic;
signal \N__18603\ : std_logic;
signal \N__18602\ : std_logic;
signal \N__18601\ : std_logic;
signal \N__18596\ : std_logic;
signal \N__18593\ : std_logic;
signal \N__18590\ : std_logic;
signal \N__18587\ : std_logic;
signal \N__18584\ : std_logic;
signal \N__18581\ : std_logic;
signal \N__18578\ : std_logic;
signal \N__18575\ : std_logic;
signal \N__18568\ : std_logic;
signal \N__18561\ : std_logic;
signal \N__18558\ : std_logic;
signal \N__18553\ : std_logic;
signal \N__18552\ : std_logic;
signal \N__18547\ : std_logic;
signal \N__18544\ : std_logic;
signal \N__18539\ : std_logic;
signal \N__18536\ : std_logic;
signal \N__18533\ : std_logic;
signal \N__18530\ : std_logic;
signal \N__18529\ : std_logic;
signal \N__18528\ : std_logic;
signal \N__18527\ : std_logic;
signal \N__18520\ : std_logic;
signal \N__18517\ : std_logic;
signal \N__18512\ : std_logic;
signal \N__18509\ : std_logic;
signal \N__18506\ : std_logic;
signal \N__18503\ : std_logic;
signal \N__18500\ : std_logic;
signal \N__18497\ : std_logic;
signal \N__18494\ : std_logic;
signal \N__18491\ : std_logic;
signal \N__18488\ : std_logic;
signal \N__18485\ : std_logic;
signal \N__18482\ : std_logic;
signal \N__18479\ : std_logic;
signal \N__18476\ : std_logic;
signal \N__18473\ : std_logic;
signal \N__18470\ : std_logic;
signal \N__18467\ : std_logic;
signal \N__18464\ : std_logic;
signal \N__18461\ : std_logic;
signal \N__18458\ : std_logic;
signal \N__18455\ : std_logic;
signal \N__18452\ : std_logic;
signal \N__18449\ : std_logic;
signal \N__18448\ : std_logic;
signal \N__18445\ : std_logic;
signal \N__18442\ : std_logic;
signal \N__18437\ : std_logic;
signal \N__18434\ : std_logic;
signal \N__18431\ : std_logic;
signal \N__18428\ : std_logic;
signal \N__18425\ : std_logic;
signal \N__18422\ : std_logic;
signal \N__18419\ : std_logic;
signal \N__18416\ : std_logic;
signal \N__18413\ : std_logic;
signal \N__18410\ : std_logic;
signal \N__18407\ : std_logic;
signal \N__18404\ : std_logic;
signal \N__18401\ : std_logic;
signal \N__18398\ : std_logic;
signal \N__18395\ : std_logic;
signal \N__18394\ : std_logic;
signal \N__18393\ : std_logic;
signal \N__18392\ : std_logic;
signal \N__18391\ : std_logic;
signal \N__18390\ : std_logic;
signal \N__18389\ : std_logic;
signal \N__18386\ : std_logic;
signal \N__18383\ : std_logic;
signal \N__18382\ : std_logic;
signal \N__18381\ : std_logic;
signal \N__18378\ : std_logic;
signal \N__18375\ : std_logic;
signal \N__18372\ : std_logic;
signal \N__18367\ : std_logic;
signal \N__18364\ : std_logic;
signal \N__18361\ : std_logic;
signal \N__18356\ : std_logic;
signal \N__18353\ : std_logic;
signal \N__18338\ : std_logic;
signal \N__18337\ : std_logic;
signal \N__18336\ : std_logic;
signal \N__18333\ : std_logic;
signal \N__18332\ : std_logic;
signal \N__18331\ : std_logic;
signal \N__18330\ : std_logic;
signal \N__18327\ : std_logic;
signal \N__18324\ : std_logic;
signal \N__18321\ : std_logic;
signal \N__18316\ : std_logic;
signal \N__18313\ : std_logic;
signal \N__18302\ : std_logic;
signal \N__18299\ : std_logic;
signal \N__18296\ : std_logic;
signal \N__18293\ : std_logic;
signal \N__18290\ : std_logic;
signal \N__18287\ : std_logic;
signal \N__18284\ : std_logic;
signal \N__18281\ : std_logic;
signal \N__18278\ : std_logic;
signal \N__18275\ : std_logic;
signal \N__18272\ : std_logic;
signal \N__18269\ : std_logic;
signal \N__18266\ : std_logic;
signal \N__18263\ : std_logic;
signal \N__18260\ : std_logic;
signal \N__18259\ : std_logic;
signal \N__18256\ : std_logic;
signal \N__18255\ : std_logic;
signal \N__18252\ : std_logic;
signal \N__18251\ : std_logic;
signal \N__18248\ : std_logic;
signal \N__18245\ : std_logic;
signal \N__18240\ : std_logic;
signal \N__18239\ : std_logic;
signal \N__18236\ : std_logic;
signal \N__18231\ : std_logic;
signal \N__18228\ : std_logic;
signal \N__18227\ : std_logic;
signal \N__18226\ : std_logic;
signal \N__18225\ : std_logic;
signal \N__18224\ : std_logic;
signal \N__18221\ : std_logic;
signal \N__18218\ : std_logic;
signal \N__18215\ : std_logic;
signal \N__18210\ : std_logic;
signal \N__18205\ : std_logic;
signal \N__18194\ : std_logic;
signal \N__18193\ : std_logic;
signal \N__18192\ : std_logic;
signal \N__18191\ : std_logic;
signal \N__18188\ : std_logic;
signal \N__18187\ : std_logic;
signal \N__18186\ : std_logic;
signal \N__18185\ : std_logic;
signal \N__18184\ : std_logic;
signal \N__18179\ : std_logic;
signal \N__18176\ : std_logic;
signal \N__18169\ : std_logic;
signal \N__18166\ : std_logic;
signal \N__18165\ : std_logic;
signal \N__18164\ : std_logic;
signal \N__18163\ : std_logic;
signal \N__18160\ : std_logic;
signal \N__18153\ : std_logic;
signal \N__18150\ : std_logic;
signal \N__18147\ : std_logic;
signal \N__18142\ : std_logic;
signal \N__18139\ : std_logic;
signal \N__18136\ : std_logic;
signal \N__18125\ : std_logic;
signal \N__18124\ : std_logic;
signal \N__18123\ : std_logic;
signal \N__18120\ : std_logic;
signal \N__18119\ : std_logic;
signal \N__18114\ : std_logic;
signal \N__18111\ : std_logic;
signal \N__18108\ : std_logic;
signal \N__18105\ : std_logic;
signal \N__18104\ : std_logic;
signal \N__18103\ : std_logic;
signal \N__18102\ : std_logic;
signal \N__18099\ : std_logic;
signal \N__18094\ : std_logic;
signal \N__18091\ : std_logic;
signal \N__18090\ : std_logic;
signal \N__18089\ : std_logic;
signal \N__18088\ : std_logic;
signal \N__18083\ : std_logic;
signal \N__18080\ : std_logic;
signal \N__18075\ : std_logic;
signal \N__18070\ : std_logic;
signal \N__18067\ : std_logic;
signal \N__18056\ : std_logic;
signal \N__18053\ : std_logic;
signal \N__18050\ : std_logic;
signal \N__18047\ : std_logic;
signal \N__18044\ : std_logic;
signal \N__18041\ : std_logic;
signal \N__18038\ : std_logic;
signal \N__18035\ : std_logic;
signal \N__18032\ : std_logic;
signal \N__18029\ : std_logic;
signal \N__18028\ : std_logic;
signal \N__18027\ : std_logic;
signal \N__18026\ : std_logic;
signal \N__18023\ : std_logic;
signal \N__18020\ : std_logic;
signal \N__18019\ : std_logic;
signal \N__18018\ : std_logic;
signal \N__18013\ : std_logic;
signal \N__18008\ : std_logic;
signal \N__18007\ : std_logic;
signal \N__18006\ : std_logic;
signal \N__18005\ : std_logic;
signal \N__18004\ : std_logic;
signal \N__18003\ : std_logic;
signal \N__18002\ : std_logic;
signal \N__17999\ : std_logic;
signal \N__17996\ : std_logic;
signal \N__17991\ : std_logic;
signal \N__17984\ : std_logic;
signal \N__17975\ : std_logic;
signal \N__17974\ : std_logic;
signal \N__17973\ : std_logic;
signal \N__17970\ : std_logic;
signal \N__17963\ : std_logic;
signal \N__17962\ : std_logic;
signal \N__17959\ : std_logic;
signal \N__17958\ : std_logic;
signal \N__17955\ : std_logic;
signal \N__17952\ : std_logic;
signal \N__17949\ : std_logic;
signal \N__17946\ : std_logic;
signal \N__17939\ : std_logic;
signal \N__17930\ : std_logic;
signal \N__17927\ : std_logic;
signal \N__17924\ : std_logic;
signal \N__17921\ : std_logic;
signal \N__17918\ : std_logic;
signal \N__17915\ : std_logic;
signal \N__17912\ : std_logic;
signal \N__17909\ : std_logic;
signal \N__17906\ : std_logic;
signal \N__17903\ : std_logic;
signal \N__17900\ : std_logic;
signal \N__17897\ : std_logic;
signal \N__17894\ : std_logic;
signal \N__17891\ : std_logic;
signal \N__17888\ : std_logic;
signal \N__17885\ : std_logic;
signal \N__17882\ : std_logic;
signal \N__17879\ : std_logic;
signal \N__17876\ : std_logic;
signal \N__17875\ : std_logic;
signal \N__17874\ : std_logic;
signal \N__17873\ : std_logic;
signal \N__17872\ : std_logic;
signal \N__17871\ : std_logic;
signal \N__17870\ : std_logic;
signal \N__17869\ : std_logic;
signal \N__17868\ : std_logic;
signal \N__17865\ : std_logic;
signal \N__17858\ : std_logic;
signal \N__17853\ : std_logic;
signal \N__17848\ : std_logic;
signal \N__17845\ : std_logic;
signal \N__17834\ : std_logic;
signal \N__17831\ : std_logic;
signal \N__17828\ : std_logic;
signal \N__17825\ : std_logic;
signal \N__17824\ : std_logic;
signal \N__17823\ : std_logic;
signal \N__17820\ : std_logic;
signal \N__17815\ : std_logic;
signal \N__17810\ : std_logic;
signal \N__17807\ : std_logic;
signal \N__17804\ : std_logic;
signal \N__17801\ : std_logic;
signal \N__17798\ : std_logic;
signal \N__17795\ : std_logic;
signal \N__17794\ : std_logic;
signal \N__17793\ : std_logic;
signal \N__17792\ : std_logic;
signal \N__17791\ : std_logic;
signal \N__17790\ : std_logic;
signal \N__17787\ : std_logic;
signal \N__17786\ : std_logic;
signal \N__17783\ : std_logic;
signal \N__17782\ : std_logic;
signal \N__17781\ : std_logic;
signal \N__17780\ : std_logic;
signal \N__17777\ : std_logic;
signal \N__17774\ : std_logic;
signal \N__17773\ : std_logic;
signal \N__17770\ : std_logic;
signal \N__17769\ : std_logic;
signal \N__17768\ : std_logic;
signal \N__17765\ : std_logic;
signal \N__17764\ : std_logic;
signal \N__17761\ : std_logic;
signal \N__17756\ : std_logic;
signal \N__17753\ : std_logic;
signal \N__17742\ : std_logic;
signal \N__17737\ : std_logic;
signal \N__17730\ : std_logic;
signal \N__17717\ : std_logic;
signal \N__17716\ : std_logic;
signal \N__17715\ : std_logic;
signal \N__17714\ : std_logic;
signal \N__17707\ : std_logic;
signal \N__17704\ : std_logic;
signal \N__17703\ : std_logic;
signal \N__17702\ : std_logic;
signal \N__17701\ : std_logic;
signal \N__17700\ : std_logic;
signal \N__17699\ : std_logic;
signal \N__17698\ : std_logic;
signal \N__17693\ : std_logic;
signal \N__17692\ : std_logic;
signal \N__17687\ : std_logic;
signal \N__17684\ : std_logic;
signal \N__17683\ : std_logic;
signal \N__17680\ : std_logic;
signal \N__17679\ : std_logic;
signal \N__17676\ : std_logic;
signal \N__17673\ : std_logic;
signal \N__17670\ : std_logic;
signal \N__17669\ : std_logic;
signal \N__17668\ : std_logic;
signal \N__17667\ : std_logic;
signal \N__17666\ : std_logic;
signal \N__17663\ : std_logic;
signal \N__17660\ : std_logic;
signal \N__17657\ : std_logic;
signal \N__17654\ : std_logic;
signal \N__17651\ : std_logic;
signal \N__17648\ : std_logic;
signal \N__17645\ : std_logic;
signal \N__17640\ : std_logic;
signal \N__17639\ : std_logic;
signal \N__17636\ : std_logic;
signal \N__17633\ : std_logic;
signal \N__17628\ : std_logic;
signal \N__17625\ : std_logic;
signal \N__17622\ : std_logic;
signal \N__17613\ : std_logic;
signal \N__17608\ : std_logic;
signal \N__17605\ : std_logic;
signal \N__17588\ : std_logic;
signal \N__17585\ : std_logic;
signal \N__17582\ : std_logic;
signal \N__17579\ : std_logic;
signal \N__17576\ : std_logic;
signal \N__17573\ : std_logic;
signal \N__17572\ : std_logic;
signal \N__17569\ : std_logic;
signal \N__17566\ : std_logic;
signal \N__17563\ : std_logic;
signal \N__17560\ : std_logic;
signal \N__17557\ : std_logic;
signal \N__17552\ : std_logic;
signal \N__17549\ : std_logic;
signal \N__17546\ : std_logic;
signal \N__17543\ : std_logic;
signal \N__17540\ : std_logic;
signal \N__17537\ : std_logic;
signal \N__17536\ : std_logic;
signal \N__17535\ : std_logic;
signal \N__17534\ : std_logic;
signal \N__17527\ : std_logic;
signal \N__17526\ : std_logic;
signal \N__17525\ : std_logic;
signal \N__17522\ : std_logic;
signal \N__17519\ : std_logic;
signal \N__17514\ : std_logic;
signal \N__17507\ : std_logic;
signal \N__17506\ : std_logic;
signal \N__17503\ : std_logic;
signal \N__17500\ : std_logic;
signal \N__17495\ : std_logic;
signal \N__17492\ : std_logic;
signal \N__17489\ : std_logic;
signal \N__17486\ : std_logic;
signal \N__17483\ : std_logic;
signal \N__17482\ : std_logic;
signal \N__17479\ : std_logic;
signal \N__17476\ : std_logic;
signal \N__17471\ : std_logic;
signal \N__17468\ : std_logic;
signal \N__17467\ : std_logic;
signal \N__17464\ : std_logic;
signal \N__17461\ : std_logic;
signal \N__17458\ : std_logic;
signal \N__17455\ : std_logic;
signal \N__17452\ : std_logic;
signal \N__17449\ : std_logic;
signal \N__17444\ : std_logic;
signal \N__17441\ : std_logic;
signal \N__17438\ : std_logic;
signal \N__17435\ : std_logic;
signal \N__17432\ : std_logic;
signal \N__17429\ : std_logic;
signal \N__17426\ : std_logic;
signal \N__17423\ : std_logic;
signal \N__17420\ : std_logic;
signal \N__17417\ : std_logic;
signal \N__17414\ : std_logic;
signal \N__17411\ : std_logic;
signal \N__17410\ : std_logic;
signal \N__17409\ : std_logic;
signal \N__17404\ : std_logic;
signal \N__17401\ : std_logic;
signal \N__17400\ : std_logic;
signal \N__17399\ : std_logic;
signal \N__17398\ : std_logic;
signal \N__17395\ : std_logic;
signal \N__17392\ : std_logic;
signal \N__17391\ : std_logic;
signal \N__17390\ : std_logic;
signal \N__17387\ : std_logic;
signal \N__17384\ : std_logic;
signal \N__17381\ : std_logic;
signal \N__17380\ : std_logic;
signal \N__17377\ : std_logic;
signal \N__17374\ : std_logic;
signal \N__17371\ : std_logic;
signal \N__17368\ : std_logic;
signal \N__17363\ : std_logic;
signal \N__17360\ : std_logic;
signal \N__17357\ : std_logic;
signal \N__17342\ : std_logic;
signal \N__17341\ : std_logic;
signal \N__17338\ : std_logic;
signal \N__17335\ : std_logic;
signal \N__17332\ : std_logic;
signal \N__17327\ : std_logic;
signal \N__17324\ : std_logic;
signal \N__17321\ : std_logic;
signal \N__17318\ : std_logic;
signal \N__17315\ : std_logic;
signal \N__17312\ : std_logic;
signal \N__17309\ : std_logic;
signal \N__17306\ : std_logic;
signal \N__17303\ : std_logic;
signal \N__17300\ : std_logic;
signal \N__17297\ : std_logic;
signal \N__17294\ : std_logic;
signal \N__17291\ : std_logic;
signal \N__17288\ : std_logic;
signal \N__17285\ : std_logic;
signal \N__17282\ : std_logic;
signal \N__17279\ : std_logic;
signal \N__17276\ : std_logic;
signal \N__17273\ : std_logic;
signal \N__17270\ : std_logic;
signal \N__17267\ : std_logic;
signal \N__17264\ : std_logic;
signal \N__17261\ : std_logic;
signal \N__17258\ : std_logic;
signal \N__17255\ : std_logic;
signal \N__17252\ : std_logic;
signal \N__17249\ : std_logic;
signal \N__17246\ : std_logic;
signal \N__17243\ : std_logic;
signal \N__17240\ : std_logic;
signal \N__17237\ : std_logic;
signal \N__17234\ : std_logic;
signal \N__17231\ : std_logic;
signal \N__17228\ : std_logic;
signal \N__17225\ : std_logic;
signal \N__17222\ : std_logic;
signal \N__17219\ : std_logic;
signal \N__17216\ : std_logic;
signal \N__17213\ : std_logic;
signal \N__17210\ : std_logic;
signal \N__17207\ : std_logic;
signal \N__17204\ : std_logic;
signal \N__17201\ : std_logic;
signal \N__17198\ : std_logic;
signal \N__17195\ : std_logic;
signal \N__17192\ : std_logic;
signal \N__17189\ : std_logic;
signal \N__17186\ : std_logic;
signal \N__17183\ : std_logic;
signal \N__17180\ : std_logic;
signal \N__17177\ : std_logic;
signal \N__17176\ : std_logic;
signal \N__17175\ : std_logic;
signal \N__17174\ : std_logic;
signal \N__17173\ : std_logic;
signal \N__17172\ : std_logic;
signal \N__17171\ : std_logic;
signal \N__17170\ : std_logic;
signal \N__17167\ : std_logic;
signal \N__17154\ : std_logic;
signal \N__17151\ : std_logic;
signal \N__17148\ : std_logic;
signal \N__17145\ : std_logic;
signal \N__17142\ : std_logic;
signal \N__17139\ : std_logic;
signal \N__17136\ : std_logic;
signal \N__17133\ : std_logic;
signal \N__17126\ : std_logic;
signal \N__17123\ : std_logic;
signal \N__17120\ : std_logic;
signal \N__17117\ : std_logic;
signal \N__17116\ : std_logic;
signal \N__17115\ : std_logic;
signal \N__17114\ : std_logic;
signal \N__17113\ : std_logic;
signal \N__17112\ : std_logic;
signal \N__17109\ : std_logic;
signal \N__17108\ : std_logic;
signal \N__17105\ : std_logic;
signal \N__17102\ : std_logic;
signal \N__17099\ : std_logic;
signal \N__17094\ : std_logic;
signal \N__17089\ : std_logic;
signal \N__17088\ : std_logic;
signal \N__17087\ : std_logic;
signal \N__17084\ : std_logic;
signal \N__17081\ : std_logic;
signal \N__17074\ : std_logic;
signal \N__17069\ : std_logic;
signal \N__17060\ : std_logic;
signal \N__17057\ : std_logic;
signal \N__17054\ : std_logic;
signal \N__17051\ : std_logic;
signal \N__17048\ : std_logic;
signal \N__17045\ : std_logic;
signal \N__17042\ : std_logic;
signal \N__17039\ : std_logic;
signal \N__17036\ : std_logic;
signal \N__17033\ : std_logic;
signal \N__17032\ : std_logic;
signal \N__17031\ : std_logic;
signal \N__17030\ : std_logic;
signal \N__17021\ : std_logic;
signal \N__17020\ : std_logic;
signal \N__17019\ : std_logic;
signal \N__17018\ : std_logic;
signal \N__17017\ : std_logic;
signal \N__17014\ : std_logic;
signal \N__17013\ : std_logic;
signal \N__17012\ : std_logic;
signal \N__17011\ : std_logic;
signal \N__17004\ : std_logic;
signal \N__17001\ : std_logic;
signal \N__17000\ : std_logic;
signal \N__16997\ : std_logic;
signal \N__16994\ : std_logic;
signal \N__16991\ : std_logic;
signal \N__16988\ : std_logic;
signal \N__16985\ : std_logic;
signal \N__16982\ : std_logic;
signal \N__16979\ : std_logic;
signal \N__16976\ : std_logic;
signal \N__16969\ : std_logic;
signal \N__16958\ : std_logic;
signal \N__16957\ : std_logic;
signal \N__16954\ : std_logic;
signal \N__16953\ : std_logic;
signal \N__16952\ : std_logic;
signal \N__16951\ : std_logic;
signal \N__16950\ : std_logic;
signal \N__16947\ : std_logic;
signal \N__16946\ : std_logic;
signal \N__16943\ : std_logic;
signal \N__16940\ : std_logic;
signal \N__16937\ : std_logic;
signal \N__16936\ : std_logic;
signal \N__16935\ : std_logic;
signal \N__16930\ : std_logic;
signal \N__16927\ : std_logic;
signal \N__16924\ : std_logic;
signal \N__16921\ : std_logic;
signal \N__16916\ : std_logic;
signal \N__16911\ : std_logic;
signal \N__16906\ : std_logic;
signal \N__16895\ : std_logic;
signal \N__16892\ : std_logic;
signal \N__16889\ : std_logic;
signal \N__16886\ : std_logic;
signal \N__16883\ : std_logic;
signal \N__16880\ : std_logic;
signal \N__16877\ : std_logic;
signal \N__16874\ : std_logic;
signal \N__16871\ : std_logic;
signal \N__16868\ : std_logic;
signal \N__16865\ : std_logic;
signal \N__16862\ : std_logic;
signal \N__16859\ : std_logic;
signal \N__16856\ : std_logic;
signal \N__16855\ : std_logic;
signal \N__16852\ : std_logic;
signal \N__16849\ : std_logic;
signal \N__16844\ : std_logic;
signal \N__16841\ : std_logic;
signal \N__16838\ : std_logic;
signal \N__16835\ : std_logic;
signal \N__16832\ : std_logic;
signal \N__16829\ : std_logic;
signal \N__16826\ : std_logic;
signal \N__16823\ : std_logic;
signal \N__16820\ : std_logic;
signal \N__16817\ : std_logic;
signal \N__16814\ : std_logic;
signal \N__16811\ : std_logic;
signal \N__16808\ : std_logic;
signal \N__16805\ : std_logic;
signal \N__16804\ : std_logic;
signal \N__16803\ : std_logic;
signal \N__16800\ : std_logic;
signal \N__16797\ : std_logic;
signal \N__16794\ : std_logic;
signal \N__16787\ : std_logic;
signal \N__16784\ : std_logic;
signal \N__16781\ : std_logic;
signal \N__16778\ : std_logic;
signal \N__16775\ : std_logic;
signal \N__16772\ : std_logic;
signal \N__16769\ : std_logic;
signal \N__16766\ : std_logic;
signal \N__16763\ : std_logic;
signal \N__16760\ : std_logic;
signal \N__16757\ : std_logic;
signal \N__16754\ : std_logic;
signal \N__16751\ : std_logic;
signal \N__16748\ : std_logic;
signal \N__16745\ : std_logic;
signal \N__16742\ : std_logic;
signal \N__16739\ : std_logic;
signal \N__16736\ : std_logic;
signal \N__16733\ : std_logic;
signal \N__16732\ : std_logic;
signal \N__16729\ : std_logic;
signal \N__16726\ : std_logic;
signal \N__16725\ : std_logic;
signal \N__16724\ : std_logic;
signal \N__16723\ : std_logic;
signal \N__16722\ : std_logic;
signal \N__16719\ : std_logic;
signal \N__16716\ : std_logic;
signal \N__16713\ : std_logic;
signal \N__16706\ : std_logic;
signal \N__16697\ : std_logic;
signal \N__16694\ : std_logic;
signal \N__16691\ : std_logic;
signal \N__16688\ : std_logic;
signal \N__16685\ : std_logic;
signal \N__16682\ : std_logic;
signal \N__16679\ : std_logic;
signal \N__16678\ : std_logic;
signal \N__16677\ : std_logic;
signal \N__16674\ : std_logic;
signal \N__16673\ : std_logic;
signal \N__16670\ : std_logic;
signal \N__16667\ : std_logic;
signal \N__16664\ : std_logic;
signal \N__16661\ : std_logic;
signal \N__16656\ : std_logic;
signal \N__16651\ : std_logic;
signal \N__16648\ : std_logic;
signal \N__16645\ : std_logic;
signal \N__16642\ : std_logic;
signal \N__16639\ : std_logic;
signal \N__16634\ : std_logic;
signal \N__16633\ : std_logic;
signal \N__16628\ : std_logic;
signal \N__16625\ : std_logic;
signal \N__16622\ : std_logic;
signal \N__16619\ : std_logic;
signal \N__16616\ : std_logic;
signal \N__16613\ : std_logic;
signal \N__16610\ : std_logic;
signal \N__16607\ : std_logic;
signal \N__16604\ : std_logic;
signal \N__16601\ : std_logic;
signal \N__16598\ : std_logic;
signal \N__16595\ : std_logic;
signal \N__16592\ : std_logic;
signal \N__16589\ : std_logic;
signal \N__16586\ : std_logic;
signal \N__16583\ : std_logic;
signal \N__16580\ : std_logic;
signal \N__16577\ : std_logic;
signal \N__16574\ : std_logic;
signal \N__16571\ : std_logic;
signal \N__16568\ : std_logic;
signal \N__16565\ : std_logic;
signal \N__16562\ : std_logic;
signal \N__16559\ : std_logic;
signal \N__16556\ : std_logic;
signal \N__16553\ : std_logic;
signal \N__16550\ : std_logic;
signal \N__16547\ : std_logic;
signal \N__16544\ : std_logic;
signal \N__16541\ : std_logic;
signal \N__16538\ : std_logic;
signal \N__16535\ : std_logic;
signal \N__16532\ : std_logic;
signal \N__16529\ : std_logic;
signal \N__16526\ : std_logic;
signal \N__16523\ : std_logic;
signal \N__16520\ : std_logic;
signal \N__16517\ : std_logic;
signal \N__16514\ : std_logic;
signal \N__16511\ : std_logic;
signal \N__16508\ : std_logic;
signal \N__16505\ : std_logic;
signal \N__16502\ : std_logic;
signal \N__16499\ : std_logic;
signal \N__16496\ : std_logic;
signal \N__16493\ : std_logic;
signal \N__16490\ : std_logic;
signal \N__16487\ : std_logic;
signal \N__16484\ : std_logic;
signal \N__16481\ : std_logic;
signal \N__16480\ : std_logic;
signal \N__16479\ : std_logic;
signal \N__16478\ : std_logic;
signal \N__16475\ : std_logic;
signal \N__16474\ : std_logic;
signal \N__16473\ : std_logic;
signal \N__16470\ : std_logic;
signal \N__16467\ : std_logic;
signal \N__16466\ : std_logic;
signal \N__16465\ : std_logic;
signal \N__16462\ : std_logic;
signal \N__16459\ : std_logic;
signal \N__16458\ : std_logic;
signal \N__16455\ : std_logic;
signal \N__16452\ : std_logic;
signal \N__16445\ : std_logic;
signal \N__16442\ : std_logic;
signal \N__16437\ : std_logic;
signal \N__16434\ : std_logic;
signal \N__16431\ : std_logic;
signal \N__16418\ : std_logic;
signal \N__16415\ : std_logic;
signal \N__16412\ : std_logic;
signal \N__16409\ : std_logic;
signal \N__16406\ : std_logic;
signal \N__16405\ : std_logic;
signal \N__16402\ : std_logic;
signal \N__16401\ : std_logic;
signal \N__16400\ : std_logic;
signal \N__16397\ : std_logic;
signal \N__16396\ : std_logic;
signal \N__16395\ : std_logic;
signal \N__16394\ : std_logic;
signal \N__16391\ : std_logic;
signal \N__16388\ : std_logic;
signal \N__16381\ : std_logic;
signal \N__16378\ : std_logic;
signal \N__16375\ : std_logic;
signal \N__16374\ : std_logic;
signal \N__16371\ : std_logic;
signal \N__16368\ : std_logic;
signal \N__16361\ : std_logic;
signal \N__16358\ : std_logic;
signal \N__16349\ : std_logic;
signal \N__16346\ : std_logic;
signal \N__16343\ : std_logic;
signal \N__16340\ : std_logic;
signal \N__16337\ : std_logic;
signal \N__16334\ : std_logic;
signal \N__16331\ : std_logic;
signal \N__16330\ : std_logic;
signal \N__16327\ : std_logic;
signal \N__16324\ : std_logic;
signal \N__16321\ : std_logic;
signal \N__16318\ : std_logic;
signal \N__16315\ : std_logic;
signal \N__16312\ : std_logic;
signal \N__16309\ : std_logic;
signal \N__16304\ : std_logic;
signal \N__16301\ : std_logic;
signal \N__16298\ : std_logic;
signal \N__16295\ : std_logic;
signal \N__16292\ : std_logic;
signal \N__16289\ : std_logic;
signal \N__16286\ : std_logic;
signal \N__16283\ : std_logic;
signal \N__16280\ : std_logic;
signal \N__16277\ : std_logic;
signal \N__16274\ : std_logic;
signal \N__16271\ : std_logic;
signal \N__16270\ : std_logic;
signal \N__16267\ : std_logic;
signal \N__16264\ : std_logic;
signal \N__16259\ : std_logic;
signal \N__16256\ : std_logic;
signal \N__16253\ : std_logic;
signal \N__16250\ : std_logic;
signal \N__16247\ : std_logic;
signal \N__16244\ : std_logic;
signal \N__16241\ : std_logic;
signal \N__16238\ : std_logic;
signal \N__16235\ : std_logic;
signal \N__16232\ : std_logic;
signal \N__16229\ : std_logic;
signal \N__16228\ : std_logic;
signal \N__16225\ : std_logic;
signal \N__16224\ : std_logic;
signal \N__16223\ : std_logic;
signal \N__16222\ : std_logic;
signal \N__16221\ : std_logic;
signal \N__16218\ : std_logic;
signal \N__16217\ : std_logic;
signal \N__16214\ : std_logic;
signal \N__16211\ : std_logic;
signal \N__16206\ : std_logic;
signal \N__16203\ : std_logic;
signal \N__16202\ : std_logic;
signal \N__16199\ : std_logic;
signal \N__16196\ : std_logic;
signal \N__16187\ : std_logic;
signal \N__16184\ : std_logic;
signal \N__16175\ : std_logic;
signal \N__16174\ : std_logic;
signal \N__16173\ : std_logic;
signal \N__16172\ : std_logic;
signal \N__16171\ : std_logic;
signal \N__16170\ : std_logic;
signal \N__16169\ : std_logic;
signal \N__16168\ : std_logic;
signal \N__16165\ : std_logic;
signal \N__16162\ : std_logic;
signal \N__16159\ : std_logic;
signal \N__16152\ : std_logic;
signal \N__16151\ : std_logic;
signal \N__16150\ : std_logic;
signal \N__16147\ : std_logic;
signal \N__16144\ : std_logic;
signal \N__16141\ : std_logic;
signal \N__16138\ : std_logic;
signal \N__16133\ : std_logic;
signal \N__16128\ : std_logic;
signal \N__16115\ : std_logic;
signal \N__16114\ : std_logic;
signal \N__16113\ : std_logic;
signal \N__16112\ : std_logic;
signal \N__16111\ : std_logic;
signal \N__16108\ : std_logic;
signal \N__16105\ : std_logic;
signal \N__16102\ : std_logic;
signal \N__16101\ : std_logic;
signal \N__16100\ : std_logic;
signal \N__16097\ : std_logic;
signal \N__16094\ : std_logic;
signal \N__16091\ : std_logic;
signal \N__16088\ : std_logic;
signal \N__16085\ : std_logic;
signal \N__16078\ : std_logic;
signal \N__16077\ : std_logic;
signal \N__16076\ : std_logic;
signal \N__16069\ : std_logic;
signal \N__16064\ : std_logic;
signal \N__16059\ : std_logic;
signal \N__16056\ : std_logic;
signal \N__16051\ : std_logic;
signal \N__16046\ : std_logic;
signal \N__16045\ : std_logic;
signal \N__16044\ : std_logic;
signal \N__16041\ : std_logic;
signal \N__16038\ : std_logic;
signal \N__16037\ : std_logic;
signal \N__16034\ : std_logic;
signal \N__16031\ : std_logic;
signal \N__16028\ : std_logic;
signal \N__16025\ : std_logic;
signal \N__16024\ : std_logic;
signal \N__16023\ : std_logic;
signal \N__16020\ : std_logic;
signal \N__16017\ : std_logic;
signal \N__16014\ : std_logic;
signal \N__16011\ : std_logic;
signal \N__16008\ : std_logic;
signal \N__16005\ : std_logic;
signal \N__15992\ : std_logic;
signal \N__15989\ : std_logic;
signal \N__15986\ : std_logic;
signal \N__15983\ : std_logic;
signal \N__15980\ : std_logic;
signal \N__15977\ : std_logic;
signal \N__15974\ : std_logic;
signal \N__15971\ : std_logic;
signal \N__15968\ : std_logic;
signal \N__15965\ : std_logic;
signal \N__15962\ : std_logic;
signal \N__15959\ : std_logic;
signal \N__15956\ : std_logic;
signal \N__15953\ : std_logic;
signal \N__15950\ : std_logic;
signal \N__15947\ : std_logic;
signal \N__15946\ : std_logic;
signal \N__15945\ : std_logic;
signal \N__15942\ : std_logic;
signal \N__15937\ : std_logic;
signal \N__15934\ : std_logic;
signal \N__15931\ : std_logic;
signal \N__15926\ : std_logic;
signal \N__15923\ : std_logic;
signal \N__15920\ : std_logic;
signal \N__15917\ : std_logic;
signal \N__15914\ : std_logic;
signal \N__15911\ : std_logic;
signal \N__15910\ : std_logic;
signal \N__15907\ : std_logic;
signal \N__15904\ : std_logic;
signal \N__15903\ : std_logic;
signal \N__15902\ : std_logic;
signal \N__15901\ : std_logic;
signal \N__15896\ : std_logic;
signal \N__15893\ : std_logic;
signal \N__15890\ : std_logic;
signal \N__15887\ : std_logic;
signal \N__15884\ : std_logic;
signal \N__15879\ : std_logic;
signal \N__15872\ : std_logic;
signal \N__15871\ : std_logic;
signal \N__15868\ : std_logic;
signal \N__15867\ : std_logic;
signal \N__15866\ : std_logic;
signal \N__15865\ : std_logic;
signal \N__15862\ : std_logic;
signal \N__15859\ : std_logic;
signal \N__15854\ : std_logic;
signal \N__15851\ : std_logic;
signal \N__15848\ : std_logic;
signal \N__15847\ : std_logic;
signal \N__15846\ : std_logic;
signal \N__15845\ : std_logic;
signal \N__15844\ : std_logic;
signal \N__15841\ : std_logic;
signal \N__15838\ : std_logic;
signal \N__15835\ : std_logic;
signal \N__15832\ : std_logic;
signal \N__15829\ : std_logic;
signal \N__15822\ : std_logic;
signal \N__15809\ : std_logic;
signal \N__15806\ : std_logic;
signal \N__15803\ : std_logic;
signal \N__15800\ : std_logic;
signal \N__15797\ : std_logic;
signal \N__15794\ : std_logic;
signal \N__15791\ : std_logic;
signal \N__15788\ : std_logic;
signal \N__15787\ : std_logic;
signal \N__15782\ : std_logic;
signal \N__15779\ : std_logic;
signal \N__15776\ : std_logic;
signal \N__15775\ : std_logic;
signal \N__15770\ : std_logic;
signal \N__15767\ : std_logic;
signal \N__15764\ : std_logic;
signal \N__15761\ : std_logic;
signal \N__15758\ : std_logic;
signal \N__15755\ : std_logic;
signal \N__15752\ : std_logic;
signal \N__15749\ : std_logic;
signal \N__15746\ : std_logic;
signal \N__15743\ : std_logic;
signal \N__15742\ : std_logic;
signal \N__15739\ : std_logic;
signal \N__15736\ : std_logic;
signal \N__15731\ : std_logic;
signal \N__15728\ : std_logic;
signal \N__15725\ : std_logic;
signal \N__15722\ : std_logic;
signal \N__15721\ : std_logic;
signal \N__15720\ : std_logic;
signal \N__15719\ : std_logic;
signal \N__15716\ : std_logic;
signal \N__15711\ : std_logic;
signal \N__15708\ : std_logic;
signal \N__15705\ : std_logic;
signal \N__15702\ : std_logic;
signal \N__15699\ : std_logic;
signal \N__15696\ : std_logic;
signal \N__15693\ : std_logic;
signal \N__15686\ : std_logic;
signal \N__15685\ : std_logic;
signal \N__15684\ : std_logic;
signal \N__15683\ : std_logic;
signal \N__15682\ : std_logic;
signal \N__15681\ : std_logic;
signal \N__15680\ : std_logic;
signal \N__15679\ : std_logic;
signal \N__15678\ : std_logic;
signal \N__15677\ : std_logic;
signal \N__15674\ : std_logic;
signal \N__15671\ : std_logic;
signal \N__15668\ : std_logic;
signal \N__15665\ : std_logic;
signal \N__15660\ : std_logic;
signal \N__15655\ : std_logic;
signal \N__15652\ : std_logic;
signal \N__15645\ : std_logic;
signal \N__15642\ : std_logic;
signal \N__15639\ : std_logic;
signal \N__15634\ : std_logic;
signal \N__15633\ : std_logic;
signal \N__15632\ : std_logic;
signal \N__15629\ : std_logic;
signal \N__15626\ : std_logic;
signal \N__15621\ : std_logic;
signal \N__15618\ : std_logic;
signal \N__15613\ : std_logic;
signal \N__15608\ : std_logic;
signal \N__15599\ : std_logic;
signal \N__15598\ : std_logic;
signal \N__15597\ : std_logic;
signal \N__15596\ : std_logic;
signal \N__15595\ : std_logic;
signal \N__15594\ : std_logic;
signal \N__15581\ : std_logic;
signal \N__15578\ : std_logic;
signal \N__15577\ : std_logic;
signal \N__15576\ : std_logic;
signal \N__15575\ : std_logic;
signal \N__15572\ : std_logic;
signal \N__15567\ : std_logic;
signal \N__15566\ : std_logic;
signal \N__15565\ : std_logic;
signal \N__15564\ : std_logic;
signal \N__15563\ : std_logic;
signal \N__15560\ : std_logic;
signal \N__15559\ : std_logic;
signal \N__15554\ : std_logic;
signal \N__15541\ : std_logic;
signal \N__15536\ : std_logic;
signal \N__15535\ : std_logic;
signal \N__15534\ : std_logic;
signal \N__15531\ : std_logic;
signal \N__15526\ : std_logic;
signal \N__15521\ : std_logic;
signal \N__15518\ : std_logic;
signal \N__15515\ : std_logic;
signal \N__15512\ : std_logic;
signal \N__15509\ : std_logic;
signal \N__15506\ : std_logic;
signal \N__15503\ : std_logic;
signal \N__15500\ : std_logic;
signal \N__15497\ : std_logic;
signal \N__15494\ : std_logic;
signal \N__15491\ : std_logic;
signal \N__15490\ : std_logic;
signal \N__15487\ : std_logic;
signal \N__15484\ : std_logic;
signal \N__15481\ : std_logic;
signal \N__15478\ : std_logic;
signal \N__15477\ : std_logic;
signal \N__15474\ : std_logic;
signal \N__15471\ : std_logic;
signal \N__15470\ : std_logic;
signal \N__15469\ : std_logic;
signal \N__15466\ : std_logic;
signal \N__15463\ : std_logic;
signal \N__15460\ : std_logic;
signal \N__15457\ : std_logic;
signal \N__15454\ : std_logic;
signal \N__15451\ : std_logic;
signal \N__15440\ : std_logic;
signal \N__15439\ : std_logic;
signal \N__15434\ : std_logic;
signal \N__15431\ : std_logic;
signal \N__15428\ : std_logic;
signal \N__15425\ : std_logic;
signal \N__15422\ : std_logic;
signal \N__15419\ : std_logic;
signal \N__15416\ : std_logic;
signal \N__15413\ : std_logic;
signal \N__15412\ : std_logic;
signal \N__15409\ : std_logic;
signal \N__15406\ : std_logic;
signal \N__15403\ : std_logic;
signal \N__15400\ : std_logic;
signal \N__15395\ : std_logic;
signal \N__15392\ : std_logic;
signal \N__15389\ : std_logic;
signal \N__15386\ : std_logic;
signal \N__15383\ : std_logic;
signal \N__15380\ : std_logic;
signal \N__15377\ : std_logic;
signal \N__15376\ : std_logic;
signal \N__15375\ : std_logic;
signal \N__15374\ : std_logic;
signal \N__15373\ : std_logic;
signal \N__15372\ : std_logic;
signal \N__15371\ : std_logic;
signal \N__15370\ : std_logic;
signal \N__15369\ : std_logic;
signal \N__15366\ : std_logic;
signal \N__15363\ : std_logic;
signal \N__15360\ : std_logic;
signal \N__15357\ : std_logic;
signal \N__15350\ : std_logic;
signal \N__15345\ : std_logic;
signal \N__15332\ : std_logic;
signal \N__15329\ : std_logic;
signal \N__15326\ : std_logic;
signal \N__15325\ : std_logic;
signal \N__15324\ : std_logic;
signal \N__15321\ : std_logic;
signal \N__15318\ : std_logic;
signal \N__15317\ : std_logic;
signal \N__15316\ : std_logic;
signal \N__15315\ : std_logic;
signal \N__15312\ : std_logic;
signal \N__15301\ : std_logic;
signal \N__15296\ : std_logic;
signal \N__15293\ : std_logic;
signal \N__15290\ : std_logic;
signal \N__15287\ : std_logic;
signal \N__15284\ : std_logic;
signal \N__15281\ : std_logic;
signal \N__15278\ : std_logic;
signal \N__15275\ : std_logic;
signal \N__15274\ : std_logic;
signal \N__15271\ : std_logic;
signal \N__15268\ : std_logic;
signal \N__15263\ : std_logic;
signal \N__15260\ : std_logic;
signal \N__15257\ : std_logic;
signal \N__15254\ : std_logic;
signal \N__15251\ : std_logic;
signal \N__15248\ : std_logic;
signal \N__15245\ : std_logic;
signal \N__15242\ : std_logic;
signal \N__15239\ : std_logic;
signal \N__15236\ : std_logic;
signal \N__15235\ : std_logic;
signal \N__15234\ : std_logic;
signal \N__15231\ : std_logic;
signal \N__15228\ : std_logic;
signal \N__15225\ : std_logic;
signal \N__15224\ : std_logic;
signal \N__15219\ : std_logic;
signal \N__15216\ : std_logic;
signal \N__15215\ : std_logic;
signal \N__15214\ : std_logic;
signal \N__15213\ : std_logic;
signal \N__15210\ : std_logic;
signal \N__15207\ : std_logic;
signal \N__15204\ : std_logic;
signal \N__15197\ : std_logic;
signal \N__15194\ : std_logic;
signal \N__15185\ : std_logic;
signal \N__15184\ : std_logic;
signal \N__15183\ : std_logic;
signal \N__15182\ : std_logic;
signal \N__15181\ : std_logic;
signal \N__15180\ : std_logic;
signal \N__15177\ : std_logic;
signal \N__15174\ : std_logic;
signal \N__15165\ : std_logic;
signal \N__15162\ : std_logic;
signal \N__15157\ : std_logic;
signal \N__15154\ : std_logic;
signal \N__15151\ : std_logic;
signal \N__15146\ : std_logic;
signal \N__15145\ : std_logic;
signal \N__15140\ : std_logic;
signal \N__15139\ : std_logic;
signal \N__15138\ : std_logic;
signal \N__15135\ : std_logic;
signal \N__15132\ : std_logic;
signal \N__15129\ : std_logic;
signal \N__15126\ : std_logic;
signal \N__15119\ : std_logic;
signal \N__15116\ : std_logic;
signal \N__15113\ : std_logic;
signal \N__15110\ : std_logic;
signal \N__15107\ : std_logic;
signal \N__15104\ : std_logic;
signal \N__15103\ : std_logic;
signal \N__15100\ : std_logic;
signal \N__15097\ : std_logic;
signal \N__15094\ : std_logic;
signal \N__15091\ : std_logic;
signal \N__15086\ : std_logic;
signal \N__15083\ : std_logic;
signal \N__15080\ : std_logic;
signal \N__15077\ : std_logic;
signal \N__15074\ : std_logic;
signal \N__15073\ : std_logic;
signal \N__15070\ : std_logic;
signal \N__15067\ : std_logic;
signal \N__15062\ : std_logic;
signal \N__15061\ : std_logic;
signal \N__15060\ : std_logic;
signal \N__15059\ : std_logic;
signal \N__15058\ : std_logic;
signal \N__15055\ : std_logic;
signal \N__15054\ : std_logic;
signal \N__15053\ : std_logic;
signal \N__15046\ : std_logic;
signal \N__15043\ : std_logic;
signal \N__15036\ : std_logic;
signal \N__15029\ : std_logic;
signal \N__15028\ : std_logic;
signal \N__15027\ : std_logic;
signal \N__15026\ : std_logic;
signal \N__15023\ : std_logic;
signal \N__15022\ : std_logic;
signal \N__15021\ : std_logic;
signal \N__15020\ : std_logic;
signal \N__15017\ : std_logic;
signal \N__15008\ : std_logic;
signal \N__15003\ : std_logic;
signal \N__14998\ : std_logic;
signal \N__14993\ : std_logic;
signal \N__14990\ : std_logic;
signal \N__14989\ : std_logic;
signal \N__14988\ : std_logic;
signal \N__14987\ : std_logic;
signal \N__14986\ : std_logic;
signal \N__14985\ : std_logic;
signal \N__14984\ : std_logic;
signal \N__14981\ : std_logic;
signal \N__14978\ : std_logic;
signal \N__14975\ : std_logic;
signal \N__14966\ : std_logic;
signal \N__14957\ : std_logic;
signal \N__14956\ : std_logic;
signal \N__14955\ : std_logic;
signal \N__14954\ : std_logic;
signal \N__14953\ : std_logic;
signal \N__14952\ : std_logic;
signal \N__14949\ : std_logic;
signal \N__14942\ : std_logic;
signal \N__14939\ : std_logic;
signal \N__14936\ : std_logic;
signal \N__14927\ : std_logic;
signal \N__14926\ : std_logic;
signal \N__14925\ : std_logic;
signal \N__14924\ : std_logic;
signal \N__14919\ : std_logic;
signal \N__14916\ : std_logic;
signal \N__14913\ : std_logic;
signal \N__14906\ : std_logic;
signal \N__14905\ : std_logic;
signal \N__14902\ : std_logic;
signal \N__14899\ : std_logic;
signal \N__14898\ : std_logic;
signal \N__14897\ : std_logic;
signal \N__14892\ : std_logic;
signal \N__14889\ : std_logic;
signal \N__14886\ : std_logic;
signal \N__14883\ : std_logic;
signal \N__14880\ : std_logic;
signal \N__14873\ : std_logic;
signal \N__14872\ : std_logic;
signal \N__14869\ : std_logic;
signal \N__14866\ : std_logic;
signal \N__14863\ : std_logic;
signal \N__14860\ : std_logic;
signal \N__14859\ : std_logic;
signal \N__14858\ : std_logic;
signal \N__14857\ : std_logic;
signal \N__14856\ : std_logic;
signal \N__14853\ : std_logic;
signal \N__14850\ : std_logic;
signal \N__14847\ : std_logic;
signal \N__14844\ : std_logic;
signal \N__14839\ : std_logic;
signal \N__14834\ : std_logic;
signal \N__14825\ : std_logic;
signal \N__14824\ : std_logic;
signal \N__14821\ : std_logic;
signal \N__14820\ : std_logic;
signal \N__14817\ : std_logic;
signal \N__14814\ : std_logic;
signal \N__14811\ : std_logic;
signal \N__14808\ : std_logic;
signal \N__14801\ : std_logic;
signal \N__14798\ : std_logic;
signal \N__14797\ : std_logic;
signal \N__14796\ : std_logic;
signal \N__14795\ : std_logic;
signal \N__14794\ : std_logic;
signal \N__14793\ : std_logic;
signal \N__14792\ : std_logic;
signal \N__14791\ : std_logic;
signal \N__14788\ : std_logic;
signal \N__14787\ : std_logic;
signal \N__14786\ : std_logic;
signal \N__14785\ : std_logic;
signal \N__14782\ : std_logic;
signal \N__14781\ : std_logic;
signal \N__14778\ : std_logic;
signal \N__14769\ : std_logic;
signal \N__14766\ : std_logic;
signal \N__14763\ : std_logic;
signal \N__14756\ : std_logic;
signal \N__14753\ : std_logic;
signal \N__14750\ : std_logic;
signal \N__14747\ : std_logic;
signal \N__14744\ : std_logic;
signal \N__14741\ : std_logic;
signal \N__14736\ : std_logic;
signal \N__14731\ : std_logic;
signal \N__14728\ : std_logic;
signal \N__14725\ : std_logic;
signal \N__14718\ : std_logic;
signal \N__14713\ : std_logic;
signal \N__14710\ : std_logic;
signal \N__14705\ : std_logic;
signal \N__14704\ : std_logic;
signal \N__14701\ : std_logic;
signal \N__14698\ : std_logic;
signal \N__14695\ : std_logic;
signal \N__14694\ : std_logic;
signal \N__14693\ : std_logic;
signal \N__14690\ : std_logic;
signal \N__14687\ : std_logic;
signal \N__14684\ : std_logic;
signal \N__14681\ : std_logic;
signal \N__14678\ : std_logic;
signal \N__14675\ : std_logic;
signal \N__14670\ : std_logic;
signal \N__14663\ : std_logic;
signal \N__14660\ : std_logic;
signal \N__14659\ : std_logic;
signal \N__14658\ : std_logic;
signal \N__14655\ : std_logic;
signal \N__14652\ : std_logic;
signal \N__14649\ : std_logic;
signal \N__14648\ : std_logic;
signal \N__14643\ : std_logic;
signal \N__14640\ : std_logic;
signal \N__14637\ : std_logic;
signal \N__14634\ : std_logic;
signal \N__14631\ : std_logic;
signal \N__14624\ : std_logic;
signal \N__14621\ : std_logic;
signal \N__14618\ : std_logic;
signal \N__14615\ : std_logic;
signal \N__14612\ : std_logic;
signal \N__14609\ : std_logic;
signal \N__14606\ : std_logic;
signal \N__14605\ : std_logic;
signal \N__14602\ : std_logic;
signal \N__14599\ : std_logic;
signal \N__14594\ : std_logic;
signal \N__14591\ : std_logic;
signal \N__14588\ : std_logic;
signal \N__14585\ : std_logic;
signal \N__14584\ : std_logic;
signal \N__14583\ : std_logic;
signal \N__14576\ : std_logic;
signal \N__14573\ : std_logic;
signal \N__14570\ : std_logic;
signal \N__14567\ : std_logic;
signal \N__14564\ : std_logic;
signal \N__14561\ : std_logic;
signal \N__14558\ : std_logic;
signal \N__14555\ : std_logic;
signal \N__14552\ : std_logic;
signal \N__14549\ : std_logic;
signal \N__14546\ : std_logic;
signal \N__14545\ : std_logic;
signal \N__14542\ : std_logic;
signal \N__14539\ : std_logic;
signal \N__14536\ : std_logic;
signal \N__14533\ : std_logic;
signal \N__14530\ : std_logic;
signal \N__14525\ : std_logic;
signal \N__14522\ : std_logic;
signal \N__14519\ : std_logic;
signal \N__14516\ : std_logic;
signal \N__14513\ : std_logic;
signal \N__14510\ : std_logic;
signal \N__14509\ : std_logic;
signal \N__14506\ : std_logic;
signal \N__14503\ : std_logic;
signal \N__14498\ : std_logic;
signal \N__14495\ : std_logic;
signal \N__14492\ : std_logic;
signal \N__14489\ : std_logic;
signal \N__14486\ : std_logic;
signal \N__14485\ : std_logic;
signal \N__14482\ : std_logic;
signal \N__14479\ : std_logic;
signal \N__14476\ : std_logic;
signal \N__14473\ : std_logic;
signal \N__14470\ : std_logic;
signal \N__14465\ : std_logic;
signal \N__14462\ : std_logic;
signal \N__14459\ : std_logic;
signal \N__14456\ : std_logic;
signal \N__14455\ : std_logic;
signal \N__14452\ : std_logic;
signal \N__14449\ : std_logic;
signal \N__14446\ : std_logic;
signal \N__14443\ : std_logic;
signal \N__14440\ : std_logic;
signal \N__14437\ : std_logic;
signal \N__14434\ : std_logic;
signal \N__14429\ : std_logic;
signal \N__14426\ : std_logic;
signal \N__14423\ : std_logic;
signal \N__14420\ : std_logic;
signal \N__14419\ : std_logic;
signal \N__14418\ : std_logic;
signal \N__14417\ : std_logic;
signal \N__14416\ : std_logic;
signal \N__14415\ : std_logic;
signal \N__14414\ : std_logic;
signal \N__14413\ : std_logic;
signal \N__14410\ : std_logic;
signal \N__14405\ : std_logic;
signal \N__14394\ : std_logic;
signal \N__14389\ : std_logic;
signal \N__14386\ : std_logic;
signal \N__14383\ : std_logic;
signal \N__14380\ : std_logic;
signal \N__14375\ : std_logic;
signal \N__14372\ : std_logic;
signal \N__14371\ : std_logic;
signal \N__14368\ : std_logic;
signal \N__14365\ : std_logic;
signal \N__14362\ : std_logic;
signal \N__14359\ : std_logic;
signal \N__14356\ : std_logic;
signal \N__14353\ : std_logic;
signal \N__14348\ : std_logic;
signal \N__14347\ : std_logic;
signal \N__14346\ : std_logic;
signal \N__14345\ : std_logic;
signal \N__14344\ : std_logic;
signal \N__14343\ : std_logic;
signal \N__14342\ : std_logic;
signal \N__14341\ : std_logic;
signal \N__14340\ : std_logic;
signal \N__14339\ : std_logic;
signal \N__14328\ : std_logic;
signal \N__14323\ : std_logic;
signal \N__14322\ : std_logic;
signal \N__14321\ : std_logic;
signal \N__14314\ : std_logic;
signal \N__14311\ : std_logic;
signal \N__14308\ : std_logic;
signal \N__14303\ : std_logic;
signal \N__14300\ : std_logic;
signal \N__14299\ : std_logic;
signal \N__14298\ : std_logic;
signal \N__14295\ : std_logic;
signal \N__14292\ : std_logic;
signal \N__14287\ : std_logic;
signal \N__14282\ : std_logic;
signal \N__14279\ : std_logic;
signal \N__14270\ : std_logic;
signal \N__14269\ : std_logic;
signal \N__14266\ : std_logic;
signal \N__14261\ : std_logic;
signal \N__14258\ : std_logic;
signal \N__14255\ : std_logic;
signal \N__14254\ : std_logic;
signal \N__14251\ : std_logic;
signal \N__14248\ : std_logic;
signal \N__14243\ : std_logic;
signal \N__14242\ : std_logic;
signal \N__14241\ : std_logic;
signal \N__14238\ : std_logic;
signal \N__14235\ : std_logic;
signal \N__14232\ : std_logic;
signal \N__14231\ : std_logic;
signal \N__14228\ : std_logic;
signal \N__14225\ : std_logic;
signal \N__14222\ : std_logic;
signal \N__14219\ : std_logic;
signal \N__14216\ : std_logic;
signal \N__14209\ : std_logic;
signal \N__14204\ : std_logic;
signal \N__14201\ : std_logic;
signal \N__14200\ : std_logic;
signal \N__14199\ : std_logic;
signal \N__14198\ : std_logic;
signal \N__14195\ : std_logic;
signal \N__14192\ : std_logic;
signal \N__14189\ : std_logic;
signal \N__14186\ : std_logic;
signal \N__14181\ : std_logic;
signal \N__14178\ : std_logic;
signal \N__14171\ : std_logic;
signal \N__14168\ : std_logic;
signal \N__14165\ : std_logic;
signal \N__14162\ : std_logic;
signal \N__14159\ : std_logic;
signal \N__14156\ : std_logic;
signal \N__14153\ : std_logic;
signal \N__14150\ : std_logic;
signal \N__14147\ : std_logic;
signal \N__14144\ : std_logic;
signal \N__14141\ : std_logic;
signal \N__14138\ : std_logic;
signal \N__14135\ : std_logic;
signal \N__14132\ : std_logic;
signal \N__14129\ : std_logic;
signal \N__14126\ : std_logic;
signal \N__14123\ : std_logic;
signal \N__14120\ : std_logic;
signal \N__14117\ : std_logic;
signal \N__14114\ : std_logic;
signal \N__14111\ : std_logic;
signal \N__14108\ : std_logic;
signal \N__14105\ : std_logic;
signal \N__14102\ : std_logic;
signal \N__14099\ : std_logic;
signal \N__14096\ : std_logic;
signal \N__14095\ : std_logic;
signal \N__14094\ : std_logic;
signal \N__14089\ : std_logic;
signal \N__14086\ : std_logic;
signal \N__14083\ : std_logic;
signal \N__14078\ : std_logic;
signal \N__14075\ : std_logic;
signal \N__14072\ : std_logic;
signal \N__14069\ : std_logic;
signal \N__14066\ : std_logic;
signal \N__14063\ : std_logic;
signal \N__14060\ : std_logic;
signal \N__14059\ : std_logic;
signal \N__14056\ : std_logic;
signal \N__14053\ : std_logic;
signal \N__14050\ : std_logic;
signal \N__14047\ : std_logic;
signal \N__14044\ : std_logic;
signal \N__14041\ : std_logic;
signal \N__14038\ : std_logic;
signal \N__14033\ : std_logic;
signal \N__14030\ : std_logic;
signal \N__14027\ : std_logic;
signal \N__14026\ : std_logic;
signal \N__14023\ : std_logic;
signal \N__14020\ : std_logic;
signal \N__14017\ : std_logic;
signal \N__14014\ : std_logic;
signal \N__14011\ : std_logic;
signal \N__14006\ : std_logic;
signal \N__14003\ : std_logic;
signal \N__14000\ : std_logic;
signal \N__13999\ : std_logic;
signal \N__13996\ : std_logic;
signal \N__13993\ : std_logic;
signal \N__13990\ : std_logic;
signal \N__13987\ : std_logic;
signal \N__13984\ : std_logic;
signal \N__13981\ : std_logic;
signal \N__13978\ : std_logic;
signal \N__13973\ : std_logic;
signal \N__13970\ : std_logic;
signal \N__13967\ : std_logic;
signal \N__13964\ : std_logic;
signal \N__13963\ : std_logic;
signal \N__13962\ : std_logic;
signal \N__13959\ : std_logic;
signal \N__13954\ : std_logic;
signal \N__13949\ : std_logic;
signal \N__13946\ : std_logic;
signal \N__13943\ : std_logic;
signal \N__13940\ : std_logic;
signal \N__13937\ : std_logic;
signal \N__13936\ : std_logic;
signal \N__13933\ : std_logic;
signal \N__13930\ : std_logic;
signal \N__13927\ : std_logic;
signal \N__13924\ : std_logic;
signal \N__13919\ : std_logic;
signal \N__13916\ : std_logic;
signal \N__13913\ : std_logic;
signal \N__13912\ : std_logic;
signal \N__13909\ : std_logic;
signal \N__13906\ : std_logic;
signal \N__13903\ : std_logic;
signal \N__13900\ : std_logic;
signal \N__13895\ : std_logic;
signal \N__13894\ : std_logic;
signal \N__13893\ : std_logic;
signal \N__13892\ : std_logic;
signal \N__13889\ : std_logic;
signal \N__13886\ : std_logic;
signal \N__13881\ : std_logic;
signal \N__13874\ : std_logic;
signal \N__13871\ : std_logic;
signal \N__13868\ : std_logic;
signal \N__13867\ : std_logic;
signal \N__13864\ : std_logic;
signal \N__13861\ : std_logic;
signal \N__13858\ : std_logic;
signal \N__13853\ : std_logic;
signal \N__13852\ : std_logic;
signal \N__13851\ : std_logic;
signal \N__13848\ : std_logic;
signal \N__13845\ : std_logic;
signal \N__13842\ : std_logic;
signal \N__13835\ : std_logic;
signal \N__13832\ : std_logic;
signal \N__13829\ : std_logic;
signal \N__13828\ : std_logic;
signal \N__13823\ : std_logic;
signal \N__13820\ : std_logic;
signal \N__13817\ : std_logic;
signal \N__13816\ : std_logic;
signal \N__13811\ : std_logic;
signal \N__13808\ : std_logic;
signal \N__13805\ : std_logic;
signal \N__13804\ : std_logic;
signal \N__13803\ : std_logic;
signal \N__13802\ : std_logic;
signal \N__13801\ : std_logic;
signal \N__13800\ : std_logic;
signal \N__13797\ : std_logic;
signal \N__13796\ : std_logic;
signal \N__13793\ : std_logic;
signal \N__13790\ : std_logic;
signal \N__13787\ : std_logic;
signal \N__13778\ : std_logic;
signal \N__13769\ : std_logic;
signal \N__13766\ : std_logic;
signal \N__13763\ : std_logic;
signal \N__13760\ : std_logic;
signal \N__13759\ : std_logic;
signal \N__13758\ : std_logic;
signal \N__13757\ : std_logic;
signal \N__13754\ : std_logic;
signal \N__13751\ : std_logic;
signal \N__13746\ : std_logic;
signal \N__13745\ : std_logic;
signal \N__13744\ : std_logic;
signal \N__13743\ : std_logic;
signal \N__13742\ : std_logic;
signal \N__13741\ : std_logic;
signal \N__13734\ : std_logic;
signal \N__13723\ : std_logic;
signal \N__13718\ : std_logic;
signal \N__13715\ : std_logic;
signal \N__13712\ : std_logic;
signal \N__13709\ : std_logic;
signal \N__13706\ : std_logic;
signal \N__13703\ : std_logic;
signal \N__13700\ : std_logic;
signal \N__13697\ : std_logic;
signal \N__13694\ : std_logic;
signal \N__13691\ : std_logic;
signal \N__13688\ : std_logic;
signal \N__13687\ : std_logic;
signal \N__13686\ : std_logic;
signal \N__13683\ : std_logic;
signal \N__13680\ : std_logic;
signal \N__13675\ : std_logic;
signal \N__13670\ : std_logic;
signal \N__13669\ : std_logic;
signal \N__13668\ : std_logic;
signal \N__13667\ : std_logic;
signal \N__13666\ : std_logic;
signal \N__13665\ : std_logic;
signal \N__13662\ : std_logic;
signal \N__13659\ : std_logic;
signal \N__13650\ : std_logic;
signal \N__13643\ : std_logic;
signal \N__13642\ : std_logic;
signal \N__13639\ : std_logic;
signal \N__13638\ : std_logic;
signal \N__13635\ : std_logic;
signal \N__13632\ : std_logic;
signal \N__13629\ : std_logic;
signal \N__13626\ : std_logic;
signal \N__13623\ : std_logic;
signal \N__13620\ : std_logic;
signal \N__13619\ : std_logic;
signal \N__13612\ : std_logic;
signal \N__13609\ : std_logic;
signal \N__13604\ : std_logic;
signal \N__13603\ : std_logic;
signal \N__13602\ : std_logic;
signal \N__13601\ : std_logic;
signal \N__13598\ : std_logic;
signal \N__13595\ : std_logic;
signal \N__13592\ : std_logic;
signal \N__13589\ : std_logic;
signal \N__13586\ : std_logic;
signal \N__13583\ : std_logic;
signal \N__13578\ : std_logic;
signal \N__13575\ : std_logic;
signal \N__13568\ : std_logic;
signal \N__13565\ : std_logic;
signal \N__13562\ : std_logic;
signal \N__13559\ : std_logic;
signal \N__13556\ : std_logic;
signal \N__13553\ : std_logic;
signal \N__13552\ : std_logic;
signal \N__13549\ : std_logic;
signal \N__13546\ : std_logic;
signal \N__13545\ : std_logic;
signal \N__13542\ : std_logic;
signal \N__13539\ : std_logic;
signal \N__13536\ : std_logic;
signal \N__13535\ : std_logic;
signal \N__13532\ : std_logic;
signal \N__13529\ : std_logic;
signal \N__13526\ : std_logic;
signal \N__13523\ : std_logic;
signal \N__13514\ : std_logic;
signal \N__13513\ : std_logic;
signal \N__13510\ : std_logic;
signal \N__13509\ : std_logic;
signal \N__13508\ : std_logic;
signal \N__13505\ : std_logic;
signal \N__13502\ : std_logic;
signal \N__13499\ : std_logic;
signal \N__13496\ : std_logic;
signal \N__13493\ : std_logic;
signal \N__13488\ : std_logic;
signal \N__13481\ : std_logic;
signal \N__13480\ : std_logic;
signal \N__13477\ : std_logic;
signal \N__13474\ : std_logic;
signal \N__13471\ : std_logic;
signal \N__13468\ : std_logic;
signal \N__13463\ : std_logic;
signal \N__13460\ : std_logic;
signal \N__13459\ : std_logic;
signal \N__13456\ : std_logic;
signal \N__13453\ : std_logic;
signal \N__13450\ : std_logic;
signal \N__13447\ : std_logic;
signal \N__13444\ : std_logic;
signal \N__13441\ : std_logic;
signal \N__13436\ : std_logic;
signal \N__13433\ : std_logic;
signal \N__13430\ : std_logic;
signal \N__13427\ : std_logic;
signal \N__13424\ : std_logic;
signal \N__13421\ : std_logic;
signal \N__13418\ : std_logic;
signal \N__13415\ : std_logic;
signal \N__13412\ : std_logic;
signal \N__13411\ : std_logic;
signal \N__13408\ : std_logic;
signal \N__13405\ : std_logic;
signal \N__13402\ : std_logic;
signal \N__13399\ : std_logic;
signal \N__13394\ : std_logic;
signal \N__13391\ : std_logic;
signal \N__13388\ : std_logic;
signal \N__13385\ : std_logic;
signal \N__13382\ : std_logic;
signal \N__13381\ : std_logic;
signal \N__13380\ : std_logic;
signal \N__13379\ : std_logic;
signal \N__13376\ : std_logic;
signal \N__13373\ : std_logic;
signal \N__13370\ : std_logic;
signal \N__13365\ : std_logic;
signal \N__13358\ : std_logic;
signal \N__13357\ : std_logic;
signal \N__13356\ : std_logic;
signal \N__13355\ : std_logic;
signal \N__13352\ : std_logic;
signal \N__13351\ : std_logic;
signal \N__13350\ : std_logic;
signal \N__13349\ : std_logic;
signal \N__13348\ : std_logic;
signal \N__13347\ : std_logic;
signal \N__13344\ : std_logic;
signal \N__13339\ : std_logic;
signal \N__13336\ : std_logic;
signal \N__13333\ : std_logic;
signal \N__13330\ : std_logic;
signal \N__13325\ : std_logic;
signal \N__13322\ : std_logic;
signal \N__13317\ : std_logic;
signal \N__13304\ : std_logic;
signal \N__13303\ : std_logic;
signal \N__13302\ : std_logic;
signal \N__13301\ : std_logic;
signal \N__13300\ : std_logic;
signal \N__13297\ : std_logic;
signal \N__13294\ : std_logic;
signal \N__13287\ : std_logic;
signal \N__13280\ : std_logic;
signal \N__13277\ : std_logic;
signal \N__13274\ : std_logic;
signal \N__13271\ : std_logic;
signal \N__13268\ : std_logic;
signal \N__13267\ : std_logic;
signal \N__13266\ : std_logic;
signal \N__13263\ : std_logic;
signal \N__13260\ : std_logic;
signal \N__13257\ : std_logic;
signal \N__13254\ : std_logic;
signal \N__13251\ : std_logic;
signal \N__13248\ : std_logic;
signal \N__13241\ : std_logic;
signal \N__13238\ : std_logic;
signal \N__13237\ : std_logic;
signal \N__13234\ : std_logic;
signal \N__13233\ : std_logic;
signal \N__13232\ : std_logic;
signal \N__13231\ : std_logic;
signal \N__13230\ : std_logic;
signal \N__13229\ : std_logic;
signal \N__13228\ : std_logic;
signal \N__13227\ : std_logic;
signal \N__13224\ : std_logic;
signal \N__13223\ : std_logic;
signal \N__13220\ : std_logic;
signal \N__13219\ : std_logic;
signal \N__13218\ : std_logic;
signal \N__13215\ : std_logic;
signal \N__13210\ : std_logic;
signal \N__13207\ : std_logic;
signal \N__13204\ : std_logic;
signal \N__13199\ : std_logic;
signal \N__13196\ : std_logic;
signal \N__13193\ : std_logic;
signal \N__13190\ : std_logic;
signal \N__13185\ : std_logic;
signal \N__13180\ : std_logic;
signal \N__13173\ : std_logic;
signal \N__13170\ : std_logic;
signal \N__13163\ : std_logic;
signal \N__13158\ : std_logic;
signal \N__13151\ : std_logic;
signal \N__13148\ : std_logic;
signal \N__13145\ : std_logic;
signal \N__13142\ : std_logic;
signal \N__13141\ : std_logic;
signal \N__13138\ : std_logic;
signal \N__13135\ : std_logic;
signal \N__13130\ : std_logic;
signal \N__13127\ : std_logic;
signal \N__13124\ : std_logic;
signal \N__13121\ : std_logic;
signal \N__13118\ : std_logic;
signal \N__13115\ : std_logic;
signal \N__13112\ : std_logic;
signal \N__13109\ : std_logic;
signal \N__13106\ : std_logic;
signal \N__13103\ : std_logic;
signal \N__13102\ : std_logic;
signal \N__13099\ : std_logic;
signal \N__13096\ : std_logic;
signal \N__13095\ : std_logic;
signal \N__13092\ : std_logic;
signal \N__13089\ : std_logic;
signal \N__13086\ : std_logic;
signal \N__13085\ : std_logic;
signal \N__13080\ : std_logic;
signal \N__13077\ : std_logic;
signal \N__13074\ : std_logic;
signal \N__13067\ : std_logic;
signal \N__13064\ : std_logic;
signal \N__13061\ : std_logic;
signal \N__13060\ : std_logic;
signal \N__13059\ : std_logic;
signal \N__13058\ : std_logic;
signal \N__13055\ : std_logic;
signal \N__13052\ : std_logic;
signal \N__13049\ : std_logic;
signal \N__13046\ : std_logic;
signal \N__13041\ : std_logic;
signal \N__13038\ : std_logic;
signal \N__13031\ : std_logic;
signal \N__13028\ : std_logic;
signal \N__13027\ : std_logic;
signal \N__13024\ : std_logic;
signal \N__13021\ : std_logic;
signal \N__13020\ : std_logic;
signal \N__13017\ : std_logic;
signal \N__13014\ : std_logic;
signal \N__13011\ : std_logic;
signal \N__13010\ : std_logic;
signal \N__13005\ : std_logic;
signal \N__13002\ : std_logic;
signal \N__12999\ : std_logic;
signal \N__12992\ : std_logic;
signal \N__12991\ : std_logic;
signal \N__12988\ : std_logic;
signal \N__12987\ : std_logic;
signal \N__12986\ : std_logic;
signal \N__12983\ : std_logic;
signal \N__12980\ : std_logic;
signal \N__12977\ : std_logic;
signal \N__12974\ : std_logic;
signal \N__12971\ : std_logic;
signal \N__12966\ : std_logic;
signal \N__12959\ : std_logic;
signal \N__12958\ : std_logic;
signal \N__12955\ : std_logic;
signal \N__12952\ : std_logic;
signal \N__12951\ : std_logic;
signal \N__12948\ : std_logic;
signal \N__12945\ : std_logic;
signal \N__12942\ : std_logic;
signal \N__12941\ : std_logic;
signal \N__12936\ : std_logic;
signal \N__12933\ : std_logic;
signal \N__12930\ : std_logic;
signal \N__12923\ : std_logic;
signal \N__12920\ : std_logic;
signal \N__12919\ : std_logic;
signal \N__12916\ : std_logic;
signal \N__12915\ : std_logic;
signal \N__12914\ : std_logic;
signal \N__12911\ : std_logic;
signal \N__12908\ : std_logic;
signal \N__12905\ : std_logic;
signal \N__12902\ : std_logic;
signal \N__12899\ : std_logic;
signal \N__12894\ : std_logic;
signal \N__12887\ : std_logic;
signal \N__12886\ : std_logic;
signal \N__12883\ : std_logic;
signal \N__12880\ : std_logic;
signal \N__12879\ : std_logic;
signal \N__12876\ : std_logic;
signal \N__12873\ : std_logic;
signal \N__12870\ : std_logic;
signal \N__12869\ : std_logic;
signal \N__12864\ : std_logic;
signal \N__12861\ : std_logic;
signal \N__12858\ : std_logic;
signal \N__12851\ : std_logic;
signal \N__12848\ : std_logic;
signal \N__12847\ : std_logic;
signal \N__12846\ : std_logic;
signal \N__12845\ : std_logic;
signal \N__12842\ : std_logic;
signal \N__12839\ : std_logic;
signal \N__12836\ : std_logic;
signal \N__12833\ : std_logic;
signal \N__12830\ : std_logic;
signal \N__12827\ : std_logic;
signal \N__12824\ : std_logic;
signal \N__12821\ : std_logic;
signal \N__12812\ : std_logic;
signal \N__12809\ : std_logic;
signal \N__12808\ : std_logic;
signal \N__12807\ : std_logic;
signal \N__12804\ : std_logic;
signal \N__12801\ : std_logic;
signal \N__12798\ : std_logic;
signal \N__12791\ : std_logic;
signal \N__12788\ : std_logic;
signal \N__12785\ : std_logic;
signal \N__12784\ : std_logic;
signal \N__12783\ : std_logic;
signal \N__12780\ : std_logic;
signal \N__12777\ : std_logic;
signal \N__12774\ : std_logic;
signal \N__12767\ : std_logic;
signal \N__12764\ : std_logic;
signal \N__12763\ : std_logic;
signal \N__12762\ : std_logic;
signal \N__12759\ : std_logic;
signal \N__12756\ : std_logic;
signal \N__12753\ : std_logic;
signal \N__12750\ : std_logic;
signal \N__12747\ : std_logic;
signal \N__12744\ : std_logic;
signal \N__12737\ : std_logic;
signal \N__12736\ : std_logic;
signal \N__12735\ : std_logic;
signal \N__12732\ : std_logic;
signal \N__12729\ : std_logic;
signal \N__12726\ : std_logic;
signal \N__12723\ : std_logic;
signal \N__12720\ : std_logic;
signal \N__12717\ : std_logic;
signal \N__12714\ : std_logic;
signal \N__12707\ : std_logic;
signal \N__12704\ : std_logic;
signal \N__12703\ : std_logic;
signal \N__12702\ : std_logic;
signal \N__12699\ : std_logic;
signal \N__12696\ : std_logic;
signal \N__12693\ : std_logic;
signal \N__12690\ : std_logic;
signal \N__12687\ : std_logic;
signal \N__12684\ : std_logic;
signal \N__12677\ : std_logic;
signal \N__12676\ : std_logic;
signal \N__12675\ : std_logic;
signal \N__12672\ : std_logic;
signal \N__12669\ : std_logic;
signal \N__12666\ : std_logic;
signal \N__12663\ : std_logic;
signal \N__12660\ : std_logic;
signal \N__12657\ : std_logic;
signal \N__12654\ : std_logic;
signal \N__12647\ : std_logic;
signal \N__12644\ : std_logic;
signal \N__12643\ : std_logic;
signal \N__12642\ : std_logic;
signal \N__12639\ : std_logic;
signal \N__12636\ : std_logic;
signal \N__12633\ : std_logic;
signal \N__12630\ : std_logic;
signal \N__12627\ : std_logic;
signal \N__12624\ : std_logic;
signal \N__12617\ : std_logic;
signal \N__12614\ : std_logic;
signal \N__12613\ : std_logic;
signal \N__12612\ : std_logic;
signal \N__12609\ : std_logic;
signal \N__12606\ : std_logic;
signal \N__12603\ : std_logic;
signal \N__12600\ : std_logic;
signal \N__12597\ : std_logic;
signal \N__12594\ : std_logic;
signal \N__12587\ : std_logic;
signal \N__12584\ : std_logic;
signal \N__12583\ : std_logic;
signal \N__12582\ : std_logic;
signal \N__12579\ : std_logic;
signal \N__12576\ : std_logic;
signal \N__12573\ : std_logic;
signal \N__12570\ : std_logic;
signal \N__12567\ : std_logic;
signal \N__12564\ : std_logic;
signal \N__12557\ : std_logic;
signal \N__12556\ : std_logic;
signal \N__12553\ : std_logic;
signal \N__12550\ : std_logic;
signal \N__12545\ : std_logic;
signal \N__12542\ : std_logic;
signal \N__12541\ : std_logic;
signal \N__12538\ : std_logic;
signal \N__12535\ : std_logic;
signal \N__12532\ : std_logic;
signal \N__12529\ : std_logic;
signal \N__12526\ : std_logic;
signal \N__12523\ : std_logic;
signal \N__12520\ : std_logic;
signal \N__12515\ : std_logic;
signal \N__12512\ : std_logic;
signal \N__12509\ : std_logic;
signal \N__12506\ : std_logic;
signal \N__12503\ : std_logic;
signal \N__12500\ : std_logic;
signal \N__12499\ : std_logic;
signal \N__12498\ : std_logic;
signal \N__12497\ : std_logic;
signal \N__12496\ : std_logic;
signal \N__12495\ : std_logic;
signal \N__12494\ : std_logic;
signal \N__12493\ : std_logic;
signal \N__12492\ : std_logic;
signal \N__12487\ : std_logic;
signal \N__12474\ : std_logic;
signal \N__12473\ : std_logic;
signal \N__12470\ : std_logic;
signal \N__12467\ : std_logic;
signal \N__12464\ : std_logic;
signal \N__12461\ : std_logic;
signal \N__12452\ : std_logic;
signal \N__12449\ : std_logic;
signal \N__12448\ : std_logic;
signal \N__12443\ : std_logic;
signal \N__12440\ : std_logic;
signal \N__12439\ : std_logic;
signal \N__12438\ : std_logic;
signal \N__12437\ : std_logic;
signal \N__12434\ : std_logic;
signal \N__12431\ : std_logic;
signal \N__12428\ : std_logic;
signal \N__12427\ : std_logic;
signal \N__12426\ : std_logic;
signal \N__12423\ : std_logic;
signal \N__12422\ : std_logic;
signal \N__12421\ : std_logic;
signal \N__12418\ : std_logic;
signal \N__12405\ : std_logic;
signal \N__12402\ : std_logic;
signal \N__12395\ : std_logic;
signal \N__12392\ : std_logic;
signal \N__12389\ : std_logic;
signal \N__12386\ : std_logic;
signal \N__12383\ : std_logic;
signal \N__12380\ : std_logic;
signal \N__12377\ : std_logic;
signal \N__12374\ : std_logic;
signal \N__12371\ : std_logic;
signal \N__12368\ : std_logic;
signal \N__12365\ : std_logic;
signal \N__12362\ : std_logic;
signal \N__12359\ : std_logic;
signal \N__12356\ : std_logic;
signal \N__12353\ : std_logic;
signal \N__12350\ : std_logic;
signal \N__12349\ : std_logic;
signal \N__12346\ : std_logic;
signal \N__12343\ : std_logic;
signal \N__12338\ : std_logic;
signal \N__12337\ : std_logic;
signal \N__12334\ : std_logic;
signal \N__12331\ : std_logic;
signal \N__12326\ : std_logic;
signal \N__12325\ : std_logic;
signal \N__12322\ : std_logic;
signal \N__12319\ : std_logic;
signal \N__12314\ : std_logic;
signal \N__12313\ : std_logic;
signal \N__12310\ : std_logic;
signal \N__12307\ : std_logic;
signal \N__12302\ : std_logic;
signal \N__12301\ : std_logic;
signal \N__12298\ : std_logic;
signal \N__12295\ : std_logic;
signal \N__12292\ : std_logic;
signal \N__12287\ : std_logic;
signal \N__12284\ : std_logic;
signal \N__12281\ : std_logic;
signal \N__12278\ : std_logic;
signal \N__12277\ : std_logic;
signal \N__12276\ : std_logic;
signal \N__12273\ : std_logic;
signal \N__12266\ : std_logic;
signal \N__12265\ : std_logic;
signal \N__12264\ : std_logic;
signal \N__12261\ : std_logic;
signal \N__12258\ : std_logic;
signal \N__12255\ : std_logic;
signal \N__12252\ : std_logic;
signal \N__12245\ : std_logic;
signal \N__12242\ : std_logic;
signal \N__12241\ : std_logic;
signal \N__12238\ : std_logic;
signal \N__12237\ : std_logic;
signal \N__12236\ : std_logic;
signal \N__12235\ : std_logic;
signal \N__12234\ : std_logic;
signal \N__12233\ : std_logic;
signal \N__12232\ : std_logic;
signal \N__12229\ : std_logic;
signal \N__12226\ : std_logic;
signal \N__12221\ : std_logic;
signal \N__12216\ : std_logic;
signal \N__12211\ : std_logic;
signal \N__12200\ : std_logic;
signal \N__12199\ : std_logic;
signal \N__12198\ : std_logic;
signal \N__12195\ : std_logic;
signal \N__12194\ : std_logic;
signal \N__12193\ : std_logic;
signal \N__12188\ : std_logic;
signal \N__12181\ : std_logic;
signal \N__12176\ : std_logic;
signal \N__12173\ : std_logic;
signal \N__12172\ : std_logic;
signal \N__12167\ : std_logic;
signal \N__12166\ : std_logic;
signal \N__12165\ : std_logic;
signal \N__12162\ : std_logic;
signal \N__12161\ : std_logic;
signal \N__12160\ : std_logic;
signal \N__12159\ : std_logic;
signal \N__12158\ : std_logic;
signal \N__12157\ : std_logic;
signal \N__12154\ : std_logic;
signal \N__12153\ : std_logic;
signal \N__12150\ : std_logic;
signal \N__12147\ : std_logic;
signal \N__12142\ : std_logic;
signal \N__12135\ : std_logic;
signal \N__12130\ : std_logic;
signal \N__12119\ : std_logic;
signal \N__12118\ : std_logic;
signal \N__12117\ : std_logic;
signal \N__12116\ : std_logic;
signal \N__12115\ : std_logic;
signal \N__12114\ : std_logic;
signal \N__12109\ : std_logic;
signal \N__12100\ : std_logic;
signal \N__12095\ : std_logic;
signal \N__12092\ : std_logic;
signal \N__12089\ : std_logic;
signal \N__12088\ : std_logic;
signal \N__12085\ : std_logic;
signal \N__12082\ : std_logic;
signal \N__12081\ : std_logic;
signal \N__12080\ : std_logic;
signal \N__12079\ : std_logic;
signal \N__12076\ : std_logic;
signal \N__12071\ : std_logic;
signal \N__12066\ : std_logic;
signal \N__12059\ : std_logic;
signal \N__12058\ : std_logic;
signal \N__12057\ : std_logic;
signal \N__12056\ : std_logic;
signal \N__12053\ : std_logic;
signal \N__12050\ : std_logic;
signal \N__12045\ : std_logic;
signal \N__12038\ : std_logic;
signal \N__12035\ : std_logic;
signal \N__12034\ : std_logic;
signal \N__12033\ : std_logic;
signal \N__12030\ : std_logic;
signal \N__12025\ : std_logic;
signal \N__12020\ : std_logic;
signal \N__12017\ : std_logic;
signal \N__12014\ : std_logic;
signal \N__12013\ : std_logic;
signal \N__12012\ : std_logic;
signal \N__12011\ : std_logic;
signal \N__12010\ : std_logic;
signal \N__12009\ : std_logic;
signal \N__12008\ : std_logic;
signal \N__12007\ : std_logic;
signal \N__12004\ : std_logic;
signal \N__11989\ : std_logic;
signal \N__11984\ : std_logic;
signal \N__11981\ : std_logic;
signal \N__11978\ : std_logic;
signal \N__11977\ : std_logic;
signal \N__11976\ : std_logic;
signal \N__11975\ : std_logic;
signal \N__11974\ : std_logic;
signal \N__11973\ : std_logic;
signal \N__11972\ : std_logic;
signal \N__11971\ : std_logic;
signal \N__11968\ : std_logic;
signal \N__11953\ : std_logic;
signal \N__11948\ : std_logic;
signal \N__11947\ : std_logic;
signal \N__11946\ : std_logic;
signal \N__11945\ : std_logic;
signal \N__11944\ : std_logic;
signal \N__11941\ : std_logic;
signal \N__11938\ : std_logic;
signal \N__11935\ : std_logic;
signal \N__11932\ : std_logic;
signal \N__11929\ : std_logic;
signal \N__11926\ : std_logic;
signal \N__11925\ : std_logic;
signal \N__11924\ : std_logic;
signal \N__11923\ : std_logic;
signal \N__11914\ : std_logic;
signal \N__11911\ : std_logic;
signal \N__11908\ : std_logic;
signal \N__11905\ : std_logic;
signal \N__11902\ : std_logic;
signal \N__11897\ : std_logic;
signal \N__11890\ : std_logic;
signal \N__11887\ : std_logic;
signal \N__11882\ : std_logic;
signal \N__11879\ : std_logic;
signal \N__11876\ : std_logic;
signal \N__11873\ : std_logic;
signal \N__11870\ : std_logic;
signal \N__11869\ : std_logic;
signal \N__11868\ : std_logic;
signal \N__11867\ : std_logic;
signal \N__11864\ : std_logic;
signal \N__11857\ : std_logic;
signal \N__11852\ : std_logic;
signal \N__11849\ : std_logic;
signal \N__11846\ : std_logic;
signal \N__11845\ : std_logic;
signal \N__11844\ : std_logic;
signal \N__11841\ : std_logic;
signal \N__11838\ : std_logic;
signal \N__11835\ : std_logic;
signal \N__11834\ : std_logic;
signal \N__11833\ : std_logic;
signal \N__11832\ : std_logic;
signal \N__11829\ : std_logic;
signal \N__11826\ : std_logic;
signal \N__11823\ : std_logic;
signal \N__11816\ : std_logic;
signal \N__11813\ : std_logic;
signal \N__11810\ : std_logic;
signal \N__11801\ : std_logic;
signal \N__11798\ : std_logic;
signal \N__11795\ : std_logic;
signal \N__11794\ : std_logic;
signal \N__11791\ : std_logic;
signal \N__11788\ : std_logic;
signal \N__11787\ : std_logic;
signal \N__11784\ : std_logic;
signal \N__11779\ : std_logic;
signal \N__11776\ : std_logic;
signal \N__11773\ : std_logic;
signal \N__11768\ : std_logic;
signal \N__11765\ : std_logic;
signal \N__11764\ : std_logic;
signal \N__11761\ : std_logic;
signal \N__11760\ : std_logic;
signal \N__11759\ : std_logic;
signal \N__11756\ : std_logic;
signal \N__11755\ : std_logic;
signal \N__11752\ : std_logic;
signal \N__11747\ : std_logic;
signal \N__11742\ : std_logic;
signal \N__11735\ : std_logic;
signal \N__11732\ : std_logic;
signal \N__11729\ : std_logic;
signal \N__11726\ : std_logic;
signal \N__11723\ : std_logic;
signal \N__11720\ : std_logic;
signal \N__11717\ : std_logic;
signal \N__11714\ : std_logic;
signal \N__11713\ : std_logic;
signal \N__11710\ : std_logic;
signal \N__11707\ : std_logic;
signal \N__11706\ : std_logic;
signal \N__11701\ : std_logic;
signal \N__11698\ : std_logic;
signal \N__11695\ : std_logic;
signal \N__11690\ : std_logic;
signal \N__11689\ : std_logic;
signal \N__11688\ : std_logic;
signal \N__11683\ : std_logic;
signal \N__11680\ : std_logic;
signal \N__11675\ : std_logic;
signal \N__11672\ : std_logic;
signal \N__11671\ : std_logic;
signal \N__11670\ : std_logic;
signal \N__11669\ : std_logic;
signal \N__11662\ : std_logic;
signal \N__11659\ : std_logic;
signal \N__11654\ : std_logic;
signal \N__11653\ : std_logic;
signal \N__11650\ : std_logic;
signal \N__11647\ : std_logic;
signal \N__11644\ : std_logic;
signal \N__11639\ : std_logic;
signal \N__11636\ : std_logic;
signal \N__11635\ : std_logic;
signal \N__11632\ : std_logic;
signal \N__11629\ : std_logic;
signal \N__11626\ : std_logic;
signal \N__11623\ : std_logic;
signal \N__11620\ : std_logic;
signal \N__11617\ : std_logic;
signal \N__11614\ : std_logic;
signal \N__11609\ : std_logic;
signal \N__11606\ : std_logic;
signal \N__11603\ : std_logic;
signal \N__11600\ : std_logic;
signal \N__11597\ : std_logic;
signal \N__11594\ : std_logic;
signal \N__11591\ : std_logic;
signal \N__11590\ : std_logic;
signal \N__11589\ : std_logic;
signal \N__11588\ : std_logic;
signal \N__11583\ : std_logic;
signal \N__11578\ : std_logic;
signal \N__11573\ : std_logic;
signal \N__11572\ : std_logic;
signal \N__11571\ : std_logic;
signal \N__11570\ : std_logic;
signal \N__11565\ : std_logic;
signal \N__11560\ : std_logic;
signal \N__11555\ : std_logic;
signal \N__11552\ : std_logic;
signal \N__11551\ : std_logic;
signal \N__11550\ : std_logic;
signal \N__11547\ : std_logic;
signal \N__11540\ : std_logic;
signal \N__11537\ : std_logic;
signal \N__11536\ : std_logic;
signal \N__11533\ : std_logic;
signal \N__11530\ : std_logic;
signal \N__11525\ : std_logic;
signal \N__11522\ : std_logic;
signal \N__11519\ : std_logic;
signal \N__11516\ : std_logic;
signal \N__11513\ : std_logic;
signal \N__11512\ : std_logic;
signal \N__11511\ : std_logic;
signal \N__11510\ : std_logic;
signal \N__11507\ : std_logic;
signal \N__11506\ : std_logic;
signal \N__11503\ : std_logic;
signal \N__11500\ : std_logic;
signal \N__11497\ : std_logic;
signal \N__11494\ : std_logic;
signal \N__11491\ : std_logic;
signal \N__11488\ : std_logic;
signal \N__11485\ : std_logic;
signal \N__11474\ : std_logic;
signal \N__11473\ : std_logic;
signal \N__11472\ : std_logic;
signal \N__11471\ : std_logic;
signal \N__11468\ : std_logic;
signal \N__11465\ : std_logic;
signal \N__11462\ : std_logic;
signal \N__11459\ : std_logic;
signal \N__11458\ : std_logic;
signal \N__11455\ : std_logic;
signal \N__11452\ : std_logic;
signal \N__11449\ : std_logic;
signal \N__11446\ : std_logic;
signal \N__11443\ : std_logic;
signal \N__11438\ : std_logic;
signal \N__11429\ : std_logic;
signal \N__11428\ : std_logic;
signal \N__11427\ : std_logic;
signal \N__11426\ : std_logic;
signal \N__11423\ : std_logic;
signal \N__11420\ : std_logic;
signal \N__11419\ : std_logic;
signal \N__11416\ : std_logic;
signal \N__11413\ : std_logic;
signal \N__11410\ : std_logic;
signal \N__11407\ : std_logic;
signal \N__11404\ : std_logic;
signal \N__11401\ : std_logic;
signal \N__11390\ : std_logic;
signal \N__11389\ : std_logic;
signal \N__11388\ : std_logic;
signal \N__11387\ : std_logic;
signal \N__11386\ : std_logic;
signal \N__11383\ : std_logic;
signal \N__11380\ : std_logic;
signal \N__11377\ : std_logic;
signal \N__11374\ : std_logic;
signal \N__11371\ : std_logic;
signal \N__11368\ : std_logic;
signal \N__11365\ : std_logic;
signal \N__11362\ : std_logic;
signal \N__11359\ : std_logic;
signal \N__11356\ : std_logic;
signal \N__11345\ : std_logic;
signal \N__11344\ : std_logic;
signal \N__11341\ : std_logic;
signal \N__11338\ : std_logic;
signal \N__11337\ : std_logic;
signal \N__11334\ : std_logic;
signal \N__11331\ : std_logic;
signal \N__11328\ : std_logic;
signal \N__11327\ : std_logic;
signal \N__11326\ : std_logic;
signal \N__11319\ : std_logic;
signal \N__11314\ : std_logic;
signal \N__11309\ : std_logic;
signal \N__11308\ : std_logic;
signal \N__11305\ : std_logic;
signal \N__11304\ : std_logic;
signal \N__11303\ : std_logic;
signal \N__11300\ : std_logic;
signal \N__11297\ : std_logic;
signal \N__11294\ : std_logic;
signal \N__11293\ : std_logic;
signal \N__11290\ : std_logic;
signal \N__11287\ : std_logic;
signal \N__11284\ : std_logic;
signal \N__11281\ : std_logic;
signal \N__11278\ : std_logic;
signal \N__11267\ : std_logic;
signal \N__11264\ : std_logic;
signal \N__11263\ : std_logic;
signal \N__11262\ : std_logic;
signal \N__11259\ : std_logic;
signal \N__11256\ : std_logic;
signal \N__11253\ : std_logic;
signal \N__11250\ : std_logic;
signal \N__11247\ : std_logic;
signal \N__11244\ : std_logic;
signal \N__11243\ : std_logic;
signal \N__11242\ : std_logic;
signal \N__11235\ : std_logic;
signal \N__11232\ : std_logic;
signal \N__11229\ : std_logic;
signal \N__11222\ : std_logic;
signal \N__11221\ : std_logic;
signal \N__11218\ : std_logic;
signal \N__11217\ : std_logic;
signal \N__11214\ : std_logic;
signal \N__11213\ : std_logic;
signal \N__11210\ : std_logic;
signal \N__11207\ : std_logic;
signal \N__11204\ : std_logic;
signal \N__11203\ : std_logic;
signal \N__11200\ : std_logic;
signal \N__11197\ : std_logic;
signal \N__11194\ : std_logic;
signal \N__11191\ : std_logic;
signal \N__11188\ : std_logic;
signal \N__11185\ : std_logic;
signal \N__11178\ : std_logic;
signal \N__11175\ : std_logic;
signal \N__11168\ : std_logic;
signal \N__11167\ : std_logic;
signal \N__11164\ : std_logic;
signal \N__11163\ : std_logic;
signal \N__11160\ : std_logic;
signal \N__11157\ : std_logic;
signal \N__11156\ : std_logic;
signal \N__11155\ : std_logic;
signal \N__11152\ : std_logic;
signal \N__11149\ : std_logic;
signal \N__11146\ : std_logic;
signal \N__11143\ : std_logic;
signal \N__11140\ : std_logic;
signal \N__11129\ : std_logic;
signal \N__11126\ : std_logic;
signal \N__11125\ : std_logic;
signal \N__11122\ : std_logic;
signal \N__11121\ : std_logic;
signal \N__11118\ : std_logic;
signal \N__11115\ : std_logic;
signal \N__11112\ : std_logic;
signal \N__11109\ : std_logic;
signal \N__11102\ : std_logic;
signal \N__11099\ : std_logic;
signal \N__11098\ : std_logic;
signal \N__11095\ : std_logic;
signal \N__11094\ : std_logic;
signal \N__11091\ : std_logic;
signal \N__11088\ : std_logic;
signal \N__11085\ : std_logic;
signal \N__11082\ : std_logic;
signal \N__11075\ : std_logic;
signal \N__11074\ : std_logic;
signal \N__11071\ : std_logic;
signal \N__11070\ : std_logic;
signal \N__11067\ : std_logic;
signal \N__11064\ : std_logic;
signal \N__11061\ : std_logic;
signal \N__11060\ : std_logic;
signal \N__11057\ : std_logic;
signal \N__11056\ : std_logic;
signal \N__11051\ : std_logic;
signal \N__11048\ : std_logic;
signal \N__11045\ : std_logic;
signal \N__11042\ : std_logic;
signal \N__11033\ : std_logic;
signal \N__11032\ : std_logic;
signal \N__11029\ : std_logic;
signal \N__11026\ : std_logic;
signal \N__11023\ : std_logic;
signal \N__11022\ : std_logic;
signal \N__11021\ : std_logic;
signal \N__11018\ : std_logic;
signal \N__11015\ : std_logic;
signal \N__11012\ : std_logic;
signal \N__11011\ : std_logic;
signal \N__11008\ : std_logic;
signal \N__11003\ : std_logic;
signal \N__11000\ : std_logic;
signal \N__10997\ : std_logic;
signal \N__10988\ : std_logic;
signal \N__10985\ : std_logic;
signal \N__10984\ : std_logic;
signal \N__10981\ : std_logic;
signal \N__10980\ : std_logic;
signal \N__10977\ : std_logic;
signal \N__10974\ : std_logic;
signal \N__10971\ : std_logic;
signal \N__10968\ : std_logic;
signal \N__10963\ : std_logic;
signal \N__10958\ : std_logic;
signal \N__10955\ : std_logic;
signal \N__10954\ : std_logic;
signal \N__10951\ : std_logic;
signal \N__10950\ : std_logic;
signal \N__10947\ : std_logic;
signal \N__10946\ : std_logic;
signal \N__10943\ : std_logic;
signal \N__10942\ : std_logic;
signal \N__10939\ : std_logic;
signal \N__10936\ : std_logic;
signal \N__10933\ : std_logic;
signal \N__10930\ : std_logic;
signal \N__10927\ : std_logic;
signal \N__10916\ : std_logic;
signal \N__10913\ : std_logic;
signal \N__10910\ : std_logic;
signal \N__10909\ : std_logic;
signal \N__10906\ : std_logic;
signal \N__10905\ : std_logic;
signal \N__10902\ : std_logic;
signal \N__10899\ : std_logic;
signal \N__10896\ : std_logic;
signal \N__10893\ : std_logic;
signal \N__10886\ : std_logic;
signal \N__10885\ : std_logic;
signal \N__10884\ : std_logic;
signal \N__10881\ : std_logic;
signal \N__10878\ : std_logic;
signal \N__10875\ : std_logic;
signal \N__10872\ : std_logic;
signal \N__10871\ : std_logic;
signal \N__10870\ : std_logic;
signal \N__10865\ : std_logic;
signal \N__10862\ : std_logic;
signal \N__10859\ : std_logic;
signal \N__10856\ : std_logic;
signal \N__10847\ : std_logic;
signal \N__10846\ : std_logic;
signal \N__10845\ : std_logic;
signal \N__10842\ : std_logic;
signal \N__10839\ : std_logic;
signal \N__10836\ : std_logic;
signal \N__10833\ : std_logic;
signal \N__10830\ : std_logic;
signal \N__10829\ : std_logic;
signal \N__10828\ : std_logic;
signal \N__10825\ : std_logic;
signal \N__10822\ : std_logic;
signal \N__10819\ : std_logic;
signal \N__10816\ : std_logic;
signal \N__10813\ : std_logic;
signal \N__10802\ : std_logic;
signal \N__10801\ : std_logic;
signal \N__10798\ : std_logic;
signal \N__10795\ : std_logic;
signal \N__10794\ : std_logic;
signal \N__10793\ : std_logic;
signal \N__10790\ : std_logic;
signal \N__10787\ : std_logic;
signal \N__10784\ : std_logic;
signal \N__10783\ : std_logic;
signal \N__10780\ : std_logic;
signal \N__10777\ : std_logic;
signal \N__10774\ : std_logic;
signal \N__10771\ : std_logic;
signal \N__10768\ : std_logic;
signal \N__10757\ : std_logic;
signal \N__10756\ : std_logic;
signal \N__10753\ : std_logic;
signal \N__10752\ : std_logic;
signal \N__10749\ : std_logic;
signal \N__10746\ : std_logic;
signal \N__10743\ : std_logic;
signal \N__10740\ : std_logic;
signal \N__10735\ : std_logic;
signal \N__10730\ : std_logic;
signal \N__10727\ : std_logic;
signal \N__10724\ : std_logic;
signal \N__10721\ : std_logic;
signal \N__10718\ : std_logic;
signal \N__10715\ : std_logic;
signal \N__10712\ : std_logic;
signal \N__10709\ : std_logic;
signal \N__10706\ : std_logic;
signal \N__10705\ : std_logic;
signal \N__10702\ : std_logic;
signal \N__10701\ : std_logic;
signal \N__10700\ : std_logic;
signal \N__10697\ : std_logic;
signal \N__10696\ : std_logic;
signal \N__10695\ : std_logic;
signal \N__10692\ : std_logic;
signal \N__10689\ : std_logic;
signal \N__10688\ : std_logic;
signal \N__10685\ : std_logic;
signal \N__10682\ : std_logic;
signal \N__10681\ : std_logic;
signal \N__10680\ : std_logic;
signal \N__10679\ : std_logic;
signal \N__10678\ : std_logic;
signal \N__10673\ : std_logic;
signal \N__10668\ : std_logic;
signal \N__10665\ : std_logic;
signal \N__10662\ : std_logic;
signal \N__10659\ : std_logic;
signal \N__10654\ : std_logic;
signal \N__10649\ : std_logic;
signal \N__10646\ : std_logic;
signal \N__10641\ : std_logic;
signal \N__10628\ : std_logic;
signal \N__10625\ : std_logic;
signal \N__10622\ : std_logic;
signal \N__10619\ : std_logic;
signal \N__10616\ : std_logic;
signal \N__10613\ : std_logic;
signal \N__10612\ : std_logic;
signal \N__10611\ : std_logic;
signal \N__10610\ : std_logic;
signal \N__10607\ : std_logic;
signal \N__10604\ : std_logic;
signal \N__10601\ : std_logic;
signal \N__10598\ : std_logic;
signal \N__10589\ : std_logic;
signal \N__10586\ : std_logic;
signal \N__10583\ : std_logic;
signal \N__10580\ : std_logic;
signal \N__10577\ : std_logic;
signal \N__10574\ : std_logic;
signal \N__10571\ : std_logic;
signal \N__10570\ : std_logic;
signal \N__10569\ : std_logic;
signal \N__10568\ : std_logic;
signal \N__10567\ : std_logic;
signal \N__10564\ : std_logic;
signal \N__10563\ : std_logic;
signal \N__10562\ : std_logic;
signal \N__10559\ : std_logic;
signal \N__10558\ : std_logic;
signal \N__10557\ : std_logic;
signal \N__10554\ : std_logic;
signal \N__10553\ : std_logic;
signal \N__10548\ : std_logic;
signal \N__10547\ : std_logic;
signal \N__10546\ : std_logic;
signal \N__10545\ : std_logic;
signal \N__10544\ : std_logic;
signal \N__10543\ : std_logic;
signal \N__10542\ : std_logic;
signal \N__10541\ : std_logic;
signal \N__10540\ : std_logic;
signal \N__10537\ : std_logic;
signal \N__10534\ : std_logic;
signal \N__10531\ : std_logic;
signal \N__10528\ : std_logic;
signal \N__10519\ : std_logic;
signal \N__10518\ : std_logic;
signal \N__10517\ : std_logic;
signal \N__10516\ : std_logic;
signal \N__10515\ : std_logic;
signal \N__10514\ : std_logic;
signal \N__10513\ : std_logic;
signal \N__10512\ : std_logic;
signal \N__10511\ : std_logic;
signal \N__10510\ : std_logic;
signal \N__10507\ : std_logic;
signal \N__10494\ : std_logic;
signal \N__10489\ : std_logic;
signal \N__10482\ : std_logic;
signal \N__10477\ : std_logic;
signal \N__10472\ : std_logic;
signal \N__10467\ : std_logic;
signal \N__10456\ : std_logic;
signal \N__10451\ : std_logic;
signal \N__10444\ : std_logic;
signal \N__10433\ : std_logic;
signal \N__10432\ : std_logic;
signal \N__10431\ : std_logic;
signal \N__10430\ : std_logic;
signal \N__10429\ : std_logic;
signal \N__10428\ : std_logic;
signal \N__10427\ : std_logic;
signal \N__10426\ : std_logic;
signal \N__10425\ : std_logic;
signal \N__10420\ : std_logic;
signal \N__10419\ : std_logic;
signal \N__10414\ : std_logic;
signal \N__10411\ : std_logic;
signal \N__10406\ : std_logic;
signal \N__10401\ : std_logic;
signal \N__10398\ : std_logic;
signal \N__10395\ : std_logic;
signal \N__10392\ : std_logic;
signal \N__10383\ : std_logic;
signal \N__10376\ : std_logic;
signal \N__10373\ : std_logic;
signal \N__10370\ : std_logic;
signal \N__10367\ : std_logic;
signal \N__10364\ : std_logic;
signal \N__10361\ : std_logic;
signal \N__10358\ : std_logic;
signal \N__10355\ : std_logic;
signal \N__10352\ : std_logic;
signal \N__10351\ : std_logic;
signal \N__10350\ : std_logic;
signal \N__10349\ : std_logic;
signal \N__10346\ : std_logic;
signal \N__10343\ : std_logic;
signal \N__10340\ : std_logic;
signal \N__10337\ : std_logic;
signal \N__10334\ : std_logic;
signal \N__10333\ : std_logic;
signal \N__10330\ : std_logic;
signal \N__10327\ : std_logic;
signal \N__10324\ : std_logic;
signal \N__10321\ : std_logic;
signal \N__10318\ : std_logic;
signal \N__10315\ : std_logic;
signal \N__10312\ : std_logic;
signal \N__10307\ : std_logic;
signal \N__10302\ : std_logic;
signal \N__10295\ : std_logic;
signal \N__10294\ : std_logic;
signal \N__10291\ : std_logic;
signal \N__10288\ : std_logic;
signal \N__10287\ : std_logic;
signal \N__10286\ : std_logic;
signal \N__10283\ : std_logic;
signal \N__10282\ : std_logic;
signal \N__10279\ : std_logic;
signal \N__10276\ : std_logic;
signal \N__10273\ : std_logic;
signal \N__10270\ : std_logic;
signal \N__10267\ : std_logic;
signal \N__10264\ : std_logic;
signal \N__10259\ : std_logic;
signal \N__10250\ : std_logic;
signal \N__10247\ : std_logic;
signal \N__10246\ : std_logic;
signal \N__10243\ : std_logic;
signal \N__10242\ : std_logic;
signal \N__10239\ : std_logic;
signal \N__10236\ : std_logic;
signal \N__10233\ : std_logic;
signal \N__10230\ : std_logic;
signal \N__10223\ : std_logic;
signal \N__10220\ : std_logic;
signal \N__10217\ : std_logic;
signal \N__10214\ : std_logic;
signal \N__10211\ : std_logic;
signal \N__10210\ : std_logic;
signal \N__10209\ : std_logic;
signal \N__10208\ : std_logic;
signal \N__10207\ : std_logic;
signal \N__10206\ : std_logic;
signal \N__10203\ : std_logic;
signal \N__10198\ : std_logic;
signal \N__10191\ : std_logic;
signal \N__10184\ : std_logic;
signal \N__10183\ : std_logic;
signal \N__10182\ : std_logic;
signal \N__10175\ : std_logic;
signal \N__10172\ : std_logic;
signal \N__10171\ : std_logic;
signal \N__10168\ : std_logic;
signal \N__10165\ : std_logic;
signal \N__10164\ : std_logic;
signal \N__10161\ : std_logic;
signal \N__10158\ : std_logic;
signal \N__10157\ : std_logic;
signal \N__10154\ : std_logic;
signal \N__10151\ : std_logic;
signal \N__10148\ : std_logic;
signal \N__10145\ : std_logic;
signal \N__10144\ : std_logic;
signal \N__10143\ : std_logic;
signal \N__10140\ : std_logic;
signal \N__10137\ : std_logic;
signal \N__10134\ : std_logic;
signal \N__10131\ : std_logic;
signal \N__10126\ : std_logic;
signal \N__10123\ : std_logic;
signal \N__10120\ : std_logic;
signal \N__10117\ : std_logic;
signal \N__10106\ : std_logic;
signal \N__10103\ : std_logic;
signal \N__10100\ : std_logic;
signal \N__10097\ : std_logic;
signal \N__10094\ : std_logic;
signal \N__10091\ : std_logic;
signal \N__10088\ : std_logic;
signal \N__10085\ : std_logic;
signal \N__10082\ : std_logic;
signal \N__10079\ : std_logic;
signal \N__10076\ : std_logic;
signal \N__10073\ : std_logic;
signal \N__10070\ : std_logic;
signal \N__10067\ : std_logic;
signal \N__10064\ : std_logic;
signal \N__10061\ : std_logic;
signal \N__10058\ : std_logic;
signal \N__10055\ : std_logic;
signal \N__10052\ : std_logic;
signal \N__10049\ : std_logic;
signal \N__10046\ : std_logic;
signal \N__10043\ : std_logic;
signal \N__10040\ : std_logic;
signal \N__10037\ : std_logic;
signal \N__10034\ : std_logic;
signal \N__10031\ : std_logic;
signal \N__10028\ : std_logic;
signal \N__10027\ : std_logic;
signal \N__10024\ : std_logic;
signal \N__10023\ : std_logic;
signal \N__10020\ : std_logic;
signal \N__10017\ : std_logic;
signal \N__10014\ : std_logic;
signal \N__10011\ : std_logic;
signal \N__10008\ : std_logic;
signal \N__10005\ : std_logic;
signal \N__10002\ : std_logic;
signal \N__9995\ : std_logic;
signal \N__9992\ : std_logic;
signal \N__9989\ : std_logic;
signal \N__9986\ : std_logic;
signal \N__9983\ : std_logic;
signal \N__9980\ : std_logic;
signal \N__9977\ : std_logic;
signal \N__9974\ : std_logic;
signal \N__9971\ : std_logic;
signal \N__9970\ : std_logic;
signal \N__9967\ : std_logic;
signal \N__9964\ : std_logic;
signal \N__9959\ : std_logic;
signal \N__9956\ : std_logic;
signal \N__9953\ : std_logic;
signal \N__9950\ : std_logic;
signal \N__9947\ : std_logic;
signal \N__9946\ : std_logic;
signal \N__9943\ : std_logic;
signal \N__9940\ : std_logic;
signal \N__9935\ : std_logic;
signal \N__9932\ : std_logic;
signal \N__9929\ : std_logic;
signal \N__9926\ : std_logic;
signal \N__9923\ : std_logic;
signal \N__9920\ : std_logic;
signal \N__9917\ : std_logic;
signal \N__9914\ : std_logic;
signal \N__9911\ : std_logic;
signal \N__9908\ : std_logic;
signal \N__9905\ : std_logic;
signal \N__9902\ : std_logic;
signal \N__9899\ : std_logic;
signal \N__9896\ : std_logic;
signal \N__9893\ : std_logic;
signal \N__9890\ : std_logic;
signal \N__9887\ : std_logic;
signal \N__9884\ : std_logic;
signal \N__9881\ : std_logic;
signal \N__9878\ : std_logic;
signal \N__9875\ : std_logic;
signal \N__9872\ : std_logic;
signal \N__9871\ : std_logic;
signal \N__9868\ : std_logic;
signal \N__9865\ : std_logic;
signal \N__9862\ : std_logic;
signal \N__9859\ : std_logic;
signal \N__9854\ : std_logic;
signal \N__9853\ : std_logic;
signal \N__9850\ : std_logic;
signal \N__9847\ : std_logic;
signal \N__9844\ : std_logic;
signal \N__9841\ : std_logic;
signal \N__9836\ : std_logic;
signal \N__9835\ : std_logic;
signal \N__9832\ : std_logic;
signal \N__9829\ : std_logic;
signal \N__9826\ : std_logic;
signal \N__9823\ : std_logic;
signal \N__9818\ : std_logic;
signal \N__9817\ : std_logic;
signal \N__9814\ : std_logic;
signal \N__9811\ : std_logic;
signal \N__9808\ : std_logic;
signal \N__9805\ : std_logic;
signal \N__9802\ : std_logic;
signal \N__9797\ : std_logic;
signal \N__9796\ : std_logic;
signal \N__9793\ : std_logic;
signal \N__9790\ : std_logic;
signal \N__9787\ : std_logic;
signal \N__9784\ : std_logic;
signal \N__9781\ : std_logic;
signal \N__9776\ : std_logic;
signal \N__9775\ : std_logic;
signal \N__9772\ : std_logic;
signal \N__9769\ : std_logic;
signal \N__9766\ : std_logic;
signal \N__9763\ : std_logic;
signal \N__9760\ : std_logic;
signal \N__9757\ : std_logic;
signal \N__9752\ : std_logic;
signal \N__9751\ : std_logic;
signal \N__9748\ : std_logic;
signal \N__9745\ : std_logic;
signal \N__9742\ : std_logic;
signal \N__9739\ : std_logic;
signal \N__9736\ : std_logic;
signal \N__9731\ : std_logic;
signal \N__9728\ : std_logic;
signal \N__9727\ : std_logic;
signal \N__9724\ : std_logic;
signal \N__9721\ : std_logic;
signal \N__9716\ : std_logic;
signal \N__9713\ : std_logic;
signal \N__9710\ : std_logic;
signal \N__9707\ : std_logic;
signal \N__9704\ : std_logic;
signal \N__9701\ : std_logic;
signal \N__9698\ : std_logic;
signal \N__9695\ : std_logic;
signal \N__9692\ : std_logic;
signal \N__9689\ : std_logic;
signal \N__9686\ : std_logic;
signal \N__9683\ : std_logic;
signal \N__9680\ : std_logic;
signal \N__9677\ : std_logic;
signal \N__9674\ : std_logic;
signal \N__9671\ : std_logic;
signal \N__9670\ : std_logic;
signal \N__9669\ : std_logic;
signal \N__9668\ : std_logic;
signal \N__9663\ : std_logic;
signal \N__9660\ : std_logic;
signal \N__9657\ : std_logic;
signal \N__9650\ : std_logic;
signal \N__9647\ : std_logic;
signal \N__9644\ : std_logic;
signal \N__9641\ : std_logic;
signal \N__9638\ : std_logic;
signal \N__9635\ : std_logic;
signal \N__9632\ : std_logic;
signal \N__9629\ : std_logic;
signal \N__9628\ : std_logic;
signal \N__9625\ : std_logic;
signal \N__9622\ : std_logic;
signal \N__9619\ : std_logic;
signal \N__9616\ : std_logic;
signal \N__9611\ : std_logic;
signal \N__9608\ : std_logic;
signal \N__9605\ : std_logic;
signal \N__9604\ : std_logic;
signal \N__9601\ : std_logic;
signal \N__9598\ : std_logic;
signal \N__9593\ : std_logic;
signal \N__9590\ : std_logic;
signal \N__9589\ : std_logic;
signal \N__9586\ : std_logic;
signal \N__9583\ : std_logic;
signal \N__9580\ : std_logic;
signal \N__9575\ : std_logic;
signal \N__9572\ : std_logic;
signal \N__9569\ : std_logic;
signal \N__9566\ : std_logic;
signal \N__9563\ : std_logic;
signal \N__9560\ : std_logic;
signal \N__9557\ : std_logic;
signal \N__9554\ : std_logic;
signal \N__9551\ : std_logic;
signal \N__9548\ : std_logic;
signal \N__9545\ : std_logic;
signal \N__9542\ : std_logic;
signal \N__9539\ : std_logic;
signal \N__9536\ : std_logic;
signal \N__9533\ : std_logic;
signal \N__9530\ : std_logic;
signal \N__9527\ : std_logic;
signal \N__9526\ : std_logic;
signal \N__9523\ : std_logic;
signal \N__9520\ : std_logic;
signal \N__9517\ : std_logic;
signal \N__9512\ : std_logic;
signal \N__9511\ : std_logic;
signal \N__9510\ : std_logic;
signal \N__9509\ : std_logic;
signal \N__9506\ : std_logic;
signal \N__9499\ : std_logic;
signal \N__9494\ : std_logic;
signal \N__9491\ : std_logic;
signal \N__9488\ : std_logic;
signal \N__9485\ : std_logic;
signal \N__9484\ : std_logic;
signal \N__9483\ : std_logic;
signal \N__9482\ : std_logic;
signal \N__9479\ : std_logic;
signal \N__9472\ : std_logic;
signal \N__9467\ : std_logic;
signal \N__9464\ : std_logic;
signal \N__9461\ : std_logic;
signal \N__9458\ : std_logic;
signal \N__9455\ : std_logic;
signal \N__9454\ : std_logic;
signal \N__9453\ : std_logic;
signal \N__9452\ : std_logic;
signal \N__9447\ : std_logic;
signal \N__9444\ : std_logic;
signal \N__9441\ : std_logic;
signal \N__9436\ : std_logic;
signal \N__9431\ : std_logic;
signal \N__9428\ : std_logic;
signal \N__9427\ : std_logic;
signal \N__9426\ : std_logic;
signal \N__9425\ : std_logic;
signal \N__9422\ : std_logic;
signal \N__9419\ : std_logic;
signal \N__9414\ : std_logic;
signal \N__9407\ : std_logic;
signal \N__9404\ : std_logic;
signal \N__9401\ : std_logic;
signal \N__9398\ : std_logic;
signal \N__9397\ : std_logic;
signal \N__9396\ : std_logic;
signal \N__9393\ : std_logic;
signal \N__9392\ : std_logic;
signal \N__9389\ : std_logic;
signal \N__9386\ : std_logic;
signal \N__9383\ : std_logic;
signal \N__9380\ : std_logic;
signal \N__9371\ : std_logic;
signal \N__9368\ : std_logic;
signal \N__9365\ : std_logic;
signal \N__9362\ : std_logic;
signal \N__9359\ : std_logic;
signal \N__9356\ : std_logic;
signal \N__9353\ : std_logic;
signal \N__9350\ : std_logic;
signal \N__9347\ : std_logic;
signal \N__9344\ : std_logic;
signal \N__9341\ : std_logic;
signal \N__9340\ : std_logic;
signal \N__9339\ : std_logic;
signal \N__9338\ : std_logic;
signal \N__9337\ : std_logic;
signal \N__9336\ : std_logic;
signal \N__9323\ : std_logic;
signal \N__9320\ : std_logic;
signal \N__9317\ : std_logic;
signal \N__9314\ : std_logic;
signal \N__9311\ : std_logic;
signal \N__9310\ : std_logic;
signal \N__9309\ : std_logic;
signal \N__9308\ : std_logic;
signal \N__9305\ : std_logic;
signal \N__9302\ : std_logic;
signal \N__9297\ : std_logic;
signal \N__9290\ : std_logic;
signal \N__9287\ : std_logic;
signal \N__9284\ : std_logic;
signal \N__9283\ : std_logic;
signal \N__9282\ : std_logic;
signal \N__9281\ : std_logic;
signal \N__9278\ : std_logic;
signal \N__9271\ : std_logic;
signal \N__9266\ : std_logic;
signal \N__9263\ : std_logic;
signal \N__9262\ : std_logic;
signal \N__9259\ : std_logic;
signal \N__9258\ : std_logic;
signal \N__9257\ : std_logic;
signal \N__9252\ : std_logic;
signal \N__9249\ : std_logic;
signal \N__9246\ : std_logic;
signal \N__9239\ : std_logic;
signal \N__9236\ : std_logic;
signal \N__9235\ : std_logic;
signal \N__9234\ : std_logic;
signal \N__9233\ : std_logic;
signal \N__9230\ : std_logic;
signal \N__9223\ : std_logic;
signal \N__9218\ : std_logic;
signal \N__9215\ : std_logic;
signal \N__9212\ : std_logic;
signal \N__9209\ : std_logic;
signal \N__9208\ : std_logic;
signal \N__9207\ : std_logic;
signal \N__9206\ : std_logic;
signal \N__9203\ : std_logic;
signal \N__9196\ : std_logic;
signal \N__9191\ : std_logic;
signal \N__9188\ : std_logic;
signal \N__9187\ : std_logic;
signal \N__9186\ : std_logic;
signal \N__9185\ : std_logic;
signal \N__9182\ : std_logic;
signal \N__9179\ : std_logic;
signal \N__9174\ : std_logic;
signal \N__9167\ : std_logic;
signal \N__9164\ : std_logic;
signal \N__9161\ : std_logic;
signal \N__9158\ : std_logic;
signal \N__9157\ : std_logic;
signal \N__9156\ : std_logic;
signal \N__9155\ : std_logic;
signal \N__9152\ : std_logic;
signal \N__9149\ : std_logic;
signal \N__9144\ : std_logic;
signal \N__9137\ : std_logic;
signal \N__9134\ : std_logic;
signal \N__9131\ : std_logic;
signal \N__9128\ : std_logic;
signal \N__9125\ : std_logic;
signal \N__9124\ : std_logic;
signal \N__9119\ : std_logic;
signal \N__9116\ : std_logic;
signal \N__9113\ : std_logic;
signal \N__9110\ : std_logic;
signal \N__9107\ : std_logic;
signal \N__9104\ : std_logic;
signal \N__9101\ : std_logic;
signal \N__9098\ : std_logic;
signal \N__9095\ : std_logic;
signal \N__9092\ : std_logic;
signal \N__9089\ : std_logic;
signal \N__9086\ : std_logic;
signal \N__9083\ : std_logic;
signal \N__9080\ : std_logic;
signal \N__9077\ : std_logic;
signal \N__9074\ : std_logic;
signal \N__9071\ : std_logic;
signal \N__9068\ : std_logic;
signal \N__9065\ : std_logic;
signal \N__9062\ : std_logic;
signal \N__9059\ : std_logic;
signal \N__9056\ : std_logic;
signal \N__9053\ : std_logic;
signal \N__9050\ : std_logic;
signal \N__9047\ : std_logic;
signal \N__9044\ : std_logic;
signal \N__9041\ : std_logic;
signal \N__9038\ : std_logic;
signal \N__9035\ : std_logic;
signal \N__9032\ : std_logic;
signal \N__9029\ : std_logic;
signal \N__9026\ : std_logic;
signal \N__9023\ : std_logic;
signal \N__9020\ : std_logic;
signal \N__9017\ : std_logic;
signal \N__9014\ : std_logic;
signal \N__9011\ : std_logic;
signal \N__9008\ : std_logic;
signal \N__9005\ : std_logic;
signal \N__9002\ : std_logic;
signal \N__8999\ : std_logic;
signal \N__8996\ : std_logic;
signal \N__8993\ : std_logic;
signal \N__8990\ : std_logic;
signal \N__8987\ : std_logic;
signal \N__8984\ : std_logic;
signal \N__8981\ : std_logic;
signal \N__8978\ : std_logic;
signal \N__8975\ : std_logic;
signal \N__8972\ : std_logic;
signal \N__8969\ : std_logic;
signal \N__8966\ : std_logic;
signal \N__8963\ : std_logic;
signal \N__8960\ : std_logic;
signal \N__8959\ : std_logic;
signal \N__8956\ : std_logic;
signal \N__8953\ : std_logic;
signal \N__8948\ : std_logic;
signal \N__8945\ : std_logic;
signal \N__8942\ : std_logic;
signal \N__8939\ : std_logic;
signal \N__8936\ : std_logic;
signal \N__8933\ : std_logic;
signal \N__8930\ : std_logic;
signal \N__8927\ : std_logic;
signal \N__8924\ : std_logic;
signal \N__8921\ : std_logic;
signal \N__8918\ : std_logic;
signal \N__8915\ : std_logic;
signal \N__8912\ : std_logic;
signal \N__8909\ : std_logic;
signal \N__8906\ : std_logic;
signal \N__8903\ : std_logic;
signal \N__8900\ : std_logic;
signal \N__8897\ : std_logic;
signal \N__8894\ : std_logic;
signal \N__8891\ : std_logic;
signal \N__8888\ : std_logic;
signal \N__8885\ : std_logic;
signal \N__8884\ : std_logic;
signal \N__8883\ : std_logic;
signal \N__8882\ : std_logic;
signal \N__8881\ : std_logic;
signal \N__8880\ : std_logic;
signal \N__8879\ : std_logic;
signal \N__8878\ : std_logic;
signal \N__8873\ : std_logic;
signal \N__8860\ : std_logic;
signal \N__8855\ : std_logic;
signal \N__8852\ : std_logic;
signal \N__8849\ : std_logic;
signal \N__8846\ : std_logic;
signal \N__8843\ : std_logic;
signal \N__8840\ : std_logic;
signal \N__8837\ : std_logic;
signal \N__8834\ : std_logic;
signal \N__8831\ : std_logic;
signal \N__8828\ : std_logic;
signal \N__8825\ : std_logic;
signal \N__8822\ : std_logic;
signal \N__8819\ : std_logic;
signal \N__8816\ : std_logic;
signal \N__8813\ : std_logic;
signal \N__8810\ : std_logic;
signal \N__8807\ : std_logic;
signal \N__8804\ : std_logic;
signal \N__8801\ : std_logic;
signal \N__8798\ : std_logic;
signal \N__8795\ : std_logic;
signal \N__8792\ : std_logic;
signal \N__8789\ : std_logic;
signal \N__8786\ : std_logic;
signal \N__8783\ : std_logic;
signal \N__8780\ : std_logic;
signal \N__8777\ : std_logic;
signal \N__8774\ : std_logic;
signal \N__8771\ : std_logic;
signal \N__8768\ : std_logic;
signal \N__8765\ : std_logic;
signal \N__8762\ : std_logic;
signal \N__8759\ : std_logic;
signal \N__8756\ : std_logic;
signal \N__8753\ : std_logic;
signal \N__8750\ : std_logic;
signal \N__8747\ : std_logic;
signal \N__8744\ : std_logic;
signal \N__8741\ : std_logic;
signal \N__8738\ : std_logic;
signal \N__8735\ : std_logic;
signal \N__8732\ : std_logic;
signal \N__8729\ : std_logic;
signal \N__8726\ : std_logic;
signal \N__8723\ : std_logic;
signal \N__8720\ : std_logic;
signal \N__8717\ : std_logic;
signal \N__8714\ : std_logic;
signal \N__8711\ : std_logic;
signal \N__8708\ : std_logic;
signal \N__8705\ : std_logic;
signal \N__8702\ : std_logic;
signal \N__8699\ : std_logic;
signal \N__8696\ : std_logic;
signal \N__8693\ : std_logic;
signal \N__8690\ : std_logic;
signal \N__8687\ : std_logic;
signal \N__8684\ : std_logic;
signal \N__8681\ : std_logic;
signal \N__8678\ : std_logic;
signal \N__8675\ : std_logic;
signal \N__8672\ : std_logic;
signal \N__8669\ : std_logic;
signal \N__8666\ : std_logic;
signal \N__8663\ : std_logic;
signal \N__8662\ : std_logic;
signal \N__8659\ : std_logic;
signal \N__8656\ : std_logic;
signal \N__8653\ : std_logic;
signal \N__8648\ : std_logic;
signal \N__8647\ : std_logic;
signal \N__8644\ : std_logic;
signal \N__8641\ : std_logic;
signal \N__8636\ : std_logic;
signal \N__8635\ : std_logic;
signal \N__8632\ : std_logic;
signal \N__8629\ : std_logic;
signal \N__8624\ : std_logic;
signal \N__8623\ : std_logic;
signal \N__8620\ : std_logic;
signal \N__8617\ : std_logic;
signal \N__8612\ : std_logic;
signal \N__8609\ : std_logic;
signal \N__8606\ : std_logic;
signal \N__8603\ : std_logic;
signal \N__8600\ : std_logic;
signal \N__8597\ : std_logic;
signal \N__8594\ : std_logic;
signal \N__8591\ : std_logic;
signal \N__8588\ : std_logic;
signal \N__8585\ : std_logic;
signal \N__8582\ : std_logic;
signal \N__8579\ : std_logic;
signal \N__8576\ : std_logic;
signal \N__8573\ : std_logic;
signal \N__8570\ : std_logic;
signal \N__8567\ : std_logic;
signal \N__8564\ : std_logic;
signal \N__8561\ : std_logic;
signal \N__8558\ : std_logic;
signal \N__8555\ : std_logic;
signal \N__8552\ : std_logic;
signal \N__8549\ : std_logic;
signal \N__8546\ : std_logic;
signal \N__8543\ : std_logic;
signal \N__8542\ : std_logic;
signal \N__8539\ : std_logic;
signal \N__8536\ : std_logic;
signal \N__8535\ : std_logic;
signal \N__8534\ : std_logic;
signal \N__8533\ : std_logic;
signal \N__8526\ : std_logic;
signal \N__8521\ : std_logic;
signal \N__8516\ : std_logic;
signal \N__8513\ : std_logic;
signal \N__8512\ : std_logic;
signal \N__8511\ : std_logic;
signal \N__8510\ : std_logic;
signal \N__8509\ : std_logic;
signal \N__8508\ : std_logic;
signal \N__8505\ : std_logic;
signal \N__8496\ : std_logic;
signal \N__8493\ : std_logic;
signal \N__8486\ : std_logic;
signal \N__8483\ : std_logic;
signal \N__8480\ : std_logic;
signal \N__8477\ : std_logic;
signal \N__8474\ : std_logic;
signal \N__8471\ : std_logic;
signal \N__8468\ : std_logic;
signal \N__8465\ : std_logic;
signal \N__8462\ : std_logic;
signal \N__8461\ : std_logic;
signal \N__8460\ : std_logic;
signal \N__8457\ : std_logic;
signal \N__8452\ : std_logic;
signal \N__8447\ : std_logic;
signal \N__8446\ : std_logic;
signal \N__8445\ : std_logic;
signal \N__8444\ : std_logic;
signal \N__8441\ : std_logic;
signal \N__8436\ : std_logic;
signal \N__8433\ : std_logic;
signal \N__8426\ : std_logic;
signal \N__8425\ : std_logic;
signal \N__8424\ : std_logic;
signal \N__8423\ : std_logic;
signal \N__8420\ : std_logic;
signal \N__8415\ : std_logic;
signal \N__8414\ : std_logic;
signal \N__8413\ : std_logic;
signal \N__8412\ : std_logic;
signal \N__8411\ : std_logic;
signal \N__8408\ : std_logic;
signal \N__8403\ : std_logic;
signal \N__8394\ : std_logic;
signal \N__8387\ : std_logic;
signal \N__8386\ : std_logic;
signal \N__8383\ : std_logic;
signal \N__8380\ : std_logic;
signal \N__8379\ : std_logic;
signal \N__8378\ : std_logic;
signal \N__8373\ : std_logic;
signal \N__8368\ : std_logic;
signal \N__8363\ : std_logic;
signal \N__8362\ : std_logic;
signal \N__8359\ : std_logic;
signal \N__8356\ : std_logic;
signal \N__8355\ : std_logic;
signal \N__8354\ : std_logic;
signal \N__8353\ : std_logic;
signal \N__8352\ : std_logic;
signal \N__8351\ : std_logic;
signal \N__8350\ : std_logic;
signal \N__8341\ : std_logic;
signal \N__8338\ : std_logic;
signal \N__8331\ : std_logic;
signal \N__8328\ : std_logic;
signal \N__8321\ : std_logic;
signal \N__8318\ : std_logic;
signal \N__8315\ : std_logic;
signal \N__8312\ : std_logic;
signal \N__8309\ : std_logic;
signal \N__8306\ : std_logic;
signal \N__8303\ : std_logic;
signal \N__8300\ : std_logic;
signal \N__8297\ : std_logic;
signal \N__8294\ : std_logic;
signal \N__8291\ : std_logic;
signal \N__8288\ : std_logic;
signal \N__8285\ : std_logic;
signal \N__8282\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \b2v_inst.cuenta_pixel_RNO_0Z0Z_1\ : std_logic;
signal \b2v_inst.g0_10_a3_0_4\ : std_logic;
signal \b2v_inst.g0_10_a3_0_7_cascade_\ : std_logic;
signal \b2v_inst.g0_10_a3_0_5\ : std_logic;
signal \b2v_inst.g0_10_a3_5_cascade_\ : std_logic;
signal \b2v_inst.g0_10_a3_4\ : std_logic;
signal \b2v_inst.un1_cuenta_pixel_c6\ : std_logic;
signal \b2v_inst.un1_cuenta_pixel_c6_cascade_\ : std_logic;
signal \b2v_inst.cuenta_pixelZ0Z_7\ : std_logic;
signal \b2v_inst.cuenta_pixelZ0Z_2\ : std_logic;
signal \b2v_inst.N_6_i\ : std_logic;
signal \b2v_inst.g0_6_1_cascade_\ : std_logic;
signal \b2v_inst.N_4\ : std_logic;
signal \b2v_inst.un11_cuenta_pixel_6_cascade_\ : std_logic;
signal \b2v_inst.un11_cuenta_pixel_6\ : std_logic;
signal \b2v_inst.cuenta_pixel_RNI3FD32_0Z0Z_5\ : std_logic;
signal \b2v_inst.cuenta_pixelZ0Z_3\ : std_logic;
signal \b2v_inst.un1_cuenta_pixel_c3\ : std_logic;
signal \b2v_inst.cuenta_pixelZ0Z_4\ : std_logic;
signal \bfn_1_15_0_\ : std_logic;
signal \b2v_inst.eventos_cry_0\ : std_logic;
signal \b2v_inst.eventos_cry_1\ : std_logic;
signal \b2v_inst.eventos_cry_2\ : std_logic;
signal \b2v_inst.eventos_cry_3\ : std_logic;
signal \b2v_inst.eventos_cry_4\ : std_logic;
signal \b2v_inst.eventos_cry_5\ : std_logic;
signal \b2v_inst.eventos_cry_6\ : std_logic;
signal \b2v_inst.eventosZ0Z_3\ : std_logic;
signal \b2v_inst.eventosZ0Z_4\ : std_logic;
signal \b2v_inst.eventosZ0Z_0\ : std_logic;
signal \b2v_inst.eventosZ0Z_5\ : std_logic;
signal \b2v_inst.N_47_i\ : std_logic;
signal \b2v_inst.reg_ancho_1_i_0\ : std_logic;
signal \bfn_1_17_0_\ : std_logic;
signal \b2v_inst.reg_ancho_1_i_1\ : std_logic;
signal \b2v_inst.un3_valor_max1_cry_0\ : std_logic;
signal \b2v_inst.reg_ancho_1_i_2\ : std_logic;
signal \b2v_inst.un3_valor_max1_cry_1\ : std_logic;
signal \b2v_inst.reg_ancho_1_i_3\ : std_logic;
signal \b2v_inst.un3_valor_max1_cry_2\ : std_logic;
signal \b2v_inst.reg_ancho_1_i_4\ : std_logic;
signal \b2v_inst.un3_valor_max1_cry_3\ : std_logic;
signal \b2v_inst.reg_ancho_1_i_5\ : std_logic;
signal \b2v_inst.un3_valor_max1_cry_4\ : std_logic;
signal \b2v_inst.reg_ancho_1_i_6\ : std_logic;
signal \b2v_inst.un3_valor_max1_cry_5\ : std_logic;
signal \b2v_inst.reg_ancho_1_i_7\ : std_logic;
signal \b2v_inst.un3_valor_max1_cry_6\ : std_logic;
signal \b2v_inst.un3_valor_max1\ : std_logic;
signal \bfn_1_18_0_\ : std_logic;
signal \bfn_1_19_0_\ : std_logic;
signal \b2v_inst.valor_max_final5_3_cry_0\ : std_logic;
signal \b2v_inst.valor_max_final5_3_cry_1\ : std_logic;
signal \b2v_inst.valor_max_final5_3_cry_2\ : std_logic;
signal \b2v_inst.valor_max_final5_3_cry_3\ : std_logic;
signal \b2v_inst.valor_max_final5_3_cry_4\ : std_logic;
signal \b2v_inst.valor_max_final5_3_cry_5\ : std_logic;
signal \b2v_inst.valor_max_final5_3_cry_6\ : std_logic;
signal \b2v_inst.valor_max_final53\ : std_logic;
signal \bfn_1_20_0_\ : std_logic;
signal \b2v_inst.g0_10_1\ : std_logic;
signal \b2v_inst.g0_10_a3_7\ : std_logic;
signal \bfn_2_11_0_\ : std_logic;
signal \b2v_inst.un1_pix_count_anterior_0_data_tmp_0\ : std_logic;
signal \b2v_inst.un1_pix_count_anterior_0_data_tmp_1\ : std_logic;
signal \b2v_inst.un1_pix_count_anterior_0_data_tmp_2\ : std_logic;
signal \b2v_inst.un1_pix_count_anterior_0_data_tmp_3\ : std_logic;
signal \b2v_inst.un1_pix_count_anterior_0_data_tmp_4\ : std_logic;
signal \b2v_inst.un1_pix_count_anterior_0_data_tmp_5\ : std_logic;
signal \b2v_inst.un1_pix_count_anterior_0_N_2\ : std_logic;
signal \b2v_inst.un1_pix_count_anterior_0_I_15_c_RNOZ0\ : std_logic;
signal \b2v_inst.pix_count_anteriorZ0Z_4\ : std_logic;
signal \b2v_inst.pix_count_anteriorZ0Z_5\ : std_logic;
signal \b2v_inst.pix_count_anteriorZ0Z_1\ : std_logic;
signal \b2v_inst.un1_pix_count_anterior_0_I_1_c_RNOZ0\ : std_logic;
signal \b2v_inst.pix_count_anteriorZ0Z_0\ : std_logic;
signal \b2v_inst.pix_count_anteriorZ0Z_12\ : std_logic;
signal \b2v_inst.un1_pix_count_anterior_0_I_39_c_RNOZ0\ : std_logic;
signal \b2v_inst.un1_pix_count_anterior_0_I_21_c_RNOZ0\ : std_logic;
signal \b2v_inst.pix_count_anteriorZ0Z_6\ : std_logic;
signal \b2v_inst4.un1_pix_count_int_0_sqmuxa_8_cascade_\ : std_logic;
signal \b2v_inst.pix_count_anteriorZ0Z_7\ : std_logic;
signal \b2v_inst.pix_count_anteriorZ0Z_8\ : std_logic;
signal \b2v_inst.un1_pix_count_anterior_0_I_51_c_RNOZ0\ : std_logic;
signal \b2v_inst.pix_count_anteriorZ0Z_9\ : std_logic;
signal \b2v_inst.un1_state_17_0\ : std_logic;
signal \b2v_inst.ignorar_anchoZ0Z_1\ : std_logic;
signal \b2v_inst.data_a_escribir_RNO_3Z0Z_4_cascade_\ : std_logic;
signal \b2v_inst.data_a_escribir_RNO_3Z0Z_0_cascade_\ : std_logic;
signal \b2v_inst.un1_reg_anterior_iv_0_0_0_0\ : std_logic;
signal \b2v_inst.un1_m3_2_0\ : std_logic;
signal \b2v_inst.data_a_escribir_RNO_1Z0Z_0_cascade_\ : std_logic;
signal \b2v_inst.un1_reg_anterior_iv_0_0_1_1_3\ : std_logic;
signal \b2v_inst.N_315_cascade_\ : std_logic;
signal \b2v_inst.un1_reg_anterior_iv_0_0_1_3\ : std_logic;
signal \b2v_inst.un1_reg_anterior_iv_0_0_a2_6_0_1_cascade_\ : std_logic;
signal \b2v_inst.N_317\ : std_logic;
signal \b2v_inst.un1_reg_anterior_iv_0_0_a2_4_tz_1_2\ : std_logic;
signal \b2v_inst.eventosZ0Z_2\ : std_logic;
signal \b2v_inst.N_320_tz_cascade_\ : std_logic;
signal \b2v_inst.un1_m3_0_m3_ns_1_cascade_\ : std_logic;
signal \b2v_inst.N_318\ : std_logic;
signal \b2v_inst.data_a_escribir_RNO_0Z0Z_4\ : std_logic;
signal \b2v_inst.un1_reg_anterior_iv_0_0_0_4\ : std_logic;
signal \N_211_i\ : std_logic;
signal \N_219_i\ : std_logic;
signal \N_217_i\ : std_logic;
signal \N_215_i\ : std_logic;
signal \b2v_inst.state_ns_i_i_a2_4Z0Z_6\ : std_logic;
signal \b2v_inst.state_ns_i_i_a2_4Z0Z_6_cascade_\ : std_logic;
signal \b2v_inst.N_497_cascade_\ : std_logic;
signal \b2v_inst.N_361\ : std_logic;
signal \b2v_inst.state_ns_i_i_a2_5Z0Z_6\ : std_logic;
signal \b2v_inst.N_254_i\ : std_logic;
signal \b2v_inst.pix_count_anteriorZ0Z_2\ : std_logic;
signal \b2v_inst.un1_pix_count_anterior_0_I_27_c_RNOZ0\ : std_logic;
signal \b2v_inst.pix_count_anteriorZ0Z_3\ : std_logic;
signal \b2v_inst.pix_count_anteriorZ0Z_10\ : std_logic;
signal \b2v_inst.un1_pix_count_anterior_0_I_9_c_RNOZ0\ : std_logic;
signal \b2v_inst.pix_count_anteriorZ0Z_11\ : std_logic;
signal \b2v_inst.N_254_i_g\ : std_logic;
signal \SYNTHESIZED_WIRE_2_0\ : std_logic;
signal \b2v_inst4.pix_count_int_RNO_0Z0Z_0\ : std_logic;
signal \bfn_3_13_0_\ : std_logic;
signal \SYNTHESIZED_WIRE_2_1\ : std_logic;
signal \b2v_inst4.un1_pix_count_int_cry_0\ : std_logic;
signal \SYNTHESIZED_WIRE_2_2\ : std_logic;
signal \b2v_inst4.un1_pix_count_int_cry_1\ : std_logic;
signal \SYNTHESIZED_WIRE_2_3\ : std_logic;
signal \b2v_inst4.pix_count_int_RNO_0Z0Z_3\ : std_logic;
signal \b2v_inst4.un1_pix_count_int_cry_2\ : std_logic;
signal \SYNTHESIZED_WIRE_2_4\ : std_logic;
signal \b2v_inst4.un1_pix_count_int_cry_3\ : std_logic;
signal \SYNTHESIZED_WIRE_2_5\ : std_logic;
signal \b2v_inst4.pix_count_int_RNO_0Z0Z_5\ : std_logic;
signal \b2v_inst4.un1_pix_count_int_cry_4\ : std_logic;
signal \SYNTHESIZED_WIRE_2_6\ : std_logic;
signal \b2v_inst4.un1_pix_count_int_cry_5\ : std_logic;
signal \SYNTHESIZED_WIRE_2_7\ : std_logic;
signal \b2v_inst4.pix_count_int_RNO_0Z0Z_7\ : std_logic;
signal \b2v_inst4.un1_pix_count_int_cry_6\ : std_logic;
signal \b2v_inst4.un1_pix_count_int_cry_7\ : std_logic;
signal \SYNTHESIZED_WIRE_2_8\ : std_logic;
signal \b2v_inst4.pix_count_int_RNO_0Z0Z_8\ : std_logic;
signal \bfn_3_14_0_\ : std_logic;
signal \b2v_inst4.un1_pix_count_int_cry_8\ : std_logic;
signal \SYNTHESIZED_WIRE_2_10\ : std_logic;
signal \b2v_inst4.un1_pix_count_int_cry_9\ : std_logic;
signal \SYNTHESIZED_WIRE_2_11\ : std_logic;
signal \b2v_inst4.pix_count_int_RNO_0Z0Z_11\ : std_logic;
signal \b2v_inst4.un1_pix_count_int_cry_10\ : std_logic;
signal \SYNTHESIZED_WIRE_2_12\ : std_logic;
signal \b2v_inst4.un1_pix_count_int_cry_11\ : std_logic;
signal \b2v_inst4.pix_count_int_RNO_0Z0Z_12\ : std_logic;
signal \b2v_inst.data_a_escribir9_0_and\ : std_logic;
signal \bfn_3_15_0_\ : std_logic;
signal \b2v_inst.data_a_escribir9_1_and\ : std_logic;
signal \b2v_inst.data_a_escribir9_0\ : std_logic;
signal \b2v_inst.data_a_escribir9_2_and\ : std_logic;
signal \b2v_inst.data_a_escribir9_1\ : std_logic;
signal \b2v_inst.data_a_escribir9_3_and\ : std_logic;
signal \b2v_inst.data_a_escribir9_2\ : std_logic;
signal \b2v_inst.data_a_escribir9_3\ : std_logic;
signal \b2v_inst.data_a_escribir9_4\ : std_logic;
signal \b2v_inst.data_a_escribir9_5\ : std_logic;
signal \b2v_inst.data_a_escribir9_6\ : std_logic;
signal \b2v_inst.data_a_escribir10\ : std_logic;
signal \bfn_3_16_0_\ : std_logic;
signal \b2v_inst.eventosZ0Z_7\ : std_logic;
signal \b2v_inst.eventosZ0Z_1\ : std_logic;
signal \b2v_inst.eventosZ0Z_6\ : std_logic;
signal \b2v_inst.un1_reg_anterior_iv_0_0_2_1_1_cascade_\ : std_logic;
signal \b2v_inst.data_a_escribir_RNO_4Z0Z_1_cascade_\ : std_logic;
signal \b2v_inst.un1_reg_anterior_iv_0_0_0_1\ : std_logic;
signal \b2v_inst.data_a_escribir_RNO_0Z0Z_1\ : std_logic;
signal \b2v_inst.data_a_escribir_RNO_1Z0Z_1_cascade_\ : std_logic;
signal \b2v_inst.N_497\ : std_logic;
signal \b2v_inst.un1_reg_anterior_iv_0_0_2_tz_2\ : std_logic;
signal \b2v_inst.data_a_escribir_RNO_1Z0Z_2_cascade_\ : std_logic;
signal \b2v_inst.un1_reg_anterior_iv_0_0_1_2\ : std_logic;
signal \b2v_inst.data_a_escribir_RNO_4Z0Z_5_cascade_\ : std_logic;
signal \b2v_inst.un1_reg_anterior_iv_0_0_2_1_5_cascade_\ : std_logic;
signal \b2v_inst.un1_reg_anterior_iv_0_0_a2_4_0_1\ : std_logic;
signal \b2v_inst.un1_reg_anterior_iv_0_0_0_5\ : std_logic;
signal \b2v_inst.data_a_escribir_RNO_0Z0Z_5_cascade_\ : std_logic;
signal \b2v_inst.data_a_escribir_RNO_1Z0Z_5\ : std_logic;
signal \b2v_inst.reg_anterior_i_0\ : std_logic;
signal \bfn_3_19_0_\ : std_logic;
signal \b2v_inst.reg_anterior_i_1\ : std_logic;
signal \b2v_inst.valor_max_final5_1_cry_0\ : std_logic;
signal \b2v_inst.reg_anterior_i_2\ : std_logic;
signal \b2v_inst.valor_max_final5_1_cry_1\ : std_logic;
signal \b2v_inst.reg_anterior_i_3\ : std_logic;
signal \b2v_inst.valor_max_final5_1_cry_2\ : std_logic;
signal \b2v_inst.reg_anterior_i_4\ : std_logic;
signal \b2v_inst.valor_max_final5_1_cry_3\ : std_logic;
signal \b2v_inst.reg_anterior_i_5\ : std_logic;
signal \b2v_inst.valor_max_final5_1_cry_4\ : std_logic;
signal \b2v_inst.reg_anterior_i_6\ : std_logic;
signal \b2v_inst.valor_max_final5_1_cry_5\ : std_logic;
signal \b2v_inst.reg_anterior_i_7\ : std_logic;
signal \b2v_inst.valor_max_final5_1_cry_6\ : std_logic;
signal \b2v_inst.valor_max_final51\ : std_logic;
signal \b2v_inst.valor_max_final53_THRU_CO\ : std_logic;
signal \b2v_inst.un1_m3_0_m3_ns_1\ : std_logic;
signal \bfn_3_20_0_\ : std_logic;
signal \b2v_inst.un1_reg_anterior_iv_0_0_2_tz_4\ : std_logic;
signal \b2v_inst3.fsm_state_ns_0_0_0_1_cascade_\ : std_logic;
signal \N_230_cascade_\ : std_logic;
signal \b2v_inst3.N_434\ : std_logic;
signal \b2v_inst3.N_490\ : std_logic;
signal \b2v_inst3.fsm_state_ns_i_i_1_0_cascade_\ : std_logic;
signal \b2v_inst3.un1_m2_0_a2_2_cascade_\ : std_logic;
signal \b2v_inst3.un1_cycle_counter_5_c5\ : std_logic;
signal \b2v_inst3.un1_cycle_counter_5_c5_cascade_\ : std_logic;
signal \SYNTHESIZED_WIRE_10_0\ : std_logic;
signal \SYNTHESIZED_WIRE_3_0\ : std_logic;
signal \SYNTHESIZED_WIRE_3_1\ : std_logic;
signal \SYNTHESIZED_WIRE_3_2\ : std_logic;
signal \SYNTHESIZED_WIRE_3_3\ : std_logic;
signal \SYNTHESIZED_WIRE_3_4\ : std_logic;
signal \SYNTHESIZED_WIRE_3_5\ : std_logic;
signal \SYNTHESIZED_WIRE_3_6\ : std_logic;
signal \SYNTHESIZED_WIRE_3_7\ : std_logic;
signal \b2v_inst4.pix_count_int_0_sqmuxa\ : std_logic;
signal \b2v_inst.we_0_a2_0_a2_4_cascade_\ : std_logic;
signal \SYNTHESIZED_WIRE_4\ : std_logic;
signal \b2v_inst.we_0_a2_0_a2_3\ : std_logic;
signal \N_458_cascade_\ : std_logic;
signal \b2v_inst.N_429_cascade_\ : std_logic;
signal \b2v_inst.un1_pix_count_anterior_0_N_2_THRU_CO\ : std_logic;
signal \b2v_inst.stateZ0Z_3\ : std_logic;
signal \b2v_inst.stateZ0Z_2\ : std_logic;
signal \b2v_inst.data_a_escribir9_4_and\ : std_logic;
signal \b2v_inst.data_a_escribir9_5_and\ : std_logic;
signal \b2v_inst.un3_valor_max1_THRU_CO\ : std_logic;
signal \b2v_inst.data_a_escribir_RNO_3Z0Z_6\ : std_logic;
signal \b2v_inst.un1_reg_anterior_iv_0_0_a2_6_0_1\ : std_logic;
signal \b2v_inst.un1_m3_0_0\ : std_logic;
signal \b2v_inst.un1_reg_anterior_iv_0_0_0_6\ : std_logic;
signal \b2v_inst.data_a_escribir_RNO_1Z0Z_6_cascade_\ : std_logic;
signal \b2v_inst.data_a_escribir10_THRU_CO\ : std_logic;
signal \b2v_inst.N_264\ : std_logic;
signal \b2v_inst.un1_reg_anterior_iv_0_0_0_7\ : std_logic;
signal \b2v_inst.un1_reg_anterior_iv_0_0_3_0_7_cascade_\ : std_logic;
signal \b2v_inst.un1_reg_anterior_iv_0_0_2_0_tz_7\ : std_logic;
signal \b2v_inst.un1_reset_inv_2_0\ : std_logic;
signal \b2v_inst.reg_ancho_1Z0Z_0\ : std_logic;
signal \b2v_inst.reg_ancho_3Z0Z_0\ : std_logic;
signal \bfn_5_17_0_\ : std_logic;
signal \b2v_inst.reg_ancho_1Z0Z_1\ : std_logic;
signal \b2v_inst.reg_ancho_3Z0Z_1\ : std_logic;
signal \b2v_inst.valor_max_final5_0_cry_0\ : std_logic;
signal \b2v_inst.reg_ancho_3Z0Z_2\ : std_logic;
signal \b2v_inst.reg_ancho_1Z0Z_2\ : std_logic;
signal \b2v_inst.valor_max_final5_0_cry_1\ : std_logic;
signal \b2v_inst.reg_ancho_1Z0Z_3\ : std_logic;
signal \b2v_inst.reg_ancho_3Z0Z_3\ : std_logic;
signal \b2v_inst.valor_max_final5_0_cry_2\ : std_logic;
signal \b2v_inst.reg_ancho_1Z0Z_4\ : std_logic;
signal \b2v_inst.reg_ancho_3Z0Z_4\ : std_logic;
signal \b2v_inst.valor_max_final5_0_cry_3\ : std_logic;
signal \b2v_inst.reg_ancho_1Z0Z_5\ : std_logic;
signal \b2v_inst.valor_max_final5_0_cry_4\ : std_logic;
signal \b2v_inst.reg_ancho_1Z0Z_6\ : std_logic;
signal \b2v_inst.valor_max_final5_0_cry_5\ : std_logic;
signal \b2v_inst.reg_ancho_1Z0Z_7\ : std_logic;
signal \b2v_inst.reg_ancho_3Z0Z_7\ : std_logic;
signal \b2v_inst.valor_max_final5_0_cry_6\ : std_logic;
signal \b2v_inst.valor_max_final50\ : std_logic;
signal \bfn_5_18_0_\ : std_logic;
signal \b2v_inst.valor_max_final50_THRU_CO\ : std_logic;
signal \b2v_inst.data_a_escribir9_6_and\ : std_logic;
signal \b2v_inst.reg_ancho_2Z0Z_0\ : std_logic;
signal \bfn_5_19_0_\ : std_logic;
signal \b2v_inst.reg_ancho_2Z0Z_1\ : std_logic;
signal \b2v_inst.valor_max_final5_2_cry_0\ : std_logic;
signal \b2v_inst.reg_ancho_2Z0Z_2\ : std_logic;
signal \b2v_inst.valor_max_final5_2_cry_1\ : std_logic;
signal \b2v_inst.reg_ancho_2Z0Z_3\ : std_logic;
signal \b2v_inst.valor_max_final5_2_cry_2\ : std_logic;
signal \b2v_inst.reg_ancho_2Z0Z_4\ : std_logic;
signal \b2v_inst.valor_max_final5_2_cry_3\ : std_logic;
signal \b2v_inst.reg_ancho_2Z0Z_5\ : std_logic;
signal \b2v_inst.valor_max_final5_2_cry_4\ : std_logic;
signal \b2v_inst.reg_ancho_2Z0Z_6\ : std_logic;
signal \b2v_inst.valor_max_final5_2_cry_5\ : std_logic;
signal \b2v_inst.reg_ancho_2Z0Z_7\ : std_logic;
signal \b2v_inst.valor_max_final5_2_cry_6\ : std_logic;
signal \b2v_inst.valor_max_final52\ : std_logic;
signal \bfn_5_20_0_\ : std_logic;
signal \b2v_inst.valor_max_final52_THRU_CO\ : std_logic;
signal \b2v_inst3.un1_bit_counter_3_c2\ : std_logic;
signal \b2v_inst3.un1_bit_counter_3_c2_cascade_\ : std_logic;
signal \b2v_inst3.N_258\ : std_logic;
signal \b2v_inst3.N_258_cascade_\ : std_logic;
signal \b2v_inst3.bit_counterZ0Z_2\ : std_logic;
signal \b2v_inst3.bit_counterZ1Z_1\ : std_logic;
signal \b2v_inst3.N_102_2_cascade_\ : std_logic;
signal \b2v_inst3.bit_counterZ0Z_3\ : std_logic;
signal \b2v_inst3.N_436\ : std_logic;
signal uart_tx_o : std_logic;
signal \b2v_inst4.stateZ0Z_0\ : std_logic;
signal \b2v_inst3.cycle_counterZ0Z_6\ : std_logic;
signal \b2v_inst3.cycle_counterZ0Z_5\ : std_logic;
signal \b2v_inst3.cycle_counterZ0Z_7\ : std_logic;
signal \b2v_inst3.next_bit_0_a3_4_cascade_\ : std_logic;
signal \b2v_inst3.next_bit_0_a3_3\ : std_logic;
signal \SYNTHESIZED_WIRE_7\ : std_logic;
signal \b2v_inst3.N_105_7_cascade_\ : std_logic;
signal \b2v_inst3.fsm_stateZ0Z_0\ : std_logic;
signal \b2v_inst3.cycle_counterZ0Z_1\ : std_logic;
signal \b2v_inst3.fsm_stateZ0Z_1\ : std_logic;
signal \b2v_inst3.cycle_counterZ0Z_0\ : std_logic;
signal \b2v_inst3.un1_cycle_counter_5_c2\ : std_logic;
signal \b2v_inst3.cycle_counterZ0Z_2\ : std_logic;
signal \b2v_inst3.cycle_counterZ0Z_3\ : std_logic;
signal \b2v_inst3.un1_cycle_counter_5_c2_cascade_\ : std_logic;
signal \b2v_inst3.cycle_counterZ0Z_4\ : std_logic;
signal \b2v_inst4.un1_pix_count_int_0_sqmuxa_9\ : std_logic;
signal \b2v_inst4.un1_pix_count_int_0_sqmuxa_11\ : std_logic;
signal \b2v_inst4.un1_pix_count_int_0_sqmuxa_10\ : std_logic;
signal \b2v_inst4.pix_count_int_RNO_0Z0Z_9\ : std_logic;
signal \SYNTHESIZED_WIRE_2_9\ : std_logic;
signal \b2v_inst.cuenta_pixelZ0Z_6\ : std_logic;
signal \b2v_inst.un11_cuenta_pixel_i_0_o2_0\ : std_logic;
signal \b2v_inst.cuenta_pixelZ0Z_5\ : std_logic;
signal \b2v_inst.cuenta_pixelZ0Z_0\ : std_logic;
signal \b2v_inst.cuenta_pixelZ0Z_1\ : std_logic;
signal \b2v_inst.cuenta_pixel_4_i_a2_0_6\ : std_logic;
signal \N_213_i\ : std_logic;
signal \N_209_i\ : std_logic;
signal \N_207_i\ : std_logic;
signal \SYNTHESIZED_WIRE_10_2\ : std_logic;
signal \SYNTHESIZED_WIRE_10_3\ : std_logic;
signal \SYNTHESIZED_WIRE_10_4\ : std_logic;
signal \SYNTHESIZED_WIRE_10_5\ : std_logic;
signal \SYNTHESIZED_WIRE_10_6\ : std_logic;
signal \SYNTHESIZED_WIRE_10_7\ : std_logic;
signal \b2v_inst.addr_ram_1_iv_i_2_5_cascade_\ : std_logic;
signal \N_54\ : std_logic;
signal \b2v_inst.addr_ram_1_iv_i_1_5\ : std_logic;
signal \b2v_inst.N_341\ : std_logic;
signal \b2v_inst.N_404_cascade_\ : std_logic;
signal \b2v_inst.reg_ancho_3Z0Z_6\ : std_logic;
signal \b2v_inst.reg_ancho_3Z0Z_5\ : std_logic;
signal \b2v_inst.reg_ancho_3_i_0\ : std_logic;
signal \bfn_6_17_0_\ : std_logic;
signal \b2v_inst.reg_ancho_3_i_1\ : std_logic;
signal \b2v_inst.un3_valor_max2_cry_0\ : std_logic;
signal \b2v_inst.reg_ancho_3_i_2\ : std_logic;
signal \b2v_inst.un3_valor_max2_cry_1\ : std_logic;
signal \b2v_inst.reg_ancho_3_i_3\ : std_logic;
signal \b2v_inst.un3_valor_max2_cry_2\ : std_logic;
signal \b2v_inst.reg_ancho_3_i_4\ : std_logic;
signal \b2v_inst.un3_valor_max2_cry_3\ : std_logic;
signal \b2v_inst.reg_ancho_3_i_5\ : std_logic;
signal \b2v_inst.un3_valor_max2_cry_4\ : std_logic;
signal \b2v_inst.reg_ancho_3_i_6\ : std_logic;
signal \b2v_inst.un3_valor_max2_cry_5\ : std_logic;
signal \b2v_inst.reg_ancho_3_i_7\ : std_logic;
signal \b2v_inst.un3_valor_max2_cry_6\ : std_logic;
signal \b2v_inst.un3_valor_max2\ : std_logic;
signal \bfn_6_18_0_\ : std_logic;
signal \b2v_inst.un3_valor_max2_THRU_CO\ : std_logic;
signal reset_i : std_logic;
signal \b2v_inst3.un2_n_fsm_state_0_sqmuxa_2_0_i\ : std_logic;
signal \b2v_inst1.r_RX_Bytece_0_6\ : std_logic;
signal \SYNTHESIZED_WIRE_1_0\ : std_logic;
signal \b2v_inst.reg_anteriorZ0Z_0\ : std_logic;
signal \SYNTHESIZED_WIRE_1_1\ : std_logic;
signal \b2v_inst.reg_anteriorZ0Z_1\ : std_logic;
signal \SYNTHESIZED_WIRE_1_2\ : std_logic;
signal \b2v_inst.reg_anteriorZ0Z_2\ : std_logic;
signal \SYNTHESIZED_WIRE_1_3\ : std_logic;
signal \b2v_inst.reg_anteriorZ0Z_3\ : std_logic;
signal \SYNTHESIZED_WIRE_1_7\ : std_logic;
signal \b2v_inst.reg_anteriorZ0Z_7\ : std_logic;
signal \b2v_inst.data_a_escribir9_7_and\ : std_logic;
signal \SYNTHESIZED_WIRE_1_4\ : std_logic;
signal \b2v_inst.reg_anteriorZ0Z_4\ : std_logic;
signal b2v_inst_data_a_escribir_1 : std_logic;
signal b2v_inst_data_a_escribir_0 : std_logic;
signal \b2v_inst3.data_to_sendZ0Z_1\ : std_logic;
signal \b2v_inst3.data_to_sendZ0Z_0\ : std_logic;
signal b2v_inst_data_a_escribir_2 : std_logic;
signal \b2v_inst3.data_to_sendZ0Z_2\ : std_logic;
signal \b2v_inst3.fsm_state_RNIEPSN1Z0Z_0\ : std_logic;
signal \b2v_inst3.N_105_7\ : std_logic;
signal \b2v_inst3.bit_counterZ0Z_0\ : std_logic;
signal \b2v_inst.state_ns_a2_0_a2_0_1_2\ : std_logic;
signal \b2v_inst.cuenta_5_i_a2_2_0_1_cascade_\ : std_logic;
signal \b2v_inst.un4_cuenta_c4_cascade_\ : std_logic;
signal \b2v_inst.cuentaZ0Z_3\ : std_logic;
signal \b2v_inst.cuentaZ0Z_2\ : std_logic;
signal \b2v_inst.un2_cuentalto7_3_cascade_\ : std_logic;
signal \b2v_inst.N_351_0_cascade_\ : std_logic;
signal \b2v_inst.cuenta_fastZ0Z_4\ : std_logic;
signal \b2v_inst.cuenta_RNIQ56K_0Z0Z_3\ : std_logic;
signal \b2v_inst.N_376_1\ : std_logic;
signal \b2v_inst.cuenta_RNIQI4FZ0Z_2\ : std_logic;
signal \b2v_inst.cuenta_RNIR03AZ0Z_1\ : std_logic;
signal \b2v_inst.N_376_1_cascade_\ : std_logic;
signal \b2v_inst.cuentaZ0Z_1\ : std_logic;
signal \b2v_inst.cuenta_5_i_a2_0_3\ : std_logic;
signal \b2v_inst.cuentaZ0Z_0\ : std_logic;
signal \b2v_inst.N_377\ : std_logic;
signal \b2v_inst.N_491_cascade_\ : std_logic;
signal \b2v_inst.state_RNIFQKOZ0Z_17\ : std_logic;
signal \b2v_inst.state_RNIFQKOZ0Z_17_cascade_\ : std_logic;
signal \b2v_inst.N_236_cascade_\ : std_logic;
signal \b2v_inst.stateZ0Z_9\ : std_logic;
signal \b2v_inst.N_399_cascade_\ : std_logic;
signal \b2v_inst.addr_ram_1_iv_i_1_6\ : std_logic;
signal \b2v_inst.addr_ram_1_iv_i_2_6_cascade_\ : std_logic;
signal \N_165\ : std_logic;
signal \b2v_inst.stateZ0Z_12\ : std_logic;
signal \b2v_inst.N_235_cascade_\ : std_logic;
signal \b2v_inst.stateZ0Z_11\ : std_logic;
signal \b2v_inst.N_237_cascade_\ : std_logic;
signal \b2v_inst.addr_ram_1_iv_i_2_0\ : std_logic;
signal \b2v_inst.addr_ram_1_iv_i_1_0_cascade_\ : std_logic;
signal \N_167\ : std_logic;
signal \b2v_inst.addr_ram_1_0_iv_i_0_1\ : std_logic;
signal \N_60\ : std_logic;
signal \b2v_inst.addr_ram_1_0_iv_i_0_2_cascade_\ : std_logic;
signal \N_56\ : std_logic;
signal \b2v_inst.dir_mem_315_0_cascade_\ : std_logic;
signal \b2v_inst.dir_mem_3Z0Z_1\ : std_logic;
signal \b2v_inst.addr_ram_1_0_iv_i_1_1\ : std_logic;
signal \b2v_inst.dir_mem_3Z0Z_0\ : std_logic;
signal \b2v_inst.dir_mem_3Z0Z_5\ : std_logic;
signal \b2v_inst.dir_mem_3Z0Z_6\ : std_logic;
signal \N_205_i\ : std_logic;
signal \b2v_inst.dir_mem_2Z0Z_6\ : std_logic;
signal \b2v_inst1.r_RX_Bytece_0_3\ : std_logic;
signal \b2v_inst1.r_RX_Bytece_0_0_4\ : std_logic;
signal b2v_inst_data_a_escribir_3 : std_logic;
signal \b2v_inst3.data_to_sendZ0Z_3\ : std_logic;
signal b2v_inst_data_a_escribir_4 : std_logic;
signal \b2v_inst3.data_to_sendZ0Z_4\ : std_logic;
signal b2v_inst_data_a_escribir_5 : std_logic;
signal \b2v_inst3.data_to_sendZ0Z_5\ : std_logic;
signal b2v_inst_data_a_escribir_6 : std_logic;
signal \b2v_inst3.data_to_sendZ0Z_6\ : std_logic;
signal \N_458\ : std_logic;
signal b2v_inst_data_a_escribir_7 : std_logic;
signal \N_230\ : std_logic;
signal \b2v_inst3.data_to_sendZ0Z_7\ : std_logic;
signal \b2v_inst3.un2_n_fsm_state_0_sqmuxa_2_0_i_0\ : std_logic;
signal \SYNTHESIZED_WIRE_1_6\ : std_logic;
signal \b2v_inst.reg_anteriorZ0Z_6\ : std_logic;
signal \SYNTHESIZED_WIRE_1_5\ : std_logic;
signal \b2v_inst.reg_anteriorZ0Z_5\ : std_logic;
signal \b2v_inst.un4_cuenta_ac0_11_0_cascade_\ : std_logic;
signal \b2v_inst.N_491\ : std_logic;
signal \b2v_inst.cuenta_5_i_o2_0_0_1_cascade_\ : std_logic;
signal \b2v_inst.state_ns_a2_0_o2_1_0_2_cascade_\ : std_logic;
signal \b2v_inst.cuenta_5_i_o2_0_0_1\ : std_logic;
signal \b2v_inst.state_17_rep1_RNICDKZ0Z34_cascade_\ : std_logic;
signal \b2v_inst.cuenta_RNIO2VO3Z0Z_4\ : std_logic;
signal \b2v_inst.N_374\ : std_logic;
signal \b2v_inst.cuentaZ0Z_5\ : std_logic;
signal \b2v_inst.cuentaZ0Z_4\ : std_logic;
signal \b2v_inst.un4_cuenta_ac0_9_0_cascade_\ : std_logic;
signal \b2v_inst.un4_cuenta_c4\ : std_logic;
signal \b2v_inst.cuentaZ0Z_6\ : std_logic;
signal \b2v_inst.cuentaZ0Z_7\ : std_logic;
signal \b2v_inst.N_399_i\ : std_logic;
signal \b2v_inst.N_227\ : std_logic;
signal \b2v_inst.N_232\ : std_logic;
signal \b2v_inst.N_232_cascade_\ : std_logic;
signal \b2v_inst.stateZ0Z_7\ : std_logic;
signal \b2v_inst.stateZ0Z_14\ : std_logic;
signal \b2v_inst.stateZ0Z_6\ : std_logic;
signal \b2v_inst.state_RNITETBZ0Z_0\ : std_logic;
signal \b2v_inst.N_351_cascade_\ : std_logic;
signal \b2v_inst.addr_ram_1_iv_i_1_3\ : std_logic;
signal \b2v_inst.addr_ram_1_iv_i_2_3_cascade_\ : std_logic;
signal \N_58\ : std_logic;
signal \b2v_inst.stateZ0Z_0\ : std_logic;
signal \b2v_inst.stateZ0Z_10\ : std_logic;
signal \b2v_inst.stateZ0Z_1\ : std_logic;
signal \b2v_inst.dir_mem_3Z0Z_4\ : std_logic;
signal \b2v_inst.addr_ram_1_0_iv_i_1_4_cascade_\ : std_logic;
signal \N_163\ : std_logic;
signal \b2v_inst.g0_11_1_cascade_\ : std_logic;
signal \b2v_inst.dir_mem_1Z0Z_4\ : std_logic;
signal \b2v_inst.N_235\ : std_logic;
signal \b2v_inst.addr_ram_1_0_iv_i_0_4\ : std_logic;
signal \b2v_inst.dir_mem_315_0\ : std_logic;
signal \b2v_inst.dir_mem_3Z0Z_3\ : std_logic;
signal \b2v_inst.dir_mem_3Z0Z_7\ : std_logic;
signal \b2v_inst.N_138_i\ : std_logic;
signal \b2v_inst1.r_RX_Bytece_0_5\ : std_logic;
signal \b2v_inst.dir_mem_3_RNO_0Z0Z_3\ : std_logic;
signal \b2v_inst1.r_RX_Bytece_0_0_1_cascade_\ : std_logic;
signal \SYNTHESIZED_WIRE_10_1\ : std_logic;
signal \b2v_inst.dir_mem_2_RNO_0Z0Z_6\ : std_logic;
signal \SYNTHESIZED_WIRE_9\ : std_logic;
signal \b2v_inst.stateZ0Z_16\ : std_logic;
signal \b2v_inst.ignorar_anteriorZ0\ : std_logic;
signal \b2v_inst.un1_state_19_0\ : std_logic;
signal \b2v_inst.N_5\ : std_logic;
signal \b2v_inst.N_7_1_cascade_\ : std_logic;
signal \b2v_inst.g2_2_cascade_\ : std_logic;
signal \b2v_inst.g1\ : std_logic;
signal \b2v_inst.un2_indice_21_s0_0_6\ : std_logic;
signal \b2v_inst.N_253_cascade_\ : std_logic;
signal \b2v_inst.state_fastZ0Z_17\ : std_logic;
signal \b2v_inst.state_fastZ0Z_15\ : std_logic;
signal \b2v_inst.N_253_i_cascade_\ : std_logic;
signal \b2v_inst.un2_indice_3_0_iv_0_a2_5_sx_2\ : std_logic;
signal \b2v_inst.N_452_cascade_\ : std_logic;
signal \b2v_inst.stateZ0Z_13\ : std_logic;
signal \b2v_inst.g2_3\ : std_logic;
signal \b2v_inst.borradoZ0\ : std_logic;
signal \b2v_inst.stateZ0Z_5\ : std_logic;
signal \b2v_inst.g4_0_cascade_\ : std_logic;
signal \b2v_inst.g0_0\ : std_logic;
signal \b2v_inst.state_ns_a2_0_o2_1_0_2\ : std_logic;
signal \b2v_inst.cuenta_RNI4SC81Z0Z_7\ : std_logic;
signal \b2v_inst.state_ns_a2_0_o2_0_2\ : std_logic;
signal \b2v_inst.stateZ0Z_8\ : std_logic;
signal \b2v_inst.dir_mem_2_RNO_0Z0Z_3_cascade_\ : std_logic;
signal \b2v_inst.dir_mem_2Z0Z_3\ : std_logic;
signal \b2v_inst.un1_dir_mem_3_ns_1_4\ : std_logic;
signal \b2v_inst.dir_mem_2_RNO_0Z0Z_7\ : std_logic;
signal \b2v_inst.N_237\ : std_logic;
signal \b2v_inst.dir_mem_2Z0Z_7\ : std_logic;
signal \b2v_inst.N_239\ : std_logic;
signal \b2v_inst.addr_ram_1_0_iv_i_1_7_cascade_\ : std_logic;
signal \b2v_inst.addr_ram_1_0_iv_i_0_7\ : std_logic;
signal \N_50\ : std_logic;
signal \b2v_inst.g0_2_6_cascade_\ : std_logic;
signal \b2v_inst.g0_2_8\ : std_logic;
signal \b2v_inst.i4_mux_cascade_\ : std_logic;
signal \b2v_inst.dir_mem_1Z0Z_6\ : std_logic;
signal \b2v_inst.un2_dir_mem_3_c5\ : std_logic;
signal \b2v_inst.un2_dir_mem_3_ac0_3\ : std_logic;
signal \b2v_inst.un2_dir_mem_3_ac0_3_cascade_\ : std_logic;
signal \b2v_inst.un1_dir_mem_3_ns_1_5\ : std_logic;
signal \b2v_inst.m7_1\ : std_logic;
signal \b2v_inst.un8_dir_mem_3_c4_cascade_\ : std_logic;
signal \b2v_inst.un8_dir_mem_3_c6\ : std_logic;
signal \b2v_inst.un2_indice_1_1_4_cascade_\ : std_logic;
signal \b2v_inst.dir_mem_2Z0Z_4\ : std_logic;
signal \b2v_inst.dir_mem_2Z0Z_1\ : std_logic;
signal \b2v_inst.dir_mem_2Z0Z_2\ : std_logic;
signal \b2v_inst.dir_mem_215_0_cascade_\ : std_logic;
signal \b2v_inst.dir_mem_2Z0Z_0\ : std_logic;
signal \b2v_inst.dir_mem_215_0\ : std_logic;
signal \b2v_inst.dir_mem_2Z0Z_5\ : std_logic;
signal \b2v_inst.N_136_i\ : std_logic;
signal \b2v_inst1.N_14\ : std_logic;
signal \b2v_inst.dir_mem_RNIGVEE1Z0Z_0\ : std_logic;
signal \bfn_10_10_0_\ : std_logic;
signal \b2v_inst.dir_mem_RNII5PO1Z0Z_1\ : std_logic;
signal \b2v_inst.un2_indice_cry_0\ : std_logic;
signal \b2v_inst.dir_mem_RNIL33H1Z0Z_2\ : std_logic;
signal \b2v_inst.un2_indice_cry_1\ : std_logic;
signal \b2v_inst.dir_mem_RNIN53H1Z0Z_3\ : std_logic;
signal \b2v_inst.un2_indice_cry_2\ : std_logic;
signal \b2v_inst.un2_indice_cry_3\ : std_logic;
signal \b2v_inst.un2_indice_cry_4\ : std_logic;
signal \b2v_inst.dir_mem_RNITB3H1Z0Z_6\ : std_logic;
signal \b2v_inst.un2_indice_20_6\ : std_logic;
signal \b2v_inst.un2_indice_cry_5\ : std_logic;
signal \b2v_inst.un2_indice_cry_6\ : std_logic;
signal \b2v_inst.un2_indice_21_s0_1_cascade_\ : std_logic;
signal \b2v_inst.un2_indice_21_s0_1\ : std_logic;
signal \b2v_inst.un2_indice_20_1\ : std_logic;
signal \b2v_inst.dir_mem_RNO_2Z0Z_1\ : std_logic;
signal \b2v_inst.dir_mem_RNO_3Z0Z_1_cascade_\ : std_logic;
signal \b2v_inst.dir_mem_RNIP73H1Z0Z_4\ : std_logic;
signal \b2v_inst.dir_mem_RNIR93H1Z0Z_5\ : std_logic;
signal \b2v_inst.g1_0_3\ : std_logic;
signal \b2v_inst.g0_2_7\ : std_logic;
signal \b2v_inst.N_467\ : std_logic;
signal \b2v_inst.N_411_cascade_\ : std_logic;
signal \b2v_inst.un2_indice_20_5\ : std_logic;
signal \b2v_inst.un2_indice_3_iv_0_a2_2_sx_5\ : std_logic;
signal \b2v_inst.un2_indice_0_d0_c4_d\ : std_logic;
signal \b2v_inst.un2_m1_e_0_cascade_\ : std_logic;
signal \b2v_inst.dir_mem_RNO_4Z0Z_4_cascade_\ : std_logic;
signal \b2v_inst.indice_RNIA33NZ0Z_1\ : std_logic;
signal \b2v_inst.N_238\ : std_logic;
signal \b2v_inst.N_236\ : std_logic;
signal \b2v_inst.dir_mem_3Z0Z_2\ : std_logic;
signal \b2v_inst.addr_ram_1_0_iv_i_1_2\ : std_logic;
signal \b2v_inst.un10_indice_cascade_\ : std_logic;
signal \b2v_inst1.r_RX_Bytece_0_2\ : std_logic;
signal \b2v_inst1.r_RX_Byte_1_sqmuxa\ : std_logic;
signal \b2v_inst1.r_RX_Bytece_0_0_0\ : std_logic;
signal \b2v_inst.indice_3_repZ0Z1\ : std_logic;
signal \b2v_inst.un2_dir_mem_2_c4_d\ : std_logic;
signal \b2v_inst1.N_7_cascade_\ : std_logic;
signal \b2v_inst1.g0_0_i_a6_1_2\ : std_logic;
signal \b2v_inst1.N_9_cascade_\ : std_logic;
signal \b2v_inst1.g0_0_i_a6_3_5\ : std_logic;
signal \b2v_inst1.N_19_cascade_\ : std_logic;
signal \b2v_inst1.N_6\ : std_logic;
signal \b2v_inst1.r_SM_Main_1_sqmuxa_1_0\ : std_logic;
signal \b2v_inst1.g0_3_4\ : std_logic;
signal \b2v_inst1.g0_0_i_a6_2_2_cascade_\ : std_logic;
signal \b2v_inst1.g0_0_i_a6_2_1\ : std_logic;
signal \b2v_inst1.N_18\ : std_logic;
signal \b2v_inst.dir_mem_RNO_2Z0Z_4\ : std_logic;
signal \b2v_inst.un2_indice_3_0_i_1_4_cascade_\ : std_logic;
signal \b2v_inst.un2_indice_20_4\ : std_logic;
signal \b2v_inst.dir_mem_RNO_2Z0Z_7\ : std_logic;
signal \b2v_inst.un2_indice_20_7\ : std_logic;
signal \b2v_inst.un2_indice_3_0_iv_0_0_7_cascade_\ : std_logic;
signal \b2v_inst.un2_indice_21_s0_2\ : std_logic;
signal \b2v_inst.un2_indice_20_2\ : std_logic;
signal \b2v_inst.un2_indice_21_s1_2\ : std_logic;
signal \b2v_inst.un2_indice_3_0_iv_0_1_2_cascade_\ : std_logic;
signal \b2v_inst.dir_mem_RNO_3Z0Z_4\ : std_logic;
signal \b2v_inst.un2_indice_0_d1_c2\ : std_logic;
signal \b2v_inst.N_451\ : std_logic;
signal \b2v_inst.un2_indice_21_s0_3\ : std_logic;
signal \b2v_inst.un2_indice_20_3\ : std_logic;
signal \b2v_inst.un2_indice_21_s1_3\ : std_logic;
signal \b2v_inst.un2_indice_3_0_iv_0_0_3_cascade_\ : std_logic;
signal \b2v_inst.dir_mem_RNO_5Z0Z_4\ : std_logic;
signal \b2v_inst.un2_indice_3_iv_0_1_0_5\ : std_logic;
signal \b2v_inst.N_410\ : std_logic;
signal \b2v_inst.un2_indice_3_iv_0_0_1\ : std_logic;
signal \b2v_inst.N_253_i\ : std_logic;
signal \b2v_inst.stateZ0Z_17\ : std_logic;
signal \b2v_inst.un2_indice_20_0_cascade_\ : std_logic;
signal \b2v_inst.N_4_0\ : std_logic;
signal \b2v_inst.un2_cuentalto7_3\ : std_logic;
signal \b2v_inst.N_228_cascade_\ : std_logic;
signal \b2v_inst.cuenta_RNI925FZ0Z_7\ : std_logic;
signal \b2v_inst.N_234\ : std_logic;
signal \b2v_inst.un2_indice_3_0_iv_0_a2_0_8_2_2\ : std_logic;
signal \b2v_inst.N_228\ : std_logic;
signal \b2v_inst.N_383_8_cascade_\ : std_logic;
signal \b2v_inst.un2_indice_3_0_iv_0_a2_0_8_3_2\ : std_logic;
signal \b2v_inst.un10_indice_2_cascade_\ : std_logic;
signal \b2v_inst.indice_fast_RNIDAJGZ0Z_2\ : std_logic;
signal \b2v_inst.dir_mem_115lto6_1_cascade_\ : std_logic;
signal \b2v_inst.un1_dir_mem_1_mb_1_7_cascade_\ : std_logic;
signal \b2v_inst.dir_mem_1Z0Z_7\ : std_logic;
signal \b2v_inst.indiceZ0Z_4\ : std_logic;
signal \b2v_inst.un2_dir_mem_2_c5\ : std_logic;
signal \b2v_inst.N_4_0_0_cascade_\ : std_logic;
signal \b2v_inst.N_8_0\ : std_logic;
signal \b2v_inst.dir_mem_315lto8_a0_1_cascade_\ : std_logic;
signal \b2v_inst.indice_fast_RNIRFV61Z0Z_3\ : std_logic;
signal \b2v_inst.indice_0_repZ0Z1\ : std_logic;
signal \b2v_inst.indice_0_rep1_RNIFJJGZ0\ : std_logic;
signal \b2v_inst.indice_1_repZ0Z1\ : std_logic;
signal \b2v_inst.indice_fastZ0Z_2\ : std_logic;
signal \b2v_inst.dir_mem_215lt6_0_cascade_\ : std_logic;
signal \b2v_inst.dir_mem_215lt8\ : std_logic;
signal \b2v_inst1.g0_0_i_a6_3_4\ : std_logic;
signal \b2v_inst1.r_rx_byteZ0Z_7\ : std_logic;
signal \b2v_inst1.r_rx_byteZ0Z_7_cascade_\ : std_logic;
signal \b2v_inst1.r_Bit_IndexZ0Z_2\ : std_logic;
signal \b2v_inst1.r_Bit_IndexZ0Z_0\ : std_logic;
signal \b2v_inst1.r_Bit_IndexZ0Z_1\ : std_logic;
signal \b2v_inst1.N_11_0_0\ : std_logic;
signal \b2v_inst1.N_9\ : std_logic;
signal \b2v_inst1.un1_r_Clk_Count_ac0_1_out_cascade_\ : std_logic;
signal \b2v_inst1.m22_ns_1\ : std_logic;
signal \b2v_inst1.N_29_mux_cascade_\ : std_logic;
signal \b2v_inst1.N_11_cascade_\ : std_logic;
signal \b2v_inst1.g0_0_i_1\ : std_logic;
signal \b2v_inst1.N_14_0\ : std_logic;
signal \b2v_inst1.g0_0_i_0\ : std_logic;
signal \b2v_inst1.m6_2_cascade_\ : std_logic;
signal \b2v_inst1.N_10_0\ : std_logic;
signal \b2v_inst1.g0_7_1\ : std_logic;
signal \b2v_inst1.g0_i_1_cascade_\ : std_logic;
signal \b2v_inst1.N_11_0\ : std_logic;
signal \b2v_inst1.N_32_mux\ : std_logic;
signal \b2v_inst1.N_10_cascade_\ : std_logic;
signal \b2v_inst1.g2_1_cascade_\ : std_logic;
signal \b2v_inst1.g2_0\ : std_logic;
signal \b2v_inst1.m6_2\ : std_logic;
signal \b2v_inst.un2_indice_0_d1_c5\ : std_logic;
signal \b2v_inst.dir_memZ0Z_4\ : std_logic;
signal \b2v_inst.un2_indice_0_d1_ac0_7_s_0_0\ : std_logic;
signal \b2v_inst.dir_memZ0Z_3\ : std_logic;
signal \b2v_inst.dir_memZ0Z_5\ : std_logic;
signal \b2v_inst.un2_indice_0_d1_ac0_7_s_0_0_cascade_\ : std_logic;
signal \b2v_inst.dir_memZ0Z_2\ : std_logic;
signal \b2v_inst.dir_memZ0Z_7\ : std_logic;
signal \b2v_inst.un2_indice_0_d1_ac0_9_0_cascade_\ : std_logic;
signal \b2v_inst.dir_memZ0Z_6\ : std_logic;
signal \b2v_inst.un2_indice_21_s1_7\ : std_logic;
signal \b2v_inst.state_17_repZ0Z1\ : std_logic;
signal \b2v_inst.stateZ0Z_15\ : std_logic;
signal reset : std_logic;
signal \b2v_inst.N_351_0\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \b2v_inst.N_384_cascade_\ : std_logic;
signal \b2v_inst.state_17_rep1_RNIN75CZ0Z3\ : std_logic;
signal \b2v_inst.un2_indice_3_0_iv_0_0_2\ : std_logic;
signal \b2v_inst.dir_memZ0Z_0\ : std_logic;
signal \b2v_inst.dir_memZ0Z_1\ : std_logic;
signal \b2v_inst.N_253\ : std_logic;
signal \b2v_inst.un2_indice_21_s1_1\ : std_logic;
signal \b2v_inst.un10_indice_2\ : std_logic;
signal \b2v_inst.CO1\ : std_logic;
signal \b2v_inst.CO1_cascade_\ : std_logic;
signal \b2v_inst.un2_dir_mem_2_c2_cascade_\ : std_logic;
signal \b2v_inst.indice_fastZ0Z_0\ : std_logic;
signal \b2v_inst.indice_fastZ0Z_1\ : std_logic;
signal \b2v_inst.indice_2_repZ0Z1\ : std_logic;
signal \b2v_inst.indiceZ0Z_3\ : std_logic;
signal \b2v_inst.dir_mem_1_RNO_0Z0Z_3_cascade_\ : std_logic;
signal \b2v_inst.dir_mem_1Z0Z_3\ : std_logic;
signal \b2v_inst.indice_fast_RNIF91EZ0Z_0\ : std_logic;
signal \b2v_inst.dir_mem_115lto8_1\ : std_logic;
signal \b2v_inst.dir_mem_115lto6_1\ : std_logic;
signal \b2v_inst.un8_dir_mem_1_c7\ : std_logic;
signal \b2v_inst.dir_mem_115lto8_1_cascade_\ : std_logic;
signal \b2v_inst.dir_mem_115_0_cascade_\ : std_logic;
signal \b2v_inst.dir_mem_1Z0Z_0\ : std_logic;
signal \b2v_inst.indiceZ0Z_2\ : std_logic;
signal \b2v_inst.un2_dir_mem_2_c2\ : std_logic;
signal \b2v_inst.dir_mem_1Z0Z_2\ : std_logic;
signal \b2v_inst.dir_mem_1_RNO_0Z0Z_5\ : std_logic;
signal \b2v_inst.dir_mem_1Z0Z_5\ : std_logic;
signal \b2v_inst.dir_mem_115_0\ : std_logic;
signal \b2v_inst.dir_mem_1Z0Z_1\ : std_logic;
signal \b2v_inst.N_134_i\ : std_logic;
signal \b2v_inst.un8_dir_mem_3_ac0_9_0_cascade_\ : std_logic;
signal \b2v_inst.un10_indice\ : std_logic;
signal \b2v_inst.indice_4_repZ0Z1\ : std_logic;
signal \b2v_inst.indice_1_repZ0Z2\ : std_logic;
signal \b2v_inst.indice_0_repZ0Z2\ : std_logic;
signal \b2v_inst.un10_indice_2_0\ : std_logic;
signal \b2v_inst.un8_dir_mem_3_ac0_9_0\ : std_logic;
signal \b2v_inst.indiceZ0Z_7\ : std_logic;
signal \b2v_inst.un8_dir_mem_3_c4\ : std_logic;
signal \b2v_inst.indice_fastZ0Z_4\ : std_logic;
signal \b2v_inst.indice_fastZ0Z_3\ : std_logic;
signal \b2v_inst.un8_dir_mem_1_ac0_7_out\ : std_logic;
signal \b2v_inst.un8_dir_mem_2_c4\ : std_logic;
signal \b2v_inst.indiceZ0Z_6\ : std_logic;
signal \b2v_inst.indiceZ0Z_5\ : std_logic;
signal \b2v_inst.dir_mem_2_RNO_1Z0Z_6\ : std_logic;
signal \b2v_inst1.g0_i_o5_0_2\ : std_logic;
signal \b2v_inst1.g0_1_4_cascade_\ : std_logic;
signal \b2v_inst1.N_28_mux\ : std_logic;
signal \b2v_inst1.un1_r_SM_Main_3_0\ : std_logic;
signal \b2v_inst1.g0_1_cascade_\ : std_logic;
signal \b2v_inst1.N_29_mux_1\ : std_logic;
signal \b2v_inst1.N_14_0_1_cascade_\ : std_logic;
signal \b2v_inst1.g0_0_i_a6_1_5_cascade_\ : std_logic;
signal \b2v_inst1.g0_0_i_a6_1_1\ : std_logic;
signal \b2v_inst1.un1_r_Clk_Count_ac0_3_out\ : std_logic;
signal \b2v_inst1.N_29_mux\ : std_logic;
signal \b2v_inst1.r_SM_Main_1_sqmuxa_1_cascade_\ : std_logic;
signal \b2v_inst1.un1_r_SM_Main_1_sqmuxa_0\ : std_logic;
signal \b2v_inst1.un1_r_Clk_Count_ac0_1_out\ : std_logic;
signal \b2v_inst1.r_Clk_CountZ0Z_3\ : std_logic;
signal \b2v_inst1.g0_3_1_cascade_\ : std_logic;
signal \b2v_inst1.N_14_0_0\ : std_logic;
signal \b2v_inst1.N_14_0_0_cascade_\ : std_logic;
signal \b2v_inst1.N_29_mux_0\ : std_logic;
signal \b2v_inst1.r_Clk_CountZ0Z_0\ : std_logic;
signal \b2v_inst1.g3_1_cascade_\ : std_logic;
signal \b2v_inst1.r_Clk_CountZ0Z_1\ : std_logic;
signal \b2v_inst1.g3\ : std_logic;
signal \b2v_inst1.N_9_0\ : std_logic;
signal \b2v_inst1.N_13_cascade_\ : std_logic;
signal \b2v_inst1.g0_0_i_a6_3_0\ : std_logic;
signal \b2v_inst1.g0_0_i_a6_1_6\ : std_logic;
signal \b2v_inst1.g0_0_i_1_0_cascade_\ : std_logic;
signal \b2v_inst1.N_7_0\ : std_logic;
signal \b2v_inst1.r_SM_Main_d_4\ : std_logic;
signal \b2v_inst1.r_Clk_CountZ0Z_6\ : std_logic;
signal \b2v_inst1.r_Clk_CountZ0Z_5\ : std_logic;
signal \b2v_inst1.r_Clk_CountZ0Z_2\ : std_logic;
signal \b2v_inst1.g2_1_4\ : std_logic;
signal \b2v_inst1.r_SM_MainZ0Z_0\ : std_logic;
signal \b2v_inst1.r_SM_MainZ0Z_1\ : std_logic;
signal \b2v_inst1.r_SM_MainZ0Z_2\ : std_logic;
signal \b2v_inst1.N_11_1\ : std_logic;
signal \b2v_inst1.g0_0_i_a6_2_0_cascade_\ : std_logic;
signal \b2v_inst1.r_Clk_CountZ0Z_4\ : std_logic;
signal \b2v_inst1.g0_0_i_0_0\ : std_logic;
signal \b2v_inst.indiceZ0Z_0\ : std_logic;
signal \b2v_inst.indiceZ0Z_1\ : std_logic;
signal \b2v_inst.state_g_2\ : std_logic;
signal reset_i_g : std_logic;
signal uart_rx_i : std_logic;
signal \b2v_inst1.r_RX_Data_RZ0\ : std_logic;
signal \b2v_inst1.r_RX_DataZ0\ : std_logic;
signal clk : std_logic;
signal \_gnd_net_\ : std_logic;

signal uart_tx_o_wire : std_logic;
signal uart_rx_i_wire : std_logic;
signal reset_wire : std_logic;
signal clk_wire : std_logic;
signal \b2v_inst2.mem_0_mem_0_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \b2v_inst2.mem_0_mem_0_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \b2v_inst2.mem_0_mem_0_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \b2v_inst2.mem_0_mem_0_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \b2v_inst2.mem_0_mem_0_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);

begin
    uart_tx_o <= uart_tx_o_wire;
    uart_rx_i_wire <= uart_rx_i;
    reset_wire <= reset;
    clk_wire <= clk;
    \SYNTHESIZED_WIRE_1_7\ <= \b2v_inst2.mem_0_mem_0_0_0_physical_RDATA_wire\(7);
    \SYNTHESIZED_WIRE_1_6\ <= \b2v_inst2.mem_0_mem_0_0_0_physical_RDATA_wire\(6);
    \SYNTHESIZED_WIRE_1_5\ <= \b2v_inst2.mem_0_mem_0_0_0_physical_RDATA_wire\(5);
    \SYNTHESIZED_WIRE_1_4\ <= \b2v_inst2.mem_0_mem_0_0_0_physical_RDATA_wire\(4);
    \SYNTHESIZED_WIRE_1_3\ <= \b2v_inst2.mem_0_mem_0_0_0_physical_RDATA_wire\(3);
    \SYNTHESIZED_WIRE_1_2\ <= \b2v_inst2.mem_0_mem_0_0_0_physical_RDATA_wire\(2);
    \SYNTHESIZED_WIRE_1_1\ <= \b2v_inst2.mem_0_mem_0_0_0_physical_RDATA_wire\(1);
    \SYNTHESIZED_WIRE_1_0\ <= \b2v_inst2.mem_0_mem_0_0_0_physical_RDATA_wire\(0);
    \b2v_inst2.mem_0_mem_0_0_0_physical_RADDR_wire\ <= '0'&'0'&'0'&\N__16330\&\N__13937\&\N__12541\&\N__15416\&\N__15107\&\N__13999\&\N__14026\&\N__14059\;
    \b2v_inst2.mem_0_mem_0_0_0_physical_WADDR_wire\ <= '0'&'0'&'0'&\N__16334\&\N__13936\&\N__12542\&\N__15412\&\N__15103\&\N__14000\&\N__14027\&\N__14060\;
    \b2v_inst2.mem_0_mem_0_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \b2v_inst2.mem_0_mem_0_0_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__14126\&\N__12362\&\N__12374\&\N__9047\&\N__12386\&\N__9008\&\N__9020\&\N__9035\;

    \b2v_inst2.mem_0_mem_0_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 0,
            READ_MODE => 0,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \b2v_inst2.mem_0_mem_0_0_0_physical_RDATA_wire\,
            RADDR => \b2v_inst2.mem_0_mem_0_0_0_physical_RADDR_wire\,
            WADDR => \b2v_inst2.mem_0_mem_0_0_0_physical_WADDR_wire\,
            MASK => \b2v_inst2.mem_0_mem_0_0_0_physical_MASK_wire\,
            WDATA => \b2v_inst2.mem_0_mem_0_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22577\,
            RE => \N__18613\,
            WCLKE => \N__9992\,
            WCLK => \N__22483\,
            WE => \N__18620\
        );

    \ipInertedIOPad_uart_tx_o_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24159\,
            DIN => \N__24158\,
            DOUT => \N__24157\,
            PACKAGEPIN => uart_tx_o_wire
        );

    \ipInertedIOPad_uart_tx_o_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24159\,
            PADOUT => \N__24158\,
            PADIN => \N__24157\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__11735\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_uart_rx_i_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24150\,
            DIN => \N__24149\,
            DOUT => \N__24148\,
            PACKAGEPIN => uart_rx_i_wire
        );

    \ipInertedIOPad_uart_rx_i_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24150\,
            PADOUT => \N__24149\,
            PADIN => \N__24148\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => uart_rx_i,
            DIN1 => OPEN
        );

    \ipInertedIOPad_reset_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24141\,
            DIN => \N__24140\,
            DOUT => \N__24139\,
            PACKAGEPIN => reset_wire
        );

    \ipInertedIOPad_reset_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24141\,
            PADOUT => \N__24140\,
            PADIN => \N__24139\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => reset,
            DIN1 => OPEN
        );

    \ipInertedIOPad_clk_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24132\,
            DIN => \N__24131\,
            DOUT => \N__24130\,
            PACKAGEPIN => clk_wire
        );

    \ipInertedIOPad_clk_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24132\,
            PADOUT => \N__24131\,
            PADIN => \N__24130\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => clk,
            DIN1 => OPEN
        );

    \I__5972\ : InMux
    port map (
            O => \N__24113\,
            I => \N__24110\
        );

    \I__5971\ : LocalMux
    port map (
            O => \N__24110\,
            I => \N__24107\
        );

    \I__5970\ : Odrv4
    port map (
            O => \N__24107\,
            I => \b2v_inst1.g0_0_i_a6_1_6\
        );

    \I__5969\ : CascadeMux
    port map (
            O => \N__24104\,
            I => \b2v_inst1.g0_0_i_1_0_cascade_\
        );

    \I__5968\ : InMux
    port map (
            O => \N__24101\,
            I => \N__24098\
        );

    \I__5967\ : LocalMux
    port map (
            O => \N__24098\,
            I => \b2v_inst1.N_7_0\
        );

    \I__5966\ : SRMux
    port map (
            O => \N__24095\,
            I => \N__24089\
        );

    \I__5965\ : SRMux
    port map (
            O => \N__24094\,
            I => \N__24086\
        );

    \I__5964\ : SRMux
    port map (
            O => \N__24093\,
            I => \N__24083\
        );

    \I__5963\ : SRMux
    port map (
            O => \N__24092\,
            I => \N__24078\
        );

    \I__5962\ : LocalMux
    port map (
            O => \N__24089\,
            I => \N__24073\
        );

    \I__5961\ : LocalMux
    port map (
            O => \N__24086\,
            I => \N__24073\
        );

    \I__5960\ : LocalMux
    port map (
            O => \N__24083\,
            I => \N__24070\
        );

    \I__5959\ : SRMux
    port map (
            O => \N__24082\,
            I => \N__24067\
        );

    \I__5958\ : SRMux
    port map (
            O => \N__24081\,
            I => \N__24064\
        );

    \I__5957\ : LocalMux
    port map (
            O => \N__24078\,
            I => \N__24060\
        );

    \I__5956\ : Span4Mux_v
    port map (
            O => \N__24073\,
            I => \N__24057\
        );

    \I__5955\ : Span4Mux_v
    port map (
            O => \N__24070\,
            I => \N__24054\
        );

    \I__5954\ : LocalMux
    port map (
            O => \N__24067\,
            I => \N__24051\
        );

    \I__5953\ : LocalMux
    port map (
            O => \N__24064\,
            I => \N__24048\
        );

    \I__5952\ : SRMux
    port map (
            O => \N__24063\,
            I => \N__24045\
        );

    \I__5951\ : Span12Mux_s10_v
    port map (
            O => \N__24060\,
            I => \N__24042\
        );

    \I__5950\ : Sp12to4
    port map (
            O => \N__24057\,
            I => \N__24037\
        );

    \I__5949\ : Sp12to4
    port map (
            O => \N__24054\,
            I => \N__24037\
        );

    \I__5948\ : Span4Mux_v
    port map (
            O => \N__24051\,
            I => \N__24032\
        );

    \I__5947\ : Span4Mux_h
    port map (
            O => \N__24048\,
            I => \N__24032\
        );

    \I__5946\ : LocalMux
    port map (
            O => \N__24045\,
            I => \N__24029\
        );

    \I__5945\ : Odrv12
    port map (
            O => \N__24042\,
            I => \b2v_inst1.r_SM_Main_d_4\
        );

    \I__5944\ : Odrv12
    port map (
            O => \N__24037\,
            I => \b2v_inst1.r_SM_Main_d_4\
        );

    \I__5943\ : Odrv4
    port map (
            O => \N__24032\,
            I => \b2v_inst1.r_SM_Main_d_4\
        );

    \I__5942\ : Odrv12
    port map (
            O => \N__24029\,
            I => \b2v_inst1.r_SM_Main_d_4\
        );

    \I__5941\ : InMux
    port map (
            O => \N__24020\,
            I => \N__24011\
        );

    \I__5940\ : InMux
    port map (
            O => \N__24019\,
            I => \N__24006\
        );

    \I__5939\ : InMux
    port map (
            O => \N__24018\,
            I => \N__24006\
        );

    \I__5938\ : InMux
    port map (
            O => \N__24017\,
            I => \N__23998\
        );

    \I__5937\ : InMux
    port map (
            O => \N__24016\,
            I => \N__23998\
        );

    \I__5936\ : InMux
    port map (
            O => \N__24015\,
            I => \N__23993\
        );

    \I__5935\ : InMux
    port map (
            O => \N__24014\,
            I => \N__23993\
        );

    \I__5934\ : LocalMux
    port map (
            O => \N__24011\,
            I => \N__23981\
        );

    \I__5933\ : LocalMux
    port map (
            O => \N__24006\,
            I => \N__23978\
        );

    \I__5932\ : InMux
    port map (
            O => \N__24005\,
            I => \N__23973\
        );

    \I__5931\ : InMux
    port map (
            O => \N__24004\,
            I => \N__23973\
        );

    \I__5930\ : InMux
    port map (
            O => \N__24003\,
            I => \N__23970\
        );

    \I__5929\ : LocalMux
    port map (
            O => \N__23998\,
            I => \N__23965\
        );

    \I__5928\ : LocalMux
    port map (
            O => \N__23993\,
            I => \N__23965\
        );

    \I__5927\ : InMux
    port map (
            O => \N__23992\,
            I => \N__23960\
        );

    \I__5926\ : InMux
    port map (
            O => \N__23991\,
            I => \N__23960\
        );

    \I__5925\ : InMux
    port map (
            O => \N__23990\,
            I => \N__23957\
        );

    \I__5924\ : InMux
    port map (
            O => \N__23989\,
            I => \N__23950\
        );

    \I__5923\ : InMux
    port map (
            O => \N__23988\,
            I => \N__23950\
        );

    \I__5922\ : InMux
    port map (
            O => \N__23987\,
            I => \N__23950\
        );

    \I__5921\ : InMux
    port map (
            O => \N__23986\,
            I => \N__23947\
        );

    \I__5920\ : InMux
    port map (
            O => \N__23985\,
            I => \N__23942\
        );

    \I__5919\ : InMux
    port map (
            O => \N__23984\,
            I => \N__23942\
        );

    \I__5918\ : Odrv4
    port map (
            O => \N__23981\,
            I => \b2v_inst1.r_Clk_CountZ0Z_6\
        );

    \I__5917\ : Odrv4
    port map (
            O => \N__23978\,
            I => \b2v_inst1.r_Clk_CountZ0Z_6\
        );

    \I__5916\ : LocalMux
    port map (
            O => \N__23973\,
            I => \b2v_inst1.r_Clk_CountZ0Z_6\
        );

    \I__5915\ : LocalMux
    port map (
            O => \N__23970\,
            I => \b2v_inst1.r_Clk_CountZ0Z_6\
        );

    \I__5914\ : Odrv4
    port map (
            O => \N__23965\,
            I => \b2v_inst1.r_Clk_CountZ0Z_6\
        );

    \I__5913\ : LocalMux
    port map (
            O => \N__23960\,
            I => \b2v_inst1.r_Clk_CountZ0Z_6\
        );

    \I__5912\ : LocalMux
    port map (
            O => \N__23957\,
            I => \b2v_inst1.r_Clk_CountZ0Z_6\
        );

    \I__5911\ : LocalMux
    port map (
            O => \N__23950\,
            I => \b2v_inst1.r_Clk_CountZ0Z_6\
        );

    \I__5910\ : LocalMux
    port map (
            O => \N__23947\,
            I => \b2v_inst1.r_Clk_CountZ0Z_6\
        );

    \I__5909\ : LocalMux
    port map (
            O => \N__23942\,
            I => \b2v_inst1.r_Clk_CountZ0Z_6\
        );

    \I__5908\ : InMux
    port map (
            O => \N__23921\,
            I => \N__23905\
        );

    \I__5907\ : InMux
    port map (
            O => \N__23920\,
            I => \N__23905\
        );

    \I__5906\ : InMux
    port map (
            O => \N__23919\,
            I => \N__23897\
        );

    \I__5905\ : InMux
    port map (
            O => \N__23918\,
            I => \N__23894\
        );

    \I__5904\ : InMux
    port map (
            O => \N__23917\,
            I => \N__23891\
        );

    \I__5903\ : InMux
    port map (
            O => \N__23916\,
            I => \N__23886\
        );

    \I__5902\ : InMux
    port map (
            O => \N__23915\,
            I => \N__23886\
        );

    \I__5901\ : InMux
    port map (
            O => \N__23914\,
            I => \N__23883\
        );

    \I__5900\ : InMux
    port map (
            O => \N__23913\,
            I => \N__23878\
        );

    \I__5899\ : InMux
    port map (
            O => \N__23912\,
            I => \N__23878\
        );

    \I__5898\ : InMux
    port map (
            O => \N__23911\,
            I => \N__23873\
        );

    \I__5897\ : InMux
    port map (
            O => \N__23910\,
            I => \N__23873\
        );

    \I__5896\ : LocalMux
    port map (
            O => \N__23905\,
            I => \N__23870\
        );

    \I__5895\ : InMux
    port map (
            O => \N__23904\,
            I => \N__23863\
        );

    \I__5894\ : InMux
    port map (
            O => \N__23903\,
            I => \N__23863\
        );

    \I__5893\ : InMux
    port map (
            O => \N__23902\,
            I => \N__23863\
        );

    \I__5892\ : InMux
    port map (
            O => \N__23901\,
            I => \N__23858\
        );

    \I__5891\ : InMux
    port map (
            O => \N__23900\,
            I => \N__23858\
        );

    \I__5890\ : LocalMux
    port map (
            O => \N__23897\,
            I => \b2v_inst1.r_Clk_CountZ0Z_5\
        );

    \I__5889\ : LocalMux
    port map (
            O => \N__23894\,
            I => \b2v_inst1.r_Clk_CountZ0Z_5\
        );

    \I__5888\ : LocalMux
    port map (
            O => \N__23891\,
            I => \b2v_inst1.r_Clk_CountZ0Z_5\
        );

    \I__5887\ : LocalMux
    port map (
            O => \N__23886\,
            I => \b2v_inst1.r_Clk_CountZ0Z_5\
        );

    \I__5886\ : LocalMux
    port map (
            O => \N__23883\,
            I => \b2v_inst1.r_Clk_CountZ0Z_5\
        );

    \I__5885\ : LocalMux
    port map (
            O => \N__23878\,
            I => \b2v_inst1.r_Clk_CountZ0Z_5\
        );

    \I__5884\ : LocalMux
    port map (
            O => \N__23873\,
            I => \b2v_inst1.r_Clk_CountZ0Z_5\
        );

    \I__5883\ : Odrv4
    port map (
            O => \N__23870\,
            I => \b2v_inst1.r_Clk_CountZ0Z_5\
        );

    \I__5882\ : LocalMux
    port map (
            O => \N__23863\,
            I => \b2v_inst1.r_Clk_CountZ0Z_5\
        );

    \I__5881\ : LocalMux
    port map (
            O => \N__23858\,
            I => \b2v_inst1.r_Clk_CountZ0Z_5\
        );

    \I__5880\ : InMux
    port map (
            O => \N__23837\,
            I => \N__23824\
        );

    \I__5879\ : InMux
    port map (
            O => \N__23836\,
            I => \N__23824\
        );

    \I__5878\ : InMux
    port map (
            O => \N__23835\,
            I => \N__23815\
        );

    \I__5877\ : InMux
    port map (
            O => \N__23834\,
            I => \N__23815\
        );

    \I__5876\ : InMux
    port map (
            O => \N__23833\,
            I => \N__23810\
        );

    \I__5875\ : InMux
    port map (
            O => \N__23832\,
            I => \N__23810\
        );

    \I__5874\ : InMux
    port map (
            O => \N__23831\,
            I => \N__23804\
        );

    \I__5873\ : InMux
    port map (
            O => \N__23830\,
            I => \N__23804\
        );

    \I__5872\ : InMux
    port map (
            O => \N__23829\,
            I => \N__23801\
        );

    \I__5871\ : LocalMux
    port map (
            O => \N__23824\,
            I => \N__23798\
        );

    \I__5870\ : InMux
    port map (
            O => \N__23823\,
            I => \N__23793\
        );

    \I__5869\ : InMux
    port map (
            O => \N__23822\,
            I => \N__23793\
        );

    \I__5868\ : InMux
    port map (
            O => \N__23821\,
            I => \N__23790\
        );

    \I__5867\ : InMux
    port map (
            O => \N__23820\,
            I => \N__23787\
        );

    \I__5866\ : LocalMux
    port map (
            O => \N__23815\,
            I => \N__23782\
        );

    \I__5865\ : LocalMux
    port map (
            O => \N__23810\,
            I => \N__23782\
        );

    \I__5864\ : InMux
    port map (
            O => \N__23809\,
            I => \N__23779\
        );

    \I__5863\ : LocalMux
    port map (
            O => \N__23804\,
            I => \b2v_inst1.r_Clk_CountZ0Z_2\
        );

    \I__5862\ : LocalMux
    port map (
            O => \N__23801\,
            I => \b2v_inst1.r_Clk_CountZ0Z_2\
        );

    \I__5861\ : Odrv4
    port map (
            O => \N__23798\,
            I => \b2v_inst1.r_Clk_CountZ0Z_2\
        );

    \I__5860\ : LocalMux
    port map (
            O => \N__23793\,
            I => \b2v_inst1.r_Clk_CountZ0Z_2\
        );

    \I__5859\ : LocalMux
    port map (
            O => \N__23790\,
            I => \b2v_inst1.r_Clk_CountZ0Z_2\
        );

    \I__5858\ : LocalMux
    port map (
            O => \N__23787\,
            I => \b2v_inst1.r_Clk_CountZ0Z_2\
        );

    \I__5857\ : Odrv4
    port map (
            O => \N__23782\,
            I => \b2v_inst1.r_Clk_CountZ0Z_2\
        );

    \I__5856\ : LocalMux
    port map (
            O => \N__23779\,
            I => \b2v_inst1.r_Clk_CountZ0Z_2\
        );

    \I__5855\ : InMux
    port map (
            O => \N__23762\,
            I => \N__23759\
        );

    \I__5854\ : LocalMux
    port map (
            O => \N__23759\,
            I => \b2v_inst1.g2_1_4\
        );

    \I__5853\ : CascadeMux
    port map (
            O => \N__23756\,
            I => \N__23750\
        );

    \I__5852\ : InMux
    port map (
            O => \N__23755\,
            I => \N__23743\
        );

    \I__5851\ : InMux
    port map (
            O => \N__23754\,
            I => \N__23743\
        );

    \I__5850\ : InMux
    port map (
            O => \N__23753\,
            I => \N__23735\
        );

    \I__5849\ : InMux
    port map (
            O => \N__23750\,
            I => \N__23730\
        );

    \I__5848\ : InMux
    port map (
            O => \N__23749\,
            I => \N__23730\
        );

    \I__5847\ : CascadeMux
    port map (
            O => \N__23748\,
            I => \N__23724\
        );

    \I__5846\ : LocalMux
    port map (
            O => \N__23743\,
            I => \N__23721\
        );

    \I__5845\ : CascadeMux
    port map (
            O => \N__23742\,
            I => \N__23718\
        );

    \I__5844\ : InMux
    port map (
            O => \N__23741\,
            I => \N__23715\
        );

    \I__5843\ : InMux
    port map (
            O => \N__23740\,
            I => \N__23712\
        );

    \I__5842\ : InMux
    port map (
            O => \N__23739\,
            I => \N__23709\
        );

    \I__5841\ : InMux
    port map (
            O => \N__23738\,
            I => \N__23700\
        );

    \I__5840\ : LocalMux
    port map (
            O => \N__23735\,
            I => \N__23695\
        );

    \I__5839\ : LocalMux
    port map (
            O => \N__23730\,
            I => \N__23695\
        );

    \I__5838\ : InMux
    port map (
            O => \N__23729\,
            I => \N__23690\
        );

    \I__5837\ : InMux
    port map (
            O => \N__23728\,
            I => \N__23690\
        );

    \I__5836\ : InMux
    port map (
            O => \N__23727\,
            I => \N__23685\
        );

    \I__5835\ : InMux
    port map (
            O => \N__23724\,
            I => \N__23685\
        );

    \I__5834\ : Span4Mux_h
    port map (
            O => \N__23721\,
            I => \N__23682\
        );

    \I__5833\ : InMux
    port map (
            O => \N__23718\,
            I => \N__23679\
        );

    \I__5832\ : LocalMux
    port map (
            O => \N__23715\,
            I => \N__23672\
        );

    \I__5831\ : LocalMux
    port map (
            O => \N__23712\,
            I => \N__23672\
        );

    \I__5830\ : LocalMux
    port map (
            O => \N__23709\,
            I => \N__23672\
        );

    \I__5829\ : InMux
    port map (
            O => \N__23708\,
            I => \N__23667\
        );

    \I__5828\ : InMux
    port map (
            O => \N__23707\,
            I => \N__23667\
        );

    \I__5827\ : InMux
    port map (
            O => \N__23706\,
            I => \N__23664\
        );

    \I__5826\ : InMux
    port map (
            O => \N__23705\,
            I => \N__23661\
        );

    \I__5825\ : InMux
    port map (
            O => \N__23704\,
            I => \N__23656\
        );

    \I__5824\ : InMux
    port map (
            O => \N__23703\,
            I => \N__23656\
        );

    \I__5823\ : LocalMux
    port map (
            O => \N__23700\,
            I => \N__23647\
        );

    \I__5822\ : Span4Mux_h
    port map (
            O => \N__23695\,
            I => \N__23647\
        );

    \I__5821\ : LocalMux
    port map (
            O => \N__23690\,
            I => \N__23647\
        );

    \I__5820\ : LocalMux
    port map (
            O => \N__23685\,
            I => \N__23647\
        );

    \I__5819\ : Odrv4
    port map (
            O => \N__23682\,
            I => \b2v_inst1.r_SM_MainZ0Z_0\
        );

    \I__5818\ : LocalMux
    port map (
            O => \N__23679\,
            I => \b2v_inst1.r_SM_MainZ0Z_0\
        );

    \I__5817\ : Odrv4
    port map (
            O => \N__23672\,
            I => \b2v_inst1.r_SM_MainZ0Z_0\
        );

    \I__5816\ : LocalMux
    port map (
            O => \N__23667\,
            I => \b2v_inst1.r_SM_MainZ0Z_0\
        );

    \I__5815\ : LocalMux
    port map (
            O => \N__23664\,
            I => \b2v_inst1.r_SM_MainZ0Z_0\
        );

    \I__5814\ : LocalMux
    port map (
            O => \N__23661\,
            I => \b2v_inst1.r_SM_MainZ0Z_0\
        );

    \I__5813\ : LocalMux
    port map (
            O => \N__23656\,
            I => \b2v_inst1.r_SM_MainZ0Z_0\
        );

    \I__5812\ : Odrv4
    port map (
            O => \N__23647\,
            I => \b2v_inst1.r_SM_MainZ0Z_0\
        );

    \I__5811\ : InMux
    port map (
            O => \N__23630\,
            I => \N__23626\
        );

    \I__5810\ : InMux
    port map (
            O => \N__23629\,
            I => \N__23614\
        );

    \I__5809\ : LocalMux
    port map (
            O => \N__23626\,
            I => \N__23609\
        );

    \I__5808\ : CascadeMux
    port map (
            O => \N__23625\,
            I => \N__23604\
        );

    \I__5807\ : InMux
    port map (
            O => \N__23624\,
            I => \N__23600\
        );

    \I__5806\ : CascadeMux
    port map (
            O => \N__23623\,
            I => \N__23595\
        );

    \I__5805\ : InMux
    port map (
            O => \N__23622\,
            I => \N__23583\
        );

    \I__5804\ : InMux
    port map (
            O => \N__23621\,
            I => \N__23583\
        );

    \I__5803\ : InMux
    port map (
            O => \N__23620\,
            I => \N__23574\
        );

    \I__5802\ : InMux
    port map (
            O => \N__23619\,
            I => \N__23574\
        );

    \I__5801\ : InMux
    port map (
            O => \N__23618\,
            I => \N__23574\
        );

    \I__5800\ : InMux
    port map (
            O => \N__23617\,
            I => \N__23574\
        );

    \I__5799\ : LocalMux
    port map (
            O => \N__23614\,
            I => \N__23571\
        );

    \I__5798\ : InMux
    port map (
            O => \N__23613\,
            I => \N__23566\
        );

    \I__5797\ : InMux
    port map (
            O => \N__23612\,
            I => \N__23566\
        );

    \I__5796\ : Span4Mux_v
    port map (
            O => \N__23609\,
            I => \N__23563\
        );

    \I__5795\ : InMux
    port map (
            O => \N__23608\,
            I => \N__23558\
        );

    \I__5794\ : InMux
    port map (
            O => \N__23607\,
            I => \N__23558\
        );

    \I__5793\ : InMux
    port map (
            O => \N__23604\,
            I => \N__23553\
        );

    \I__5792\ : InMux
    port map (
            O => \N__23603\,
            I => \N__23553\
        );

    \I__5791\ : LocalMux
    port map (
            O => \N__23600\,
            I => \N__23550\
        );

    \I__5790\ : InMux
    port map (
            O => \N__23599\,
            I => \N__23545\
        );

    \I__5789\ : InMux
    port map (
            O => \N__23598\,
            I => \N__23545\
        );

    \I__5788\ : InMux
    port map (
            O => \N__23595\,
            I => \N__23540\
        );

    \I__5787\ : InMux
    port map (
            O => \N__23594\,
            I => \N__23540\
        );

    \I__5786\ : InMux
    port map (
            O => \N__23593\,
            I => \N__23533\
        );

    \I__5785\ : InMux
    port map (
            O => \N__23592\,
            I => \N__23533\
        );

    \I__5784\ : InMux
    port map (
            O => \N__23591\,
            I => \N__23533\
        );

    \I__5783\ : InMux
    port map (
            O => \N__23590\,
            I => \N__23526\
        );

    \I__5782\ : InMux
    port map (
            O => \N__23589\,
            I => \N__23526\
        );

    \I__5781\ : InMux
    port map (
            O => \N__23588\,
            I => \N__23526\
        );

    \I__5780\ : LocalMux
    port map (
            O => \N__23583\,
            I => \N__23519\
        );

    \I__5779\ : LocalMux
    port map (
            O => \N__23574\,
            I => \N__23519\
        );

    \I__5778\ : Span4Mux_h
    port map (
            O => \N__23571\,
            I => \N__23519\
        );

    \I__5777\ : LocalMux
    port map (
            O => \N__23566\,
            I => \b2v_inst1.r_SM_MainZ0Z_1\
        );

    \I__5776\ : Odrv4
    port map (
            O => \N__23563\,
            I => \b2v_inst1.r_SM_MainZ0Z_1\
        );

    \I__5775\ : LocalMux
    port map (
            O => \N__23558\,
            I => \b2v_inst1.r_SM_MainZ0Z_1\
        );

    \I__5774\ : LocalMux
    port map (
            O => \N__23553\,
            I => \b2v_inst1.r_SM_MainZ0Z_1\
        );

    \I__5773\ : Odrv4
    port map (
            O => \N__23550\,
            I => \b2v_inst1.r_SM_MainZ0Z_1\
        );

    \I__5772\ : LocalMux
    port map (
            O => \N__23545\,
            I => \b2v_inst1.r_SM_MainZ0Z_1\
        );

    \I__5771\ : LocalMux
    port map (
            O => \N__23540\,
            I => \b2v_inst1.r_SM_MainZ0Z_1\
        );

    \I__5770\ : LocalMux
    port map (
            O => \N__23533\,
            I => \b2v_inst1.r_SM_MainZ0Z_1\
        );

    \I__5769\ : LocalMux
    port map (
            O => \N__23526\,
            I => \b2v_inst1.r_SM_MainZ0Z_1\
        );

    \I__5768\ : Odrv4
    port map (
            O => \N__23519\,
            I => \b2v_inst1.r_SM_MainZ0Z_1\
        );

    \I__5767\ : CascadeMux
    port map (
            O => \N__23498\,
            I => \N__23491\
        );

    \I__5766\ : InMux
    port map (
            O => \N__23497\,
            I => \N__23485\
        );

    \I__5765\ : CascadeMux
    port map (
            O => \N__23496\,
            I => \N__23479\
        );

    \I__5764\ : CascadeMux
    port map (
            O => \N__23495\,
            I => \N__23476\
        );

    \I__5763\ : InMux
    port map (
            O => \N__23494\,
            I => \N__23471\
        );

    \I__5762\ : InMux
    port map (
            O => \N__23491\,
            I => \N__23468\
        );

    \I__5761\ : InMux
    port map (
            O => \N__23490\,
            I => \N__23465\
        );

    \I__5760\ : InMux
    port map (
            O => \N__23489\,
            I => \N__23462\
        );

    \I__5759\ : InMux
    port map (
            O => \N__23488\,
            I => \N__23459\
        );

    \I__5758\ : LocalMux
    port map (
            O => \N__23485\,
            I => \N__23456\
        );

    \I__5757\ : CascadeMux
    port map (
            O => \N__23484\,
            I => \N__23452\
        );

    \I__5756\ : InMux
    port map (
            O => \N__23483\,
            I => \N__23449\
        );

    \I__5755\ : InMux
    port map (
            O => \N__23482\,
            I => \N__23446\
        );

    \I__5754\ : InMux
    port map (
            O => \N__23479\,
            I => \N__23442\
        );

    \I__5753\ : InMux
    port map (
            O => \N__23476\,
            I => \N__23439\
        );

    \I__5752\ : CascadeMux
    port map (
            O => \N__23475\,
            I => \N__23436\
        );

    \I__5751\ : CascadeMux
    port map (
            O => \N__23474\,
            I => \N__23433\
        );

    \I__5750\ : LocalMux
    port map (
            O => \N__23471\,
            I => \N__23430\
        );

    \I__5749\ : LocalMux
    port map (
            O => \N__23468\,
            I => \N__23427\
        );

    \I__5748\ : LocalMux
    port map (
            O => \N__23465\,
            I => \N__23420\
        );

    \I__5747\ : LocalMux
    port map (
            O => \N__23462\,
            I => \N__23420\
        );

    \I__5746\ : LocalMux
    port map (
            O => \N__23459\,
            I => \N__23420\
        );

    \I__5745\ : Span4Mux_v
    port map (
            O => \N__23456\,
            I => \N__23417\
        );

    \I__5744\ : InMux
    port map (
            O => \N__23455\,
            I => \N__23412\
        );

    \I__5743\ : InMux
    port map (
            O => \N__23452\,
            I => \N__23412\
        );

    \I__5742\ : LocalMux
    port map (
            O => \N__23449\,
            I => \N__23409\
        );

    \I__5741\ : LocalMux
    port map (
            O => \N__23446\,
            I => \N__23406\
        );

    \I__5740\ : InMux
    port map (
            O => \N__23445\,
            I => \N__23403\
        );

    \I__5739\ : LocalMux
    port map (
            O => \N__23442\,
            I => \N__23398\
        );

    \I__5738\ : LocalMux
    port map (
            O => \N__23439\,
            I => \N__23398\
        );

    \I__5737\ : InMux
    port map (
            O => \N__23436\,
            I => \N__23395\
        );

    \I__5736\ : InMux
    port map (
            O => \N__23433\,
            I => \N__23392\
        );

    \I__5735\ : Span4Mux_v
    port map (
            O => \N__23430\,
            I => \N__23379\
        );

    \I__5734\ : Span4Mux_v
    port map (
            O => \N__23427\,
            I => \N__23379\
        );

    \I__5733\ : Span4Mux_v
    port map (
            O => \N__23420\,
            I => \N__23379\
        );

    \I__5732\ : Span4Mux_h
    port map (
            O => \N__23417\,
            I => \N__23379\
        );

    \I__5731\ : LocalMux
    port map (
            O => \N__23412\,
            I => \N__23379\
        );

    \I__5730\ : Span4Mux_v
    port map (
            O => \N__23409\,
            I => \N__23379\
        );

    \I__5729\ : Odrv4
    port map (
            O => \N__23406\,
            I => \b2v_inst1.r_SM_MainZ0Z_2\
        );

    \I__5728\ : LocalMux
    port map (
            O => \N__23403\,
            I => \b2v_inst1.r_SM_MainZ0Z_2\
        );

    \I__5727\ : Odrv4
    port map (
            O => \N__23398\,
            I => \b2v_inst1.r_SM_MainZ0Z_2\
        );

    \I__5726\ : LocalMux
    port map (
            O => \N__23395\,
            I => \b2v_inst1.r_SM_MainZ0Z_2\
        );

    \I__5725\ : LocalMux
    port map (
            O => \N__23392\,
            I => \b2v_inst1.r_SM_MainZ0Z_2\
        );

    \I__5724\ : Odrv4
    port map (
            O => \N__23379\,
            I => \b2v_inst1.r_SM_MainZ0Z_2\
        );

    \I__5723\ : InMux
    port map (
            O => \N__23366\,
            I => \N__23362\
        );

    \I__5722\ : InMux
    port map (
            O => \N__23365\,
            I => \N__23359\
        );

    \I__5721\ : LocalMux
    port map (
            O => \N__23362\,
            I => \b2v_inst1.N_11_1\
        );

    \I__5720\ : LocalMux
    port map (
            O => \N__23359\,
            I => \b2v_inst1.N_11_1\
        );

    \I__5719\ : CascadeMux
    port map (
            O => \N__23354\,
            I => \b2v_inst1.g0_0_i_a6_2_0_cascade_\
        );

    \I__5718\ : CascadeMux
    port map (
            O => \N__23351\,
            I => \N__23348\
        );

    \I__5717\ : InMux
    port map (
            O => \N__23348\,
            I => \N__23336\
        );

    \I__5716\ : InMux
    port map (
            O => \N__23347\,
            I => \N__23336\
        );

    \I__5715\ : CascadeMux
    port map (
            O => \N__23346\,
            I => \N__23333\
        );

    \I__5714\ : CascadeMux
    port map (
            O => \N__23345\,
            I => \N__23330\
        );

    \I__5713\ : CascadeMux
    port map (
            O => \N__23344\,
            I => \N__23327\
        );

    \I__5712\ : InMux
    port map (
            O => \N__23343\,
            I => \N__23324\
        );

    \I__5711\ : InMux
    port map (
            O => \N__23342\,
            I => \N__23321\
        );

    \I__5710\ : CascadeMux
    port map (
            O => \N__23341\,
            I => \N__23317\
        );

    \I__5709\ : LocalMux
    port map (
            O => \N__23336\,
            I => \N__23310\
        );

    \I__5708\ : InMux
    port map (
            O => \N__23333\,
            I => \N__23305\
        );

    \I__5707\ : InMux
    port map (
            O => \N__23330\,
            I => \N__23305\
        );

    \I__5706\ : InMux
    port map (
            O => \N__23327\,
            I => \N__23302\
        );

    \I__5705\ : LocalMux
    port map (
            O => \N__23324\,
            I => \N__23296\
        );

    \I__5704\ : LocalMux
    port map (
            O => \N__23321\,
            I => \N__23296\
        );

    \I__5703\ : CascadeMux
    port map (
            O => \N__23320\,
            I => \N__23291\
        );

    \I__5702\ : InMux
    port map (
            O => \N__23317\,
            I => \N__23286\
        );

    \I__5701\ : InMux
    port map (
            O => \N__23316\,
            I => \N__23286\
        );

    \I__5700\ : InMux
    port map (
            O => \N__23315\,
            I => \N__23282\
        );

    \I__5699\ : InMux
    port map (
            O => \N__23314\,
            I => \N__23279\
        );

    \I__5698\ : InMux
    port map (
            O => \N__23313\,
            I => \N__23276\
        );

    \I__5697\ : Span4Mux_v
    port map (
            O => \N__23310\,
            I => \N__23271\
        );

    \I__5696\ : LocalMux
    port map (
            O => \N__23305\,
            I => \N__23271\
        );

    \I__5695\ : LocalMux
    port map (
            O => \N__23302\,
            I => \N__23268\
        );

    \I__5694\ : InMux
    port map (
            O => \N__23301\,
            I => \N__23265\
        );

    \I__5693\ : Span4Mux_h
    port map (
            O => \N__23296\,
            I => \N__23262\
        );

    \I__5692\ : InMux
    port map (
            O => \N__23295\,
            I => \N__23255\
        );

    \I__5691\ : InMux
    port map (
            O => \N__23294\,
            I => \N__23255\
        );

    \I__5690\ : InMux
    port map (
            O => \N__23291\,
            I => \N__23255\
        );

    \I__5689\ : LocalMux
    port map (
            O => \N__23286\,
            I => \N__23252\
        );

    \I__5688\ : InMux
    port map (
            O => \N__23285\,
            I => \N__23249\
        );

    \I__5687\ : LocalMux
    port map (
            O => \N__23282\,
            I => \N__23238\
        );

    \I__5686\ : LocalMux
    port map (
            O => \N__23279\,
            I => \N__23238\
        );

    \I__5685\ : LocalMux
    port map (
            O => \N__23276\,
            I => \N__23238\
        );

    \I__5684\ : Span4Mux_h
    port map (
            O => \N__23271\,
            I => \N__23238\
        );

    \I__5683\ : Span4Mux_h
    port map (
            O => \N__23268\,
            I => \N__23238\
        );

    \I__5682\ : LocalMux
    port map (
            O => \N__23265\,
            I => \b2v_inst1.r_Clk_CountZ0Z_4\
        );

    \I__5681\ : Odrv4
    port map (
            O => \N__23262\,
            I => \b2v_inst1.r_Clk_CountZ0Z_4\
        );

    \I__5680\ : LocalMux
    port map (
            O => \N__23255\,
            I => \b2v_inst1.r_Clk_CountZ0Z_4\
        );

    \I__5679\ : Odrv4
    port map (
            O => \N__23252\,
            I => \b2v_inst1.r_Clk_CountZ0Z_4\
        );

    \I__5678\ : LocalMux
    port map (
            O => \N__23249\,
            I => \b2v_inst1.r_Clk_CountZ0Z_4\
        );

    \I__5677\ : Odrv4
    port map (
            O => \N__23238\,
            I => \b2v_inst1.r_Clk_CountZ0Z_4\
        );

    \I__5676\ : InMux
    port map (
            O => \N__23225\,
            I => \N__23222\
        );

    \I__5675\ : LocalMux
    port map (
            O => \N__23222\,
            I => \b2v_inst1.g0_0_i_0_0\
        );

    \I__5674\ : CascadeMux
    port map (
            O => \N__23219\,
            I => \N__23212\
        );

    \I__5673\ : InMux
    port map (
            O => \N__23218\,
            I => \N__23207\
        );

    \I__5672\ : CascadeMux
    port map (
            O => \N__23217\,
            I => \N__23203\
        );

    \I__5671\ : CascadeMux
    port map (
            O => \N__23216\,
            I => \N__23196\
        );

    \I__5670\ : CascadeMux
    port map (
            O => \N__23215\,
            I => \N__23192\
        );

    \I__5669\ : InMux
    port map (
            O => \N__23212\,
            I => \N__23185\
        );

    \I__5668\ : InMux
    port map (
            O => \N__23211\,
            I => \N__23185\
        );

    \I__5667\ : InMux
    port map (
            O => \N__23210\,
            I => \N__23185\
        );

    \I__5666\ : LocalMux
    port map (
            O => \N__23207\,
            I => \N__23182\
        );

    \I__5665\ : InMux
    port map (
            O => \N__23206\,
            I => \N__23177\
        );

    \I__5664\ : InMux
    port map (
            O => \N__23203\,
            I => \N__23177\
        );

    \I__5663\ : InMux
    port map (
            O => \N__23202\,
            I => \N__23168\
        );

    \I__5662\ : InMux
    port map (
            O => \N__23201\,
            I => \N__23168\
        );

    \I__5661\ : InMux
    port map (
            O => \N__23200\,
            I => \N__23163\
        );

    \I__5660\ : InMux
    port map (
            O => \N__23199\,
            I => \N__23158\
        );

    \I__5659\ : InMux
    port map (
            O => \N__23196\,
            I => \N__23158\
        );

    \I__5658\ : InMux
    port map (
            O => \N__23195\,
            I => \N__23153\
        );

    \I__5657\ : InMux
    port map (
            O => \N__23192\,
            I => \N__23153\
        );

    \I__5656\ : LocalMux
    port map (
            O => \N__23185\,
            I => \N__23149\
        );

    \I__5655\ : Span4Mux_v
    port map (
            O => \N__23182\,
            I => \N__23144\
        );

    \I__5654\ : LocalMux
    port map (
            O => \N__23177\,
            I => \N__23144\
        );

    \I__5653\ : InMux
    port map (
            O => \N__23176\,
            I => \N__23135\
        );

    \I__5652\ : InMux
    port map (
            O => \N__23175\,
            I => \N__23135\
        );

    \I__5651\ : InMux
    port map (
            O => \N__23174\,
            I => \N__23135\
        );

    \I__5650\ : InMux
    port map (
            O => \N__23173\,
            I => \N__23135\
        );

    \I__5649\ : LocalMux
    port map (
            O => \N__23168\,
            I => \N__23131\
        );

    \I__5648\ : InMux
    port map (
            O => \N__23167\,
            I => \N__23126\
        );

    \I__5647\ : InMux
    port map (
            O => \N__23166\,
            I => \N__23126\
        );

    \I__5646\ : LocalMux
    port map (
            O => \N__23163\,
            I => \N__23119\
        );

    \I__5645\ : LocalMux
    port map (
            O => \N__23158\,
            I => \N__23119\
        );

    \I__5644\ : LocalMux
    port map (
            O => \N__23153\,
            I => \N__23119\
        );

    \I__5643\ : InMux
    port map (
            O => \N__23152\,
            I => \N__23116\
        );

    \I__5642\ : Span12Mux_v
    port map (
            O => \N__23149\,
            I => \N__23113\
        );

    \I__5641\ : Span4Mux_h
    port map (
            O => \N__23144\,
            I => \N__23110\
        );

    \I__5640\ : LocalMux
    port map (
            O => \N__23135\,
            I => \N__23107\
        );

    \I__5639\ : InMux
    port map (
            O => \N__23134\,
            I => \N__23104\
        );

    \I__5638\ : Span4Mux_v
    port map (
            O => \N__23131\,
            I => \N__23097\
        );

    \I__5637\ : LocalMux
    port map (
            O => \N__23126\,
            I => \N__23097\
        );

    \I__5636\ : Span4Mux_h
    port map (
            O => \N__23119\,
            I => \N__23097\
        );

    \I__5635\ : LocalMux
    port map (
            O => \N__23116\,
            I => \b2v_inst.indiceZ0Z_0\
        );

    \I__5634\ : Odrv12
    port map (
            O => \N__23113\,
            I => \b2v_inst.indiceZ0Z_0\
        );

    \I__5633\ : Odrv4
    port map (
            O => \N__23110\,
            I => \b2v_inst.indiceZ0Z_0\
        );

    \I__5632\ : Odrv12
    port map (
            O => \N__23107\,
            I => \b2v_inst.indiceZ0Z_0\
        );

    \I__5631\ : LocalMux
    port map (
            O => \N__23104\,
            I => \b2v_inst.indiceZ0Z_0\
        );

    \I__5630\ : Odrv4
    port map (
            O => \N__23097\,
            I => \b2v_inst.indiceZ0Z_0\
        );

    \I__5629\ : InMux
    port map (
            O => \N__23084\,
            I => \N__23078\
        );

    \I__5628\ : InMux
    port map (
            O => \N__23083\,
            I => \N__23071\
        );

    \I__5627\ : InMux
    port map (
            O => \N__23082\,
            I => \N__23071\
        );

    \I__5626\ : InMux
    port map (
            O => \N__23081\,
            I => \N__23068\
        );

    \I__5625\ : LocalMux
    port map (
            O => \N__23078\,
            I => \N__23065\
        );

    \I__5624\ : CascadeMux
    port map (
            O => \N__23077\,
            I => \N__23060\
        );

    \I__5623\ : CascadeMux
    port map (
            O => \N__23076\,
            I => \N__23055\
        );

    \I__5622\ : LocalMux
    port map (
            O => \N__23071\,
            I => \N__23051\
        );

    \I__5621\ : LocalMux
    port map (
            O => \N__23068\,
            I => \N__23048\
        );

    \I__5620\ : Span4Mux_v
    port map (
            O => \N__23065\,
            I => \N__23045\
        );

    \I__5619\ : InMux
    port map (
            O => \N__23064\,
            I => \N__23038\
        );

    \I__5618\ : InMux
    port map (
            O => \N__23063\,
            I => \N__23038\
        );

    \I__5617\ : InMux
    port map (
            O => \N__23060\,
            I => \N__23038\
        );

    \I__5616\ : InMux
    port map (
            O => \N__23059\,
            I => \N__23029\
        );

    \I__5615\ : InMux
    port map (
            O => \N__23058\,
            I => \N__23029\
        );

    \I__5614\ : InMux
    port map (
            O => \N__23055\,
            I => \N__23029\
        );

    \I__5613\ : CascadeMux
    port map (
            O => \N__23054\,
            I => \N__23024\
        );

    \I__5612\ : Span4Mux_v
    port map (
            O => \N__23051\,
            I => \N__23012\
        );

    \I__5611\ : Span4Mux_h
    port map (
            O => \N__23048\,
            I => \N__23012\
        );

    \I__5610\ : Span4Mux_v
    port map (
            O => \N__23045\,
            I => \N__23012\
        );

    \I__5609\ : LocalMux
    port map (
            O => \N__23038\,
            I => \N__23012\
        );

    \I__5608\ : InMux
    port map (
            O => \N__23037\,
            I => \N__23007\
        );

    \I__5607\ : InMux
    port map (
            O => \N__23036\,
            I => \N__23007\
        );

    \I__5606\ : LocalMux
    port map (
            O => \N__23029\,
            I => \N__23004\
        );

    \I__5605\ : InMux
    port map (
            O => \N__23028\,
            I => \N__22997\
        );

    \I__5604\ : InMux
    port map (
            O => \N__23027\,
            I => \N__22997\
        );

    \I__5603\ : InMux
    port map (
            O => \N__23024\,
            I => \N__22997\
        );

    \I__5602\ : InMux
    port map (
            O => \N__23023\,
            I => \N__22991\
        );

    \I__5601\ : InMux
    port map (
            O => \N__23022\,
            I => \N__22991\
        );

    \I__5600\ : InMux
    port map (
            O => \N__23021\,
            I => \N__22988\
        );

    \I__5599\ : Span4Mux_h
    port map (
            O => \N__23012\,
            I => \N__22985\
        );

    \I__5598\ : LocalMux
    port map (
            O => \N__23007\,
            I => \N__22982\
        );

    \I__5597\ : Span4Mux_v
    port map (
            O => \N__23004\,
            I => \N__22977\
        );

    \I__5596\ : LocalMux
    port map (
            O => \N__22997\,
            I => \N__22977\
        );

    \I__5595\ : InMux
    port map (
            O => \N__22996\,
            I => \N__22974\
        );

    \I__5594\ : LocalMux
    port map (
            O => \N__22991\,
            I => \N__22969\
        );

    \I__5593\ : LocalMux
    port map (
            O => \N__22988\,
            I => \N__22969\
        );

    \I__5592\ : Span4Mux_h
    port map (
            O => \N__22985\,
            I => \N__22966\
        );

    \I__5591\ : Span4Mux_v
    port map (
            O => \N__22982\,
            I => \N__22961\
        );

    \I__5590\ : Span4Mux_h
    port map (
            O => \N__22977\,
            I => \N__22961\
        );

    \I__5589\ : LocalMux
    port map (
            O => \N__22974\,
            I => \b2v_inst.indiceZ0Z_1\
        );

    \I__5588\ : Odrv4
    port map (
            O => \N__22969\,
            I => \b2v_inst.indiceZ0Z_1\
        );

    \I__5587\ : Odrv4
    port map (
            O => \N__22966\,
            I => \b2v_inst.indiceZ0Z_1\
        );

    \I__5586\ : Odrv4
    port map (
            O => \N__22961\,
            I => \b2v_inst.indiceZ0Z_1\
        );

    \I__5585\ : CEMux
    port map (
            O => \N__22952\,
            I => \N__22928\
        );

    \I__5584\ : CEMux
    port map (
            O => \N__22951\,
            I => \N__22928\
        );

    \I__5583\ : CEMux
    port map (
            O => \N__22950\,
            I => \N__22928\
        );

    \I__5582\ : CEMux
    port map (
            O => \N__22949\,
            I => \N__22928\
        );

    \I__5581\ : CEMux
    port map (
            O => \N__22948\,
            I => \N__22928\
        );

    \I__5580\ : CEMux
    port map (
            O => \N__22947\,
            I => \N__22928\
        );

    \I__5579\ : CEMux
    port map (
            O => \N__22946\,
            I => \N__22928\
        );

    \I__5578\ : CEMux
    port map (
            O => \N__22945\,
            I => \N__22928\
        );

    \I__5577\ : GlobalMux
    port map (
            O => \N__22928\,
            I => \N__22925\
        );

    \I__5576\ : gio2CtrlBuf
    port map (
            O => \N__22925\,
            I => \b2v_inst.state_g_2\
        );

    \I__5575\ : SRMux
    port map (
            O => \N__22922\,
            I => \N__22778\
        );

    \I__5574\ : SRMux
    port map (
            O => \N__22921\,
            I => \N__22778\
        );

    \I__5573\ : SRMux
    port map (
            O => \N__22920\,
            I => \N__22778\
        );

    \I__5572\ : SRMux
    port map (
            O => \N__22919\,
            I => \N__22778\
        );

    \I__5571\ : SRMux
    port map (
            O => \N__22918\,
            I => \N__22778\
        );

    \I__5570\ : SRMux
    port map (
            O => \N__22917\,
            I => \N__22778\
        );

    \I__5569\ : SRMux
    port map (
            O => \N__22916\,
            I => \N__22778\
        );

    \I__5568\ : SRMux
    port map (
            O => \N__22915\,
            I => \N__22778\
        );

    \I__5567\ : SRMux
    port map (
            O => \N__22914\,
            I => \N__22778\
        );

    \I__5566\ : SRMux
    port map (
            O => \N__22913\,
            I => \N__22778\
        );

    \I__5565\ : SRMux
    port map (
            O => \N__22912\,
            I => \N__22778\
        );

    \I__5564\ : SRMux
    port map (
            O => \N__22911\,
            I => \N__22778\
        );

    \I__5563\ : SRMux
    port map (
            O => \N__22910\,
            I => \N__22778\
        );

    \I__5562\ : SRMux
    port map (
            O => \N__22909\,
            I => \N__22778\
        );

    \I__5561\ : SRMux
    port map (
            O => \N__22908\,
            I => \N__22778\
        );

    \I__5560\ : SRMux
    port map (
            O => \N__22907\,
            I => \N__22778\
        );

    \I__5559\ : SRMux
    port map (
            O => \N__22906\,
            I => \N__22778\
        );

    \I__5558\ : SRMux
    port map (
            O => \N__22905\,
            I => \N__22778\
        );

    \I__5557\ : SRMux
    port map (
            O => \N__22904\,
            I => \N__22778\
        );

    \I__5556\ : SRMux
    port map (
            O => \N__22903\,
            I => \N__22778\
        );

    \I__5555\ : SRMux
    port map (
            O => \N__22902\,
            I => \N__22778\
        );

    \I__5554\ : SRMux
    port map (
            O => \N__22901\,
            I => \N__22778\
        );

    \I__5553\ : SRMux
    port map (
            O => \N__22900\,
            I => \N__22778\
        );

    \I__5552\ : SRMux
    port map (
            O => \N__22899\,
            I => \N__22778\
        );

    \I__5551\ : SRMux
    port map (
            O => \N__22898\,
            I => \N__22778\
        );

    \I__5550\ : SRMux
    port map (
            O => \N__22897\,
            I => \N__22778\
        );

    \I__5549\ : SRMux
    port map (
            O => \N__22896\,
            I => \N__22778\
        );

    \I__5548\ : SRMux
    port map (
            O => \N__22895\,
            I => \N__22778\
        );

    \I__5547\ : SRMux
    port map (
            O => \N__22894\,
            I => \N__22778\
        );

    \I__5546\ : SRMux
    port map (
            O => \N__22893\,
            I => \N__22778\
        );

    \I__5545\ : SRMux
    port map (
            O => \N__22892\,
            I => \N__22778\
        );

    \I__5544\ : SRMux
    port map (
            O => \N__22891\,
            I => \N__22778\
        );

    \I__5543\ : SRMux
    port map (
            O => \N__22890\,
            I => \N__22778\
        );

    \I__5542\ : SRMux
    port map (
            O => \N__22889\,
            I => \N__22778\
        );

    \I__5541\ : SRMux
    port map (
            O => \N__22888\,
            I => \N__22778\
        );

    \I__5540\ : SRMux
    port map (
            O => \N__22887\,
            I => \N__22778\
        );

    \I__5539\ : SRMux
    port map (
            O => \N__22886\,
            I => \N__22778\
        );

    \I__5538\ : SRMux
    port map (
            O => \N__22885\,
            I => \N__22778\
        );

    \I__5537\ : SRMux
    port map (
            O => \N__22884\,
            I => \N__22778\
        );

    \I__5536\ : SRMux
    port map (
            O => \N__22883\,
            I => \N__22778\
        );

    \I__5535\ : SRMux
    port map (
            O => \N__22882\,
            I => \N__22778\
        );

    \I__5534\ : SRMux
    port map (
            O => \N__22881\,
            I => \N__22778\
        );

    \I__5533\ : SRMux
    port map (
            O => \N__22880\,
            I => \N__22778\
        );

    \I__5532\ : SRMux
    port map (
            O => \N__22879\,
            I => \N__22778\
        );

    \I__5531\ : SRMux
    port map (
            O => \N__22878\,
            I => \N__22778\
        );

    \I__5530\ : SRMux
    port map (
            O => \N__22877\,
            I => \N__22778\
        );

    \I__5529\ : SRMux
    port map (
            O => \N__22876\,
            I => \N__22778\
        );

    \I__5528\ : SRMux
    port map (
            O => \N__22875\,
            I => \N__22778\
        );

    \I__5527\ : GlobalMux
    port map (
            O => \N__22778\,
            I => \N__22775\
        );

    \I__5526\ : gio2CtrlBuf
    port map (
            O => \N__22775\,
            I => reset_i_g
        );

    \I__5525\ : InMux
    port map (
            O => \N__22772\,
            I => \N__22769\
        );

    \I__5524\ : LocalMux
    port map (
            O => \N__22769\,
            I => \N__22766\
        );

    \I__5523\ : Span4Mux_h
    port map (
            O => \N__22766\,
            I => \N__22763\
        );

    \I__5522\ : Span4Mux_v
    port map (
            O => \N__22763\,
            I => \N__22760\
        );

    \I__5521\ : Odrv4
    port map (
            O => \N__22760\,
            I => uart_rx_i
        );

    \I__5520\ : InMux
    port map (
            O => \N__22757\,
            I => \N__22754\
        );

    \I__5519\ : LocalMux
    port map (
            O => \N__22754\,
            I => \b2v_inst1.r_RX_Data_RZ0\
        );

    \I__5518\ : CascadeMux
    port map (
            O => \N__22751\,
            I => \N__22743\
        );

    \I__5517\ : CascadeMux
    port map (
            O => \N__22750\,
            I => \N__22740\
        );

    \I__5516\ : CascadeMux
    port map (
            O => \N__22749\,
            I => \N__22737\
        );

    \I__5515\ : CascadeMux
    port map (
            O => \N__22748\,
            I => \N__22734\
        );

    \I__5514\ : CascadeMux
    port map (
            O => \N__22747\,
            I => \N__22730\
        );

    \I__5513\ : CascadeMux
    port map (
            O => \N__22746\,
            I => \N__22727\
        );

    \I__5512\ : InMux
    port map (
            O => \N__22743\,
            I => \N__22724\
        );

    \I__5511\ : InMux
    port map (
            O => \N__22740\,
            I => \N__22715\
        );

    \I__5510\ : InMux
    port map (
            O => \N__22737\,
            I => \N__22715\
        );

    \I__5509\ : InMux
    port map (
            O => \N__22734\,
            I => \N__22715\
        );

    \I__5508\ : InMux
    port map (
            O => \N__22733\,
            I => \N__22715\
        );

    \I__5507\ : InMux
    port map (
            O => \N__22730\,
            I => \N__22710\
        );

    \I__5506\ : InMux
    port map (
            O => \N__22727\,
            I => \N__22710\
        );

    \I__5505\ : LocalMux
    port map (
            O => \N__22724\,
            I => \N__22705\
        );

    \I__5504\ : LocalMux
    port map (
            O => \N__22715\,
            I => \N__22700\
        );

    \I__5503\ : LocalMux
    port map (
            O => \N__22710\,
            I => \N__22700\
        );

    \I__5502\ : CascadeMux
    port map (
            O => \N__22709\,
            I => \N__22695\
        );

    \I__5501\ : InMux
    port map (
            O => \N__22708\,
            I => \N__22691\
        );

    \I__5500\ : Span4Mux_h
    port map (
            O => \N__22705\,
            I => \N__22686\
        );

    \I__5499\ : Span4Mux_v
    port map (
            O => \N__22700\,
            I => \N__22683\
        );

    \I__5498\ : CascadeMux
    port map (
            O => \N__22699\,
            I => \N__22680\
        );

    \I__5497\ : CascadeMux
    port map (
            O => \N__22698\,
            I => \N__22676\
        );

    \I__5496\ : InMux
    port map (
            O => \N__22695\,
            I => \N__22673\
        );

    \I__5495\ : InMux
    port map (
            O => \N__22694\,
            I => \N__22670\
        );

    \I__5494\ : LocalMux
    port map (
            O => \N__22691\,
            I => \N__22667\
        );

    \I__5493\ : InMux
    port map (
            O => \N__22690\,
            I => \N__22664\
        );

    \I__5492\ : CascadeMux
    port map (
            O => \N__22689\,
            I => \N__22661\
        );

    \I__5491\ : Span4Mux_h
    port map (
            O => \N__22686\,
            I => \N__22658\
        );

    \I__5490\ : Span4Mux_v
    port map (
            O => \N__22683\,
            I => \N__22655\
        );

    \I__5489\ : InMux
    port map (
            O => \N__22680\,
            I => \N__22650\
        );

    \I__5488\ : InMux
    port map (
            O => \N__22679\,
            I => \N__22650\
        );

    \I__5487\ : InMux
    port map (
            O => \N__22676\,
            I => \N__22647\
        );

    \I__5486\ : LocalMux
    port map (
            O => \N__22673\,
            I => \N__22642\
        );

    \I__5485\ : LocalMux
    port map (
            O => \N__22670\,
            I => \N__22642\
        );

    \I__5484\ : Span4Mux_v
    port map (
            O => \N__22667\,
            I => \N__22637\
        );

    \I__5483\ : LocalMux
    port map (
            O => \N__22664\,
            I => \N__22637\
        );

    \I__5482\ : InMux
    port map (
            O => \N__22661\,
            I => \N__22634\
        );

    \I__5481\ : Span4Mux_h
    port map (
            O => \N__22658\,
            I => \N__22631\
        );

    \I__5480\ : Span4Mux_h
    port map (
            O => \N__22655\,
            I => \N__22624\
        );

    \I__5479\ : LocalMux
    port map (
            O => \N__22650\,
            I => \N__22624\
        );

    \I__5478\ : LocalMux
    port map (
            O => \N__22647\,
            I => \N__22624\
        );

    \I__5477\ : Span4Mux_h
    port map (
            O => \N__22642\,
            I => \N__22621\
        );

    \I__5476\ : Span4Mux_h
    port map (
            O => \N__22637\,
            I => \N__22618\
        );

    \I__5475\ : LocalMux
    port map (
            O => \N__22634\,
            I => \b2v_inst1.r_RX_DataZ0\
        );

    \I__5474\ : Odrv4
    port map (
            O => \N__22631\,
            I => \b2v_inst1.r_RX_DataZ0\
        );

    \I__5473\ : Odrv4
    port map (
            O => \N__22624\,
            I => \b2v_inst1.r_RX_DataZ0\
        );

    \I__5472\ : Odrv4
    port map (
            O => \N__22621\,
            I => \b2v_inst1.r_RX_DataZ0\
        );

    \I__5471\ : Odrv4
    port map (
            O => \N__22618\,
            I => \b2v_inst1.r_RX_DataZ0\
        );

    \I__5470\ : ClkMux
    port map (
            O => \N__22607\,
            I => \N__22602\
        );

    \I__5469\ : ClkMux
    port map (
            O => \N__22606\,
            I => \N__22599\
        );

    \I__5468\ : ClkMux
    port map (
            O => \N__22605\,
            I => \N__22590\
        );

    \I__5467\ : LocalMux
    port map (
            O => \N__22602\,
            I => \N__22582\
        );

    \I__5466\ : LocalMux
    port map (
            O => \N__22599\,
            I => \N__22582\
        );

    \I__5465\ : ClkMux
    port map (
            O => \N__22598\,
            I => \N__22579\
        );

    \I__5464\ : ClkMux
    port map (
            O => \N__22597\,
            I => \N__22574\
        );

    \I__5463\ : ClkMux
    port map (
            O => \N__22596\,
            I => \N__22566\
        );

    \I__5462\ : ClkMux
    port map (
            O => \N__22595\,
            I => \N__22558\
        );

    \I__5461\ : ClkMux
    port map (
            O => \N__22594\,
            I => \N__22555\
        );

    \I__5460\ : ClkMux
    port map (
            O => \N__22593\,
            I => \N__22551\
        );

    \I__5459\ : LocalMux
    port map (
            O => \N__22590\,
            I => \N__22547\
        );

    \I__5458\ : ClkMux
    port map (
            O => \N__22589\,
            I => \N__22544\
        );

    \I__5457\ : ClkMux
    port map (
            O => \N__22588\,
            I => \N__22541\
        );

    \I__5456\ : ClkMux
    port map (
            O => \N__22587\,
            I => \N__22538\
        );

    \I__5455\ : Span4Mux_v
    port map (
            O => \N__22582\,
            I => \N__22533\
        );

    \I__5454\ : LocalMux
    port map (
            O => \N__22579\,
            I => \N__22533\
        );

    \I__5453\ : ClkMux
    port map (
            O => \N__22578\,
            I => \N__22530\
        );

    \I__5452\ : ClkMux
    port map (
            O => \N__22577\,
            I => \N__22527\
        );

    \I__5451\ : LocalMux
    port map (
            O => \N__22574\,
            I => \N__22524\
        );

    \I__5450\ : ClkMux
    port map (
            O => \N__22573\,
            I => \N__22521\
        );

    \I__5449\ : ClkMux
    port map (
            O => \N__22572\,
            I => \N__22518\
        );

    \I__5448\ : ClkMux
    port map (
            O => \N__22571\,
            I => \N__22511\
        );

    \I__5447\ : ClkMux
    port map (
            O => \N__22570\,
            I => \N__22506\
        );

    \I__5446\ : ClkMux
    port map (
            O => \N__22569\,
            I => \N__22503\
        );

    \I__5445\ : LocalMux
    port map (
            O => \N__22566\,
            I => \N__22497\
        );

    \I__5444\ : ClkMux
    port map (
            O => \N__22565\,
            I => \N__22493\
        );

    \I__5443\ : ClkMux
    port map (
            O => \N__22564\,
            I => \N__22490\
        );

    \I__5442\ : ClkMux
    port map (
            O => \N__22563\,
            I => \N__22487\
        );

    \I__5441\ : ClkMux
    port map (
            O => \N__22562\,
            I => \N__22484\
        );

    \I__5440\ : ClkMux
    port map (
            O => \N__22561\,
            I => \N__22477\
        );

    \I__5439\ : LocalMux
    port map (
            O => \N__22558\,
            I => \N__22472\
        );

    \I__5438\ : LocalMux
    port map (
            O => \N__22555\,
            I => \N__22472\
        );

    \I__5437\ : ClkMux
    port map (
            O => \N__22554\,
            I => \N__22469\
        );

    \I__5436\ : LocalMux
    port map (
            O => \N__22551\,
            I => \N__22465\
        );

    \I__5435\ : ClkMux
    port map (
            O => \N__22550\,
            I => \N__22462\
        );

    \I__5434\ : Span4Mux_v
    port map (
            O => \N__22547\,
            I => \N__22456\
        );

    \I__5433\ : LocalMux
    port map (
            O => \N__22544\,
            I => \N__22456\
        );

    \I__5432\ : LocalMux
    port map (
            O => \N__22541\,
            I => \N__22448\
        );

    \I__5431\ : LocalMux
    port map (
            O => \N__22538\,
            I => \N__22448\
        );

    \I__5430\ : Span4Mux_v
    port map (
            O => \N__22533\,
            I => \N__22444\
        );

    \I__5429\ : LocalMux
    port map (
            O => \N__22530\,
            I => \N__22439\
        );

    \I__5428\ : LocalMux
    port map (
            O => \N__22527\,
            I => \N__22439\
        );

    \I__5427\ : Span4Mux_h
    port map (
            O => \N__22524\,
            I => \N__22432\
        );

    \I__5426\ : LocalMux
    port map (
            O => \N__22521\,
            I => \N__22432\
        );

    \I__5425\ : LocalMux
    port map (
            O => \N__22518\,
            I => \N__22432\
        );

    \I__5424\ : ClkMux
    port map (
            O => \N__22517\,
            I => \N__22429\
        );

    \I__5423\ : ClkMux
    port map (
            O => \N__22516\,
            I => \N__22426\
        );

    \I__5422\ : ClkMux
    port map (
            O => \N__22515\,
            I => \N__22423\
        );

    \I__5421\ : ClkMux
    port map (
            O => \N__22514\,
            I => \N__22420\
        );

    \I__5420\ : LocalMux
    port map (
            O => \N__22511\,
            I => \N__22416\
        );

    \I__5419\ : ClkMux
    port map (
            O => \N__22510\,
            I => \N__22413\
        );

    \I__5418\ : ClkMux
    port map (
            O => \N__22509\,
            I => \N__22407\
        );

    \I__5417\ : LocalMux
    port map (
            O => \N__22506\,
            I => \N__22402\
        );

    \I__5416\ : LocalMux
    port map (
            O => \N__22503\,
            I => \N__22399\
        );

    \I__5415\ : ClkMux
    port map (
            O => \N__22502\,
            I => \N__22396\
        );

    \I__5414\ : ClkMux
    port map (
            O => \N__22501\,
            I => \N__22393\
        );

    \I__5413\ : ClkMux
    port map (
            O => \N__22500\,
            I => \N__22389\
        );

    \I__5412\ : Span4Mux_v
    port map (
            O => \N__22497\,
            I => \N__22385\
        );

    \I__5411\ : ClkMux
    port map (
            O => \N__22496\,
            I => \N__22382\
        );

    \I__5410\ : LocalMux
    port map (
            O => \N__22493\,
            I => \N__22377\
        );

    \I__5409\ : LocalMux
    port map (
            O => \N__22490\,
            I => \N__22374\
        );

    \I__5408\ : LocalMux
    port map (
            O => \N__22487\,
            I => \N__22371\
        );

    \I__5407\ : LocalMux
    port map (
            O => \N__22484\,
            I => \N__22368\
        );

    \I__5406\ : ClkMux
    port map (
            O => \N__22483\,
            I => \N__22365\
        );

    \I__5405\ : ClkMux
    port map (
            O => \N__22482\,
            I => \N__22362\
        );

    \I__5404\ : ClkMux
    port map (
            O => \N__22481\,
            I => \N__22359\
        );

    \I__5403\ : ClkMux
    port map (
            O => \N__22480\,
            I => \N__22356\
        );

    \I__5402\ : LocalMux
    port map (
            O => \N__22477\,
            I => \N__22348\
        );

    \I__5401\ : Span4Mux_v
    port map (
            O => \N__22472\,
            I => \N__22343\
        );

    \I__5400\ : LocalMux
    port map (
            O => \N__22469\,
            I => \N__22343\
        );

    \I__5399\ : ClkMux
    port map (
            O => \N__22468\,
            I => \N__22340\
        );

    \I__5398\ : Span4Mux_h
    port map (
            O => \N__22465\,
            I => \N__22335\
        );

    \I__5397\ : LocalMux
    port map (
            O => \N__22462\,
            I => \N__22335\
        );

    \I__5396\ : ClkMux
    port map (
            O => \N__22461\,
            I => \N__22332\
        );

    \I__5395\ : Span4Mux_h
    port map (
            O => \N__22456\,
            I => \N__22329\
        );

    \I__5394\ : ClkMux
    port map (
            O => \N__22455\,
            I => \N__22326\
        );

    \I__5393\ : ClkMux
    port map (
            O => \N__22454\,
            I => \N__22323\
        );

    \I__5392\ : ClkMux
    port map (
            O => \N__22453\,
            I => \N__22320\
        );

    \I__5391\ : Span4Mux_v
    port map (
            O => \N__22448\,
            I => \N__22315\
        );

    \I__5390\ : ClkMux
    port map (
            O => \N__22447\,
            I => \N__22312\
        );

    \I__5389\ : Span4Mux_h
    port map (
            O => \N__22444\,
            I => \N__22297\
        );

    \I__5388\ : Span4Mux_h
    port map (
            O => \N__22439\,
            I => \N__22297\
        );

    \I__5387\ : Span4Mux_v
    port map (
            O => \N__22432\,
            I => \N__22297\
        );

    \I__5386\ : LocalMux
    port map (
            O => \N__22429\,
            I => \N__22297\
        );

    \I__5385\ : LocalMux
    port map (
            O => \N__22426\,
            I => \N__22297\
        );

    \I__5384\ : LocalMux
    port map (
            O => \N__22423\,
            I => \N__22297\
        );

    \I__5383\ : LocalMux
    port map (
            O => \N__22420\,
            I => \N__22297\
        );

    \I__5382\ : ClkMux
    port map (
            O => \N__22419\,
            I => \N__22294\
        );

    \I__5381\ : Span4Mux_v
    port map (
            O => \N__22416\,
            I => \N__22291\
        );

    \I__5380\ : LocalMux
    port map (
            O => \N__22413\,
            I => \N__22288\
        );

    \I__5379\ : ClkMux
    port map (
            O => \N__22412\,
            I => \N__22285\
        );

    \I__5378\ : ClkMux
    port map (
            O => \N__22411\,
            I => \N__22282\
        );

    \I__5377\ : ClkMux
    port map (
            O => \N__22410\,
            I => \N__22277\
        );

    \I__5376\ : LocalMux
    port map (
            O => \N__22407\,
            I => \N__22274\
        );

    \I__5375\ : ClkMux
    port map (
            O => \N__22406\,
            I => \N__22271\
        );

    \I__5374\ : ClkMux
    port map (
            O => \N__22405\,
            I => \N__22268\
        );

    \I__5373\ : Span4Mux_v
    port map (
            O => \N__22402\,
            I => \N__22264\
        );

    \I__5372\ : Span4Mux_v
    port map (
            O => \N__22399\,
            I => \N__22256\
        );

    \I__5371\ : LocalMux
    port map (
            O => \N__22396\,
            I => \N__22256\
        );

    \I__5370\ : LocalMux
    port map (
            O => \N__22393\,
            I => \N__22256\
        );

    \I__5369\ : ClkMux
    port map (
            O => \N__22392\,
            I => \N__22253\
        );

    \I__5368\ : LocalMux
    port map (
            O => \N__22389\,
            I => \N__22248\
        );

    \I__5367\ : ClkMux
    port map (
            O => \N__22388\,
            I => \N__22245\
        );

    \I__5366\ : Span4Mux_v
    port map (
            O => \N__22385\,
            I => \N__22237\
        );

    \I__5365\ : LocalMux
    port map (
            O => \N__22382\,
            I => \N__22237\
        );

    \I__5364\ : ClkMux
    port map (
            O => \N__22381\,
            I => \N__22234\
        );

    \I__5363\ : ClkMux
    port map (
            O => \N__22380\,
            I => \N__22231\
        );

    \I__5362\ : Span4Mux_v
    port map (
            O => \N__22377\,
            I => \N__22219\
        );

    \I__5361\ : Span4Mux_h
    port map (
            O => \N__22374\,
            I => \N__22219\
        );

    \I__5360\ : Span4Mux_h
    port map (
            O => \N__22371\,
            I => \N__22219\
        );

    \I__5359\ : Span4Mux_h
    port map (
            O => \N__22368\,
            I => \N__22219\
        );

    \I__5358\ : LocalMux
    port map (
            O => \N__22365\,
            I => \N__22219\
        );

    \I__5357\ : LocalMux
    port map (
            O => \N__22362\,
            I => \N__22216\
        );

    \I__5356\ : LocalMux
    port map (
            O => \N__22359\,
            I => \N__22213\
        );

    \I__5355\ : LocalMux
    port map (
            O => \N__22356\,
            I => \N__22210\
        );

    \I__5354\ : ClkMux
    port map (
            O => \N__22355\,
            I => \N__22207\
        );

    \I__5353\ : ClkMux
    port map (
            O => \N__22354\,
            I => \N__22204\
        );

    \I__5352\ : ClkMux
    port map (
            O => \N__22353\,
            I => \N__22201\
        );

    \I__5351\ : ClkMux
    port map (
            O => \N__22352\,
            I => \N__22198\
        );

    \I__5350\ : ClkMux
    port map (
            O => \N__22351\,
            I => \N__22195\
        );

    \I__5349\ : Span4Mux_v
    port map (
            O => \N__22348\,
            I => \N__22188\
        );

    \I__5348\ : Span4Mux_v
    port map (
            O => \N__22343\,
            I => \N__22188\
        );

    \I__5347\ : LocalMux
    port map (
            O => \N__22340\,
            I => \N__22188\
        );

    \I__5346\ : Span4Mux_v
    port map (
            O => \N__22335\,
            I => \N__22182\
        );

    \I__5345\ : LocalMux
    port map (
            O => \N__22332\,
            I => \N__22182\
        );

    \I__5344\ : Span4Mux_h
    port map (
            O => \N__22329\,
            I => \N__22177\
        );

    \I__5343\ : LocalMux
    port map (
            O => \N__22326\,
            I => \N__22177\
        );

    \I__5342\ : LocalMux
    port map (
            O => \N__22323\,
            I => \N__22174\
        );

    \I__5341\ : LocalMux
    port map (
            O => \N__22320\,
            I => \N__22171\
        );

    \I__5340\ : ClkMux
    port map (
            O => \N__22319\,
            I => \N__22168\
        );

    \I__5339\ : ClkMux
    port map (
            O => \N__22318\,
            I => \N__22165\
        );

    \I__5338\ : Span4Mux_h
    port map (
            O => \N__22315\,
            I => \N__22162\
        );

    \I__5337\ : LocalMux
    port map (
            O => \N__22312\,
            I => \N__22155\
        );

    \I__5336\ : Span4Mux_v
    port map (
            O => \N__22297\,
            I => \N__22155\
        );

    \I__5335\ : LocalMux
    port map (
            O => \N__22294\,
            I => \N__22155\
        );

    \I__5334\ : Span4Mux_h
    port map (
            O => \N__22291\,
            I => \N__22150\
        );

    \I__5333\ : Span4Mux_h
    port map (
            O => \N__22288\,
            I => \N__22150\
        );

    \I__5332\ : LocalMux
    port map (
            O => \N__22285\,
            I => \N__22145\
        );

    \I__5331\ : LocalMux
    port map (
            O => \N__22282\,
            I => \N__22145\
        );

    \I__5330\ : ClkMux
    port map (
            O => \N__22281\,
            I => \N__22142\
        );

    \I__5329\ : ClkMux
    port map (
            O => \N__22280\,
            I => \N__22139\
        );

    \I__5328\ : LocalMux
    port map (
            O => \N__22277\,
            I => \N__22136\
        );

    \I__5327\ : Span4Mux_h
    port map (
            O => \N__22274\,
            I => \N__22129\
        );

    \I__5326\ : LocalMux
    port map (
            O => \N__22271\,
            I => \N__22129\
        );

    \I__5325\ : LocalMux
    port map (
            O => \N__22268\,
            I => \N__22129\
        );

    \I__5324\ : ClkMux
    port map (
            O => \N__22267\,
            I => \N__22126\
        );

    \I__5323\ : Span4Mux_h
    port map (
            O => \N__22264\,
            I => \N__22123\
        );

    \I__5322\ : ClkMux
    port map (
            O => \N__22263\,
            I => \N__22120\
        );

    \I__5321\ : Span4Mux_v
    port map (
            O => \N__22256\,
            I => \N__22115\
        );

    \I__5320\ : LocalMux
    port map (
            O => \N__22253\,
            I => \N__22115\
        );

    \I__5319\ : ClkMux
    port map (
            O => \N__22252\,
            I => \N__22111\
        );

    \I__5318\ : ClkMux
    port map (
            O => \N__22251\,
            I => \N__22108\
        );

    \I__5317\ : Span4Mux_v
    port map (
            O => \N__22248\,
            I => \N__22103\
        );

    \I__5316\ : LocalMux
    port map (
            O => \N__22245\,
            I => \N__22103\
        );

    \I__5315\ : ClkMux
    port map (
            O => \N__22244\,
            I => \N__22099\
        );

    \I__5314\ : ClkMux
    port map (
            O => \N__22243\,
            I => \N__22096\
        );

    \I__5313\ : ClkMux
    port map (
            O => \N__22242\,
            I => \N__22093\
        );

    \I__5312\ : Span4Mux_v
    port map (
            O => \N__22237\,
            I => \N__22090\
        );

    \I__5311\ : LocalMux
    port map (
            O => \N__22234\,
            I => \N__22085\
        );

    \I__5310\ : LocalMux
    port map (
            O => \N__22231\,
            I => \N__22085\
        );

    \I__5309\ : ClkMux
    port map (
            O => \N__22230\,
            I => \N__22078\
        );

    \I__5308\ : Span4Mux_v
    port map (
            O => \N__22219\,
            I => \N__22075\
        );

    \I__5307\ : Span4Mux_h
    port map (
            O => \N__22216\,
            I => \N__22072\
        );

    \I__5306\ : Span4Mux_v
    port map (
            O => \N__22213\,
            I => \N__22069\
        );

    \I__5305\ : Span4Mux_v
    port map (
            O => \N__22210\,
            I => \N__22064\
        );

    \I__5304\ : LocalMux
    port map (
            O => \N__22207\,
            I => \N__22064\
        );

    \I__5303\ : LocalMux
    port map (
            O => \N__22204\,
            I => \N__22053\
        );

    \I__5302\ : LocalMux
    port map (
            O => \N__22201\,
            I => \N__22053\
        );

    \I__5301\ : LocalMux
    port map (
            O => \N__22198\,
            I => \N__22053\
        );

    \I__5300\ : LocalMux
    port map (
            O => \N__22195\,
            I => \N__22053\
        );

    \I__5299\ : Span4Mux_h
    port map (
            O => \N__22188\,
            I => \N__22053\
        );

    \I__5298\ : ClkMux
    port map (
            O => \N__22187\,
            I => \N__22050\
        );

    \I__5297\ : Span4Mux_h
    port map (
            O => \N__22182\,
            I => \N__22047\
        );

    \I__5296\ : Span4Mux_v
    port map (
            O => \N__22177\,
            I => \N__22044\
        );

    \I__5295\ : Span4Mux_h
    port map (
            O => \N__22174\,
            I => \N__22035\
        );

    \I__5294\ : Span4Mux_v
    port map (
            O => \N__22171\,
            I => \N__22035\
        );

    \I__5293\ : LocalMux
    port map (
            O => \N__22168\,
            I => \N__22035\
        );

    \I__5292\ : LocalMux
    port map (
            O => \N__22165\,
            I => \N__22035\
        );

    \I__5291\ : Span4Mux_h
    port map (
            O => \N__22162\,
            I => \N__22030\
        );

    \I__5290\ : Span4Mux_v
    port map (
            O => \N__22155\,
            I => \N__22030\
        );

    \I__5289\ : Span4Mux_v
    port map (
            O => \N__22150\,
            I => \N__22021\
        );

    \I__5288\ : Span4Mux_v
    port map (
            O => \N__22145\,
            I => \N__22021\
        );

    \I__5287\ : LocalMux
    port map (
            O => \N__22142\,
            I => \N__22021\
        );

    \I__5286\ : LocalMux
    port map (
            O => \N__22139\,
            I => \N__22021\
        );

    \I__5285\ : Span4Mux_h
    port map (
            O => \N__22136\,
            I => \N__22014\
        );

    \I__5284\ : Span4Mux_v
    port map (
            O => \N__22129\,
            I => \N__22014\
        );

    \I__5283\ : LocalMux
    port map (
            O => \N__22126\,
            I => \N__22014\
        );

    \I__5282\ : Span4Mux_v
    port map (
            O => \N__22123\,
            I => \N__22009\
        );

    \I__5281\ : LocalMux
    port map (
            O => \N__22120\,
            I => \N__22009\
        );

    \I__5280\ : Span4Mux_v
    port map (
            O => \N__22115\,
            I => \N__22006\
        );

    \I__5279\ : ClkMux
    port map (
            O => \N__22114\,
            I => \N__22003\
        );

    \I__5278\ : LocalMux
    port map (
            O => \N__22111\,
            I => \N__21998\
        );

    \I__5277\ : LocalMux
    port map (
            O => \N__22108\,
            I => \N__21998\
        );

    \I__5276\ : Span4Mux_v
    port map (
            O => \N__22103\,
            I => \N__21995\
        );

    \I__5275\ : ClkMux
    port map (
            O => \N__22102\,
            I => \N__21992\
        );

    \I__5274\ : LocalMux
    port map (
            O => \N__22099\,
            I => \N__21989\
        );

    \I__5273\ : LocalMux
    port map (
            O => \N__22096\,
            I => \N__21986\
        );

    \I__5272\ : LocalMux
    port map (
            O => \N__22093\,
            I => \N__21983\
        );

    \I__5271\ : Span4Mux_h
    port map (
            O => \N__22090\,
            I => \N__21978\
        );

    \I__5270\ : Span4Mux_v
    port map (
            O => \N__22085\,
            I => \N__21978\
        );

    \I__5269\ : ClkMux
    port map (
            O => \N__22084\,
            I => \N__21975\
        );

    \I__5268\ : ClkMux
    port map (
            O => \N__22083\,
            I => \N__21972\
        );

    \I__5267\ : ClkMux
    port map (
            O => \N__22082\,
            I => \N__21968\
        );

    \I__5266\ : ClkMux
    port map (
            O => \N__22081\,
            I => \N__21965\
        );

    \I__5265\ : LocalMux
    port map (
            O => \N__22078\,
            I => \N__21961\
        );

    \I__5264\ : Span4Mux_h
    port map (
            O => \N__22075\,
            I => \N__21948\
        );

    \I__5263\ : Span4Mux_h
    port map (
            O => \N__22072\,
            I => \N__21948\
        );

    \I__5262\ : Span4Mux_h
    port map (
            O => \N__22069\,
            I => \N__21948\
        );

    \I__5261\ : Span4Mux_v
    port map (
            O => \N__22064\,
            I => \N__21948\
        );

    \I__5260\ : Span4Mux_v
    port map (
            O => \N__22053\,
            I => \N__21948\
        );

    \I__5259\ : LocalMux
    port map (
            O => \N__22050\,
            I => \N__21948\
        );

    \I__5258\ : Span4Mux_v
    port map (
            O => \N__22047\,
            I => \N__21940\
        );

    \I__5257\ : Span4Mux_h
    port map (
            O => \N__22044\,
            I => \N__21940\
        );

    \I__5256\ : Span4Mux_v
    port map (
            O => \N__22035\,
            I => \N__21937\
        );

    \I__5255\ : Span4Mux_h
    port map (
            O => \N__22030\,
            I => \N__21932\
        );

    \I__5254\ : Span4Mux_v
    port map (
            O => \N__22021\,
            I => \N__21932\
        );

    \I__5253\ : Span4Mux_h
    port map (
            O => \N__22014\,
            I => \N__21923\
        );

    \I__5252\ : Span4Mux_h
    port map (
            O => \N__22009\,
            I => \N__21923\
        );

    \I__5251\ : Span4Mux_v
    port map (
            O => \N__22006\,
            I => \N__21923\
        );

    \I__5250\ : LocalMux
    port map (
            O => \N__22003\,
            I => \N__21923\
        );

    \I__5249\ : Span4Mux_v
    port map (
            O => \N__21998\,
            I => \N__21916\
        );

    \I__5248\ : Span4Mux_v
    port map (
            O => \N__21995\,
            I => \N__21916\
        );

    \I__5247\ : LocalMux
    port map (
            O => \N__21992\,
            I => \N__21916\
        );

    \I__5246\ : Span4Mux_v
    port map (
            O => \N__21989\,
            I => \N__21905\
        );

    \I__5245\ : Span4Mux_v
    port map (
            O => \N__21986\,
            I => \N__21905\
        );

    \I__5244\ : Span4Mux_v
    port map (
            O => \N__21983\,
            I => \N__21905\
        );

    \I__5243\ : Span4Mux_h
    port map (
            O => \N__21978\,
            I => \N__21905\
        );

    \I__5242\ : LocalMux
    port map (
            O => \N__21975\,
            I => \N__21905\
        );

    \I__5241\ : LocalMux
    port map (
            O => \N__21972\,
            I => \N__21902\
        );

    \I__5240\ : ClkMux
    port map (
            O => \N__21971\,
            I => \N__21899\
        );

    \I__5239\ : LocalMux
    port map (
            O => \N__21968\,
            I => \N__21894\
        );

    \I__5238\ : LocalMux
    port map (
            O => \N__21965\,
            I => \N__21894\
        );

    \I__5237\ : ClkMux
    port map (
            O => \N__21964\,
            I => \N__21891\
        );

    \I__5236\ : Span4Mux_h
    port map (
            O => \N__21961\,
            I => \N__21885\
        );

    \I__5235\ : Span4Mux_v
    port map (
            O => \N__21948\,
            I => \N__21885\
        );

    \I__5234\ : ClkMux
    port map (
            O => \N__21947\,
            I => \N__21881\
        );

    \I__5233\ : ClkMux
    port map (
            O => \N__21946\,
            I => \N__21878\
        );

    \I__5232\ : ClkMux
    port map (
            O => \N__21945\,
            I => \N__21875\
        );

    \I__5231\ : Span4Mux_h
    port map (
            O => \N__21940\,
            I => \N__21871\
        );

    \I__5230\ : Span4Mux_h
    port map (
            O => \N__21937\,
            I => \N__21866\
        );

    \I__5229\ : Span4Mux_h
    port map (
            O => \N__21932\,
            I => \N__21866\
        );

    \I__5228\ : Span4Mux_h
    port map (
            O => \N__21923\,
            I => \N__21861\
        );

    \I__5227\ : Span4Mux_v
    port map (
            O => \N__21916\,
            I => \N__21861\
        );

    \I__5226\ : Span4Mux_v
    port map (
            O => \N__21905\,
            I => \N__21850\
        );

    \I__5225\ : Span4Mux_v
    port map (
            O => \N__21902\,
            I => \N__21850\
        );

    \I__5224\ : LocalMux
    port map (
            O => \N__21899\,
            I => \N__21850\
        );

    \I__5223\ : Span4Mux_v
    port map (
            O => \N__21894\,
            I => \N__21850\
        );

    \I__5222\ : LocalMux
    port map (
            O => \N__21891\,
            I => \N__21850\
        );

    \I__5221\ : ClkMux
    port map (
            O => \N__21890\,
            I => \N__21847\
        );

    \I__5220\ : Span4Mux_h
    port map (
            O => \N__21885\,
            I => \N__21844\
        );

    \I__5219\ : ClkMux
    port map (
            O => \N__21884\,
            I => \N__21841\
        );

    \I__5218\ : LocalMux
    port map (
            O => \N__21881\,
            I => \N__21838\
        );

    \I__5217\ : LocalMux
    port map (
            O => \N__21878\,
            I => \N__21833\
        );

    \I__5216\ : LocalMux
    port map (
            O => \N__21875\,
            I => \N__21833\
        );

    \I__5215\ : ClkMux
    port map (
            O => \N__21874\,
            I => \N__21830\
        );

    \I__5214\ : Span4Mux_h
    port map (
            O => \N__21871\,
            I => \N__21827\
        );

    \I__5213\ : Span4Mux_h
    port map (
            O => \N__21866\,
            I => \N__21824\
        );

    \I__5212\ : Span4Mux_h
    port map (
            O => \N__21861\,
            I => \N__21821\
        );

    \I__5211\ : Sp12to4
    port map (
            O => \N__21850\,
            I => \N__21818\
        );

    \I__5210\ : LocalMux
    port map (
            O => \N__21847\,
            I => \N__21811\
        );

    \I__5209\ : Sp12to4
    port map (
            O => \N__21844\,
            I => \N__21811\
        );

    \I__5208\ : LocalMux
    port map (
            O => \N__21841\,
            I => \N__21811\
        );

    \I__5207\ : Span4Mux_h
    port map (
            O => \N__21838\,
            I => \N__21804\
        );

    \I__5206\ : Span4Mux_v
    port map (
            O => \N__21833\,
            I => \N__21804\
        );

    \I__5205\ : LocalMux
    port map (
            O => \N__21830\,
            I => \N__21804\
        );

    \I__5204\ : Span4Mux_h
    port map (
            O => \N__21827\,
            I => \N__21801\
        );

    \I__5203\ : Span4Mux_h
    port map (
            O => \N__21824\,
            I => \N__21798\
        );

    \I__5202\ : Sp12to4
    port map (
            O => \N__21821\,
            I => \N__21793\
        );

    \I__5201\ : Span12Mux_h
    port map (
            O => \N__21818\,
            I => \N__21793\
        );

    \I__5200\ : Span12Mux_v
    port map (
            O => \N__21811\,
            I => \N__21788\
        );

    \I__5199\ : Sp12to4
    port map (
            O => \N__21804\,
            I => \N__21788\
        );

    \I__5198\ : IoSpan4Mux
    port map (
            O => \N__21801\,
            I => \N__21785\
        );

    \I__5197\ : Span4Mux_h
    port map (
            O => \N__21798\,
            I => \N__21782\
        );

    \I__5196\ : Span12Mux_h
    port map (
            O => \N__21793\,
            I => \N__21779\
        );

    \I__5195\ : Span12Mux_h
    port map (
            O => \N__21788\,
            I => \N__21776\
        );

    \I__5194\ : Odrv4
    port map (
            O => \N__21785\,
            I => clk
        );

    \I__5193\ : Odrv4
    port map (
            O => \N__21782\,
            I => clk
        );

    \I__5192\ : Odrv12
    port map (
            O => \N__21779\,
            I => clk
        );

    \I__5191\ : Odrv12
    port map (
            O => \N__21776\,
            I => clk
        );

    \I__5190\ : InMux
    port map (
            O => \N__21767\,
            I => \N__21763\
        );

    \I__5189\ : InMux
    port map (
            O => \N__21766\,
            I => \N__21760\
        );

    \I__5188\ : LocalMux
    port map (
            O => \N__21763\,
            I => \N__21757\
        );

    \I__5187\ : LocalMux
    port map (
            O => \N__21760\,
            I => \b2v_inst1.N_29_mux\
        );

    \I__5186\ : Odrv4
    port map (
            O => \N__21757\,
            I => \b2v_inst1.N_29_mux\
        );

    \I__5185\ : CascadeMux
    port map (
            O => \N__21752\,
            I => \b2v_inst1.r_SM_Main_1_sqmuxa_1_cascade_\
        );

    \I__5184\ : InMux
    port map (
            O => \N__21749\,
            I => \N__21742\
        );

    \I__5183\ : InMux
    port map (
            O => \N__21748\,
            I => \N__21742\
        );

    \I__5182\ : InMux
    port map (
            O => \N__21747\,
            I => \N__21739\
        );

    \I__5181\ : LocalMux
    port map (
            O => \N__21742\,
            I => \b2v_inst1.un1_r_SM_Main_1_sqmuxa_0\
        );

    \I__5180\ : LocalMux
    port map (
            O => \N__21739\,
            I => \b2v_inst1.un1_r_SM_Main_1_sqmuxa_0\
        );

    \I__5179\ : InMux
    port map (
            O => \N__21734\,
            I => \N__21729\
        );

    \I__5178\ : InMux
    port map (
            O => \N__21733\,
            I => \N__21726\
        );

    \I__5177\ : InMux
    port map (
            O => \N__21732\,
            I => \N__21720\
        );

    \I__5176\ : LocalMux
    port map (
            O => \N__21729\,
            I => \N__21715\
        );

    \I__5175\ : LocalMux
    port map (
            O => \N__21726\,
            I => \N__21715\
        );

    \I__5174\ : InMux
    port map (
            O => \N__21725\,
            I => \N__21712\
        );

    \I__5173\ : InMux
    port map (
            O => \N__21724\,
            I => \N__21709\
        );

    \I__5172\ : InMux
    port map (
            O => \N__21723\,
            I => \N__21706\
        );

    \I__5171\ : LocalMux
    port map (
            O => \N__21720\,
            I => \b2v_inst1.un1_r_Clk_Count_ac0_1_out\
        );

    \I__5170\ : Odrv4
    port map (
            O => \N__21715\,
            I => \b2v_inst1.un1_r_Clk_Count_ac0_1_out\
        );

    \I__5169\ : LocalMux
    port map (
            O => \N__21712\,
            I => \b2v_inst1.un1_r_Clk_Count_ac0_1_out\
        );

    \I__5168\ : LocalMux
    port map (
            O => \N__21709\,
            I => \b2v_inst1.un1_r_Clk_Count_ac0_1_out\
        );

    \I__5167\ : LocalMux
    port map (
            O => \N__21706\,
            I => \b2v_inst1.un1_r_Clk_Count_ac0_1_out\
        );

    \I__5166\ : CascadeMux
    port map (
            O => \N__21695\,
            I => \N__21686\
        );

    \I__5165\ : InMux
    port map (
            O => \N__21694\,
            I => \N__21681\
        );

    \I__5164\ : InMux
    port map (
            O => \N__21693\,
            I => \N__21681\
        );

    \I__5163\ : CascadeMux
    port map (
            O => \N__21692\,
            I => \N__21678\
        );

    \I__5162\ : CascadeMux
    port map (
            O => \N__21691\,
            I => \N__21675\
        );

    \I__5161\ : InMux
    port map (
            O => \N__21690\,
            I => \N__21670\
        );

    \I__5160\ : InMux
    port map (
            O => \N__21689\,
            I => \N__21670\
        );

    \I__5159\ : InMux
    port map (
            O => \N__21686\,
            I => \N__21667\
        );

    \I__5158\ : LocalMux
    port map (
            O => \N__21681\,
            I => \N__21663\
        );

    \I__5157\ : InMux
    port map (
            O => \N__21678\,
            I => \N__21653\
        );

    \I__5156\ : InMux
    port map (
            O => \N__21675\,
            I => \N__21650\
        );

    \I__5155\ : LocalMux
    port map (
            O => \N__21670\,
            I => \N__21647\
        );

    \I__5154\ : LocalMux
    port map (
            O => \N__21667\,
            I => \N__21644\
        );

    \I__5153\ : CascadeMux
    port map (
            O => \N__21666\,
            I => \N__21640\
        );

    \I__5152\ : Span4Mux_h
    port map (
            O => \N__21663\,
            I => \N__21636\
        );

    \I__5151\ : InMux
    port map (
            O => \N__21662\,
            I => \N__21633\
        );

    \I__5150\ : InMux
    port map (
            O => \N__21661\,
            I => \N__21626\
        );

    \I__5149\ : InMux
    port map (
            O => \N__21660\,
            I => \N__21626\
        );

    \I__5148\ : InMux
    port map (
            O => \N__21659\,
            I => \N__21626\
        );

    \I__5147\ : InMux
    port map (
            O => \N__21658\,
            I => \N__21623\
        );

    \I__5146\ : InMux
    port map (
            O => \N__21657\,
            I => \N__21620\
        );

    \I__5145\ : InMux
    port map (
            O => \N__21656\,
            I => \N__21617\
        );

    \I__5144\ : LocalMux
    port map (
            O => \N__21653\,
            I => \N__21612\
        );

    \I__5143\ : LocalMux
    port map (
            O => \N__21650\,
            I => \N__21612\
        );

    \I__5142\ : Span4Mux_h
    port map (
            O => \N__21647\,
            I => \N__21607\
        );

    \I__5141\ : Span4Mux_h
    port map (
            O => \N__21644\,
            I => \N__21607\
        );

    \I__5140\ : InMux
    port map (
            O => \N__21643\,
            I => \N__21600\
        );

    \I__5139\ : InMux
    port map (
            O => \N__21640\,
            I => \N__21600\
        );

    \I__5138\ : InMux
    port map (
            O => \N__21639\,
            I => \N__21600\
        );

    \I__5137\ : Odrv4
    port map (
            O => \N__21636\,
            I => \b2v_inst1.r_Clk_CountZ0Z_3\
        );

    \I__5136\ : LocalMux
    port map (
            O => \N__21633\,
            I => \b2v_inst1.r_Clk_CountZ0Z_3\
        );

    \I__5135\ : LocalMux
    port map (
            O => \N__21626\,
            I => \b2v_inst1.r_Clk_CountZ0Z_3\
        );

    \I__5134\ : LocalMux
    port map (
            O => \N__21623\,
            I => \b2v_inst1.r_Clk_CountZ0Z_3\
        );

    \I__5133\ : LocalMux
    port map (
            O => \N__21620\,
            I => \b2v_inst1.r_Clk_CountZ0Z_3\
        );

    \I__5132\ : LocalMux
    port map (
            O => \N__21617\,
            I => \b2v_inst1.r_Clk_CountZ0Z_3\
        );

    \I__5131\ : Odrv4
    port map (
            O => \N__21612\,
            I => \b2v_inst1.r_Clk_CountZ0Z_3\
        );

    \I__5130\ : Odrv4
    port map (
            O => \N__21607\,
            I => \b2v_inst1.r_Clk_CountZ0Z_3\
        );

    \I__5129\ : LocalMux
    port map (
            O => \N__21600\,
            I => \b2v_inst1.r_Clk_CountZ0Z_3\
        );

    \I__5128\ : CascadeMux
    port map (
            O => \N__21581\,
            I => \b2v_inst1.g0_3_1_cascade_\
        );

    \I__5127\ : InMux
    port map (
            O => \N__21578\,
            I => \N__21575\
        );

    \I__5126\ : LocalMux
    port map (
            O => \N__21575\,
            I => \b2v_inst1.N_14_0_0\
        );

    \I__5125\ : CascadeMux
    port map (
            O => \N__21572\,
            I => \b2v_inst1.N_14_0_0_cascade_\
        );

    \I__5124\ : InMux
    port map (
            O => \N__21569\,
            I => \N__21566\
        );

    \I__5123\ : LocalMux
    port map (
            O => \N__21566\,
            I => \b2v_inst1.N_29_mux_0\
        );

    \I__5122\ : InMux
    port map (
            O => \N__21563\,
            I => \N__21556\
        );

    \I__5121\ : CascadeMux
    port map (
            O => \N__21562\,
            I => \N__21553\
        );

    \I__5120\ : InMux
    port map (
            O => \N__21561\,
            I => \N__21549\
        );

    \I__5119\ : InMux
    port map (
            O => \N__21560\,
            I => \N__21544\
        );

    \I__5118\ : InMux
    port map (
            O => \N__21559\,
            I => \N__21544\
        );

    \I__5117\ : LocalMux
    port map (
            O => \N__21556\,
            I => \N__21539\
        );

    \I__5116\ : InMux
    port map (
            O => \N__21553\,
            I => \N__21534\
        );

    \I__5115\ : InMux
    port map (
            O => \N__21552\,
            I => \N__21534\
        );

    \I__5114\ : LocalMux
    port map (
            O => \N__21549\,
            I => \N__21522\
        );

    \I__5113\ : LocalMux
    port map (
            O => \N__21544\,
            I => \N__21522\
        );

    \I__5112\ : InMux
    port map (
            O => \N__21543\,
            I => \N__21517\
        );

    \I__5111\ : InMux
    port map (
            O => \N__21542\,
            I => \N__21517\
        );

    \I__5110\ : Span4Mux_v
    port map (
            O => \N__21539\,
            I => \N__21512\
        );

    \I__5109\ : LocalMux
    port map (
            O => \N__21534\,
            I => \N__21512\
        );

    \I__5108\ : InMux
    port map (
            O => \N__21533\,
            I => \N__21507\
        );

    \I__5107\ : InMux
    port map (
            O => \N__21532\,
            I => \N__21507\
        );

    \I__5106\ : InMux
    port map (
            O => \N__21531\,
            I => \N__21500\
        );

    \I__5105\ : InMux
    port map (
            O => \N__21530\,
            I => \N__21500\
        );

    \I__5104\ : InMux
    port map (
            O => \N__21529\,
            I => \N__21500\
        );

    \I__5103\ : InMux
    port map (
            O => \N__21528\,
            I => \N__21495\
        );

    \I__5102\ : InMux
    port map (
            O => \N__21527\,
            I => \N__21495\
        );

    \I__5101\ : Odrv4
    port map (
            O => \N__21522\,
            I => \b2v_inst1.r_Clk_CountZ0Z_0\
        );

    \I__5100\ : LocalMux
    port map (
            O => \N__21517\,
            I => \b2v_inst1.r_Clk_CountZ0Z_0\
        );

    \I__5099\ : Odrv4
    port map (
            O => \N__21512\,
            I => \b2v_inst1.r_Clk_CountZ0Z_0\
        );

    \I__5098\ : LocalMux
    port map (
            O => \N__21507\,
            I => \b2v_inst1.r_Clk_CountZ0Z_0\
        );

    \I__5097\ : LocalMux
    port map (
            O => \N__21500\,
            I => \b2v_inst1.r_Clk_CountZ0Z_0\
        );

    \I__5096\ : LocalMux
    port map (
            O => \N__21495\,
            I => \b2v_inst1.r_Clk_CountZ0Z_0\
        );

    \I__5095\ : CascadeMux
    port map (
            O => \N__21482\,
            I => \b2v_inst1.g3_1_cascade_\
        );

    \I__5094\ : InMux
    port map (
            O => \N__21479\,
            I => \N__21473\
        );

    \I__5093\ : InMux
    port map (
            O => \N__21478\,
            I => \N__21468\
        );

    \I__5092\ : InMux
    port map (
            O => \N__21477\,
            I => \N__21468\
        );

    \I__5091\ : CascadeMux
    port map (
            O => \N__21476\,
            I => \N__21464\
        );

    \I__5090\ : LocalMux
    port map (
            O => \N__21473\,
            I => \N__21457\
        );

    \I__5089\ : LocalMux
    port map (
            O => \N__21468\,
            I => \N__21457\
        );

    \I__5088\ : InMux
    port map (
            O => \N__21467\,
            I => \N__21450\
        );

    \I__5087\ : InMux
    port map (
            O => \N__21464\,
            I => \N__21445\
        );

    \I__5086\ : InMux
    port map (
            O => \N__21463\,
            I => \N__21445\
        );

    \I__5085\ : CascadeMux
    port map (
            O => \N__21462\,
            I => \N__21440\
        );

    \I__5084\ : Span4Mux_v
    port map (
            O => \N__21457\,
            I => \N__21436\
        );

    \I__5083\ : InMux
    port map (
            O => \N__21456\,
            I => \N__21431\
        );

    \I__5082\ : InMux
    port map (
            O => \N__21455\,
            I => \N__21431\
        );

    \I__5081\ : InMux
    port map (
            O => \N__21454\,
            I => \N__21426\
        );

    \I__5080\ : InMux
    port map (
            O => \N__21453\,
            I => \N__21426\
        );

    \I__5079\ : LocalMux
    port map (
            O => \N__21450\,
            I => \N__21421\
        );

    \I__5078\ : LocalMux
    port map (
            O => \N__21445\,
            I => \N__21421\
        );

    \I__5077\ : InMux
    port map (
            O => \N__21444\,
            I => \N__21416\
        );

    \I__5076\ : InMux
    port map (
            O => \N__21443\,
            I => \N__21416\
        );

    \I__5075\ : InMux
    port map (
            O => \N__21440\,
            I => \N__21411\
        );

    \I__5074\ : InMux
    port map (
            O => \N__21439\,
            I => \N__21411\
        );

    \I__5073\ : Span4Mux_h
    port map (
            O => \N__21436\,
            I => \N__21404\
        );

    \I__5072\ : LocalMux
    port map (
            O => \N__21431\,
            I => \N__21404\
        );

    \I__5071\ : LocalMux
    port map (
            O => \N__21426\,
            I => \N__21404\
        );

    \I__5070\ : Odrv4
    port map (
            O => \N__21421\,
            I => \b2v_inst1.r_Clk_CountZ0Z_1\
        );

    \I__5069\ : LocalMux
    port map (
            O => \N__21416\,
            I => \b2v_inst1.r_Clk_CountZ0Z_1\
        );

    \I__5068\ : LocalMux
    port map (
            O => \N__21411\,
            I => \b2v_inst1.r_Clk_CountZ0Z_1\
        );

    \I__5067\ : Odrv4
    port map (
            O => \N__21404\,
            I => \b2v_inst1.r_Clk_CountZ0Z_1\
        );

    \I__5066\ : InMux
    port map (
            O => \N__21395\,
            I => \N__21392\
        );

    \I__5065\ : LocalMux
    port map (
            O => \N__21392\,
            I => \N__21389\
        );

    \I__5064\ : Odrv4
    port map (
            O => \N__21389\,
            I => \b2v_inst1.g3\
        );

    \I__5063\ : InMux
    port map (
            O => \N__21386\,
            I => \N__21383\
        );

    \I__5062\ : LocalMux
    port map (
            O => \N__21383\,
            I => \N__21380\
        );

    \I__5061\ : Odrv4
    port map (
            O => \N__21380\,
            I => \b2v_inst1.N_9_0\
        );

    \I__5060\ : CascadeMux
    port map (
            O => \N__21377\,
            I => \b2v_inst1.N_13_cascade_\
        );

    \I__5059\ : InMux
    port map (
            O => \N__21374\,
            I => \N__21371\
        );

    \I__5058\ : LocalMux
    port map (
            O => \N__21371\,
            I => \N__21368\
        );

    \I__5057\ : Span4Mux_h
    port map (
            O => \N__21368\,
            I => \N__21365\
        );

    \I__5056\ : Odrv4
    port map (
            O => \N__21365\,
            I => \b2v_inst1.g0_0_i_a6_3_0\
        );

    \I__5055\ : CascadeMux
    port map (
            O => \N__21362\,
            I => \b2v_inst1.g0_1_4_cascade_\
        );

    \I__5054\ : InMux
    port map (
            O => \N__21359\,
            I => \N__21356\
        );

    \I__5053\ : LocalMux
    port map (
            O => \N__21356\,
            I => \N__21348\
        );

    \I__5052\ : CascadeMux
    port map (
            O => \N__21355\,
            I => \N__21345\
        );

    \I__5051\ : CascadeMux
    port map (
            O => \N__21354\,
            I => \N__21342\
        );

    \I__5050\ : InMux
    port map (
            O => \N__21353\,
            I => \N__21339\
        );

    \I__5049\ : InMux
    port map (
            O => \N__21352\,
            I => \N__21336\
        );

    \I__5048\ : InMux
    port map (
            O => \N__21351\,
            I => \N__21333\
        );

    \I__5047\ : Span4Mux_h
    port map (
            O => \N__21348\,
            I => \N__21330\
        );

    \I__5046\ : InMux
    port map (
            O => \N__21345\,
            I => \N__21327\
        );

    \I__5045\ : InMux
    port map (
            O => \N__21342\,
            I => \N__21324\
        );

    \I__5044\ : LocalMux
    port map (
            O => \N__21339\,
            I => \b2v_inst1.N_28_mux\
        );

    \I__5043\ : LocalMux
    port map (
            O => \N__21336\,
            I => \b2v_inst1.N_28_mux\
        );

    \I__5042\ : LocalMux
    port map (
            O => \N__21333\,
            I => \b2v_inst1.N_28_mux\
        );

    \I__5041\ : Odrv4
    port map (
            O => \N__21330\,
            I => \b2v_inst1.N_28_mux\
        );

    \I__5040\ : LocalMux
    port map (
            O => \N__21327\,
            I => \b2v_inst1.N_28_mux\
        );

    \I__5039\ : LocalMux
    port map (
            O => \N__21324\,
            I => \b2v_inst1.N_28_mux\
        );

    \I__5038\ : InMux
    port map (
            O => \N__21311\,
            I => \N__21305\
        );

    \I__5037\ : InMux
    port map (
            O => \N__21310\,
            I => \N__21305\
        );

    \I__5036\ : LocalMux
    port map (
            O => \N__21305\,
            I => \N__21302\
        );

    \I__5035\ : Odrv4
    port map (
            O => \N__21302\,
            I => \b2v_inst1.un1_r_SM_Main_3_0\
        );

    \I__5034\ : CascadeMux
    port map (
            O => \N__21299\,
            I => \b2v_inst1.g0_1_cascade_\
        );

    \I__5033\ : InMux
    port map (
            O => \N__21296\,
            I => \N__21293\
        );

    \I__5032\ : LocalMux
    port map (
            O => \N__21293\,
            I => \b2v_inst1.N_29_mux_1\
        );

    \I__5031\ : CascadeMux
    port map (
            O => \N__21290\,
            I => \b2v_inst1.N_14_0_1_cascade_\
        );

    \I__5030\ : CascadeMux
    port map (
            O => \N__21287\,
            I => \b2v_inst1.g0_0_i_a6_1_5_cascade_\
        );

    \I__5029\ : InMux
    port map (
            O => \N__21284\,
            I => \N__21281\
        );

    \I__5028\ : LocalMux
    port map (
            O => \N__21281\,
            I => \b2v_inst1.g0_0_i_a6_1_1\
        );

    \I__5027\ : CascadeMux
    port map (
            O => \N__21278\,
            I => \N__21275\
        );

    \I__5026\ : InMux
    port map (
            O => \N__21275\,
            I => \N__21272\
        );

    \I__5025\ : LocalMux
    port map (
            O => \N__21272\,
            I => \b2v_inst1.un1_r_Clk_Count_ac0_3_out\
        );

    \I__5024\ : CascadeMux
    port map (
            O => \N__21269\,
            I => \b2v_inst.un8_dir_mem_3_ac0_9_0_cascade_\
        );

    \I__5023\ : InMux
    port map (
            O => \N__21266\,
            I => \N__21262\
        );

    \I__5022\ : InMux
    port map (
            O => \N__21265\,
            I => \N__21258\
        );

    \I__5021\ : LocalMux
    port map (
            O => \N__21262\,
            I => \N__21255\
        );

    \I__5020\ : InMux
    port map (
            O => \N__21261\,
            I => \N__21252\
        );

    \I__5019\ : LocalMux
    port map (
            O => \N__21258\,
            I => \N__21248\
        );

    \I__5018\ : Span4Mux_v
    port map (
            O => \N__21255\,
            I => \N__21243\
        );

    \I__5017\ : LocalMux
    port map (
            O => \N__21252\,
            I => \N__21243\
        );

    \I__5016\ : InMux
    port map (
            O => \N__21251\,
            I => \N__21240\
        );

    \I__5015\ : Odrv4
    port map (
            O => \N__21248\,
            I => \b2v_inst.un10_indice\
        );

    \I__5014\ : Odrv4
    port map (
            O => \N__21243\,
            I => \b2v_inst.un10_indice\
        );

    \I__5013\ : LocalMux
    port map (
            O => \N__21240\,
            I => \b2v_inst.un10_indice\
        );

    \I__5012\ : InMux
    port map (
            O => \N__21233\,
            I => \N__21229\
        );

    \I__5011\ : InMux
    port map (
            O => \N__21232\,
            I => \N__21226\
        );

    \I__5010\ : LocalMux
    port map (
            O => \N__21229\,
            I => \N__21215\
        );

    \I__5009\ : LocalMux
    port map (
            O => \N__21226\,
            I => \N__21215\
        );

    \I__5008\ : InMux
    port map (
            O => \N__21225\,
            I => \N__21210\
        );

    \I__5007\ : InMux
    port map (
            O => \N__21224\,
            I => \N__21210\
        );

    \I__5006\ : InMux
    port map (
            O => \N__21223\,
            I => \N__21207\
        );

    \I__5005\ : InMux
    port map (
            O => \N__21222\,
            I => \N__21197\
        );

    \I__5004\ : InMux
    port map (
            O => \N__21221\,
            I => \N__21197\
        );

    \I__5003\ : InMux
    port map (
            O => \N__21220\,
            I => \N__21197\
        );

    \I__5002\ : Span4Mux_h
    port map (
            O => \N__21215\,
            I => \N__21190\
        );

    \I__5001\ : LocalMux
    port map (
            O => \N__21210\,
            I => \N__21190\
        );

    \I__5000\ : LocalMux
    port map (
            O => \N__21207\,
            I => \N__21190\
        );

    \I__4999\ : InMux
    port map (
            O => \N__21206\,
            I => \N__21183\
        );

    \I__4998\ : InMux
    port map (
            O => \N__21205\,
            I => \N__21183\
        );

    \I__4997\ : InMux
    port map (
            O => \N__21204\,
            I => \N__21183\
        );

    \I__4996\ : LocalMux
    port map (
            O => \N__21197\,
            I => \b2v_inst.indice_4_repZ0Z1\
        );

    \I__4995\ : Odrv4
    port map (
            O => \N__21190\,
            I => \b2v_inst.indice_4_repZ0Z1\
        );

    \I__4994\ : LocalMux
    port map (
            O => \N__21183\,
            I => \b2v_inst.indice_4_repZ0Z1\
        );

    \I__4993\ : InMux
    port map (
            O => \N__21176\,
            I => \N__21165\
        );

    \I__4992\ : InMux
    port map (
            O => \N__21175\,
            I => \N__21165\
        );

    \I__4991\ : InMux
    port map (
            O => \N__21174\,
            I => \N__21165\
        );

    \I__4990\ : InMux
    port map (
            O => \N__21173\,
            I => \N__21162\
        );

    \I__4989\ : InMux
    port map (
            O => \N__21172\,
            I => \N__21159\
        );

    \I__4988\ : LocalMux
    port map (
            O => \N__21165\,
            I => \N__21152\
        );

    \I__4987\ : LocalMux
    port map (
            O => \N__21162\,
            I => \N__21147\
        );

    \I__4986\ : LocalMux
    port map (
            O => \N__21159\,
            I => \N__21147\
        );

    \I__4985\ : InMux
    port map (
            O => \N__21158\,
            I => \N__21142\
        );

    \I__4984\ : InMux
    port map (
            O => \N__21157\,
            I => \N__21135\
        );

    \I__4983\ : InMux
    port map (
            O => \N__21156\,
            I => \N__21135\
        );

    \I__4982\ : InMux
    port map (
            O => \N__21155\,
            I => \N__21135\
        );

    \I__4981\ : Span4Mux_v
    port map (
            O => \N__21152\,
            I => \N__21128\
        );

    \I__4980\ : Span4Mux_h
    port map (
            O => \N__21147\,
            I => \N__21128\
        );

    \I__4979\ : InMux
    port map (
            O => \N__21146\,
            I => \N__21125\
        );

    \I__4978\ : InMux
    port map (
            O => \N__21145\,
            I => \N__21122\
        );

    \I__4977\ : LocalMux
    port map (
            O => \N__21142\,
            I => \N__21119\
        );

    \I__4976\ : LocalMux
    port map (
            O => \N__21135\,
            I => \N__21116\
        );

    \I__4975\ : InMux
    port map (
            O => \N__21134\,
            I => \N__21111\
        );

    \I__4974\ : InMux
    port map (
            O => \N__21133\,
            I => \N__21111\
        );

    \I__4973\ : Span4Mux_v
    port map (
            O => \N__21128\,
            I => \N__21106\
        );

    \I__4972\ : LocalMux
    port map (
            O => \N__21125\,
            I => \N__21106\
        );

    \I__4971\ : LocalMux
    port map (
            O => \N__21122\,
            I => \b2v_inst.indice_1_repZ0Z2\
        );

    \I__4970\ : Odrv12
    port map (
            O => \N__21119\,
            I => \b2v_inst.indice_1_repZ0Z2\
        );

    \I__4969\ : Odrv4
    port map (
            O => \N__21116\,
            I => \b2v_inst.indice_1_repZ0Z2\
        );

    \I__4968\ : LocalMux
    port map (
            O => \N__21111\,
            I => \b2v_inst.indice_1_repZ0Z2\
        );

    \I__4967\ : Odrv4
    port map (
            O => \N__21106\,
            I => \b2v_inst.indice_1_repZ0Z2\
        );

    \I__4966\ : CascadeMux
    port map (
            O => \N__21095\,
            I => \N__21087\
        );

    \I__4965\ : InMux
    port map (
            O => \N__21094\,
            I => \N__21080\
        );

    \I__4964\ : InMux
    port map (
            O => \N__21093\,
            I => \N__21077\
        );

    \I__4963\ : InMux
    port map (
            O => \N__21092\,
            I => \N__21072\
        );

    \I__4962\ : InMux
    port map (
            O => \N__21091\,
            I => \N__21072\
        );

    \I__4961\ : InMux
    port map (
            O => \N__21090\,
            I => \N__21069\
        );

    \I__4960\ : InMux
    port map (
            O => \N__21087\,
            I => \N__21066\
        );

    \I__4959\ : InMux
    port map (
            O => \N__21086\,
            I => \N__21063\
        );

    \I__4958\ : CascadeMux
    port map (
            O => \N__21085\,
            I => \N__21060\
        );

    \I__4957\ : InMux
    port map (
            O => \N__21084\,
            I => \N__21053\
        );

    \I__4956\ : InMux
    port map (
            O => \N__21083\,
            I => \N__21053\
        );

    \I__4955\ : LocalMux
    port map (
            O => \N__21080\,
            I => \N__21046\
        );

    \I__4954\ : LocalMux
    port map (
            O => \N__21077\,
            I => \N__21046\
        );

    \I__4953\ : LocalMux
    port map (
            O => \N__21072\,
            I => \N__21046\
        );

    \I__4952\ : LocalMux
    port map (
            O => \N__21069\,
            I => \N__21039\
        );

    \I__4951\ : LocalMux
    port map (
            O => \N__21066\,
            I => \N__21039\
        );

    \I__4950\ : LocalMux
    port map (
            O => \N__21063\,
            I => \N__21039\
        );

    \I__4949\ : InMux
    port map (
            O => \N__21060\,
            I => \N__21035\
        );

    \I__4948\ : InMux
    port map (
            O => \N__21059\,
            I => \N__21032\
        );

    \I__4947\ : InMux
    port map (
            O => \N__21058\,
            I => \N__21029\
        );

    \I__4946\ : LocalMux
    port map (
            O => \N__21053\,
            I => \N__21024\
        );

    \I__4945\ : Span4Mux_v
    port map (
            O => \N__21046\,
            I => \N__21024\
        );

    \I__4944\ : Span4Mux_v
    port map (
            O => \N__21039\,
            I => \N__21021\
        );

    \I__4943\ : InMux
    port map (
            O => \N__21038\,
            I => \N__21018\
        );

    \I__4942\ : LocalMux
    port map (
            O => \N__21035\,
            I => \b2v_inst.indice_0_repZ0Z2\
        );

    \I__4941\ : LocalMux
    port map (
            O => \N__21032\,
            I => \b2v_inst.indice_0_repZ0Z2\
        );

    \I__4940\ : LocalMux
    port map (
            O => \N__21029\,
            I => \b2v_inst.indice_0_repZ0Z2\
        );

    \I__4939\ : Odrv4
    port map (
            O => \N__21024\,
            I => \b2v_inst.indice_0_repZ0Z2\
        );

    \I__4938\ : Odrv4
    port map (
            O => \N__21021\,
            I => \b2v_inst.indice_0_repZ0Z2\
        );

    \I__4937\ : LocalMux
    port map (
            O => \N__21018\,
            I => \b2v_inst.indice_0_repZ0Z2\
        );

    \I__4936\ : InMux
    port map (
            O => \N__21005\,
            I => \N__20997\
        );

    \I__4935\ : InMux
    port map (
            O => \N__21004\,
            I => \N__20997\
        );

    \I__4934\ : InMux
    port map (
            O => \N__21003\,
            I => \N__20994\
        );

    \I__4933\ : CascadeMux
    port map (
            O => \N__21002\,
            I => \N__20991\
        );

    \I__4932\ : LocalMux
    port map (
            O => \N__20997\,
            I => \N__20987\
        );

    \I__4931\ : LocalMux
    port map (
            O => \N__20994\,
            I => \N__20984\
        );

    \I__4930\ : InMux
    port map (
            O => \N__20991\,
            I => \N__20981\
        );

    \I__4929\ : InMux
    port map (
            O => \N__20990\,
            I => \N__20978\
        );

    \I__4928\ : Span4Mux_h
    port map (
            O => \N__20987\,
            I => \N__20975\
        );

    \I__4927\ : Span4Mux_h
    port map (
            O => \N__20984\,
            I => \N__20972\
        );

    \I__4926\ : LocalMux
    port map (
            O => \N__20981\,
            I => \N__20969\
        );

    \I__4925\ : LocalMux
    port map (
            O => \N__20978\,
            I => \N__20966\
        );

    \I__4924\ : Odrv4
    port map (
            O => \N__20975\,
            I => \b2v_inst.un10_indice_2_0\
        );

    \I__4923\ : Odrv4
    port map (
            O => \N__20972\,
            I => \b2v_inst.un10_indice_2_0\
        );

    \I__4922\ : Odrv4
    port map (
            O => \N__20969\,
            I => \b2v_inst.un10_indice_2_0\
        );

    \I__4921\ : Odrv4
    port map (
            O => \N__20966\,
            I => \b2v_inst.un10_indice_2_0\
        );

    \I__4920\ : InMux
    port map (
            O => \N__20957\,
            I => \N__20954\
        );

    \I__4919\ : LocalMux
    port map (
            O => \N__20954\,
            I => \N__20950\
        );

    \I__4918\ : CascadeMux
    port map (
            O => \N__20953\,
            I => \N__20947\
        );

    \I__4917\ : Span4Mux_h
    port map (
            O => \N__20950\,
            I => \N__20944\
        );

    \I__4916\ : InMux
    port map (
            O => \N__20947\,
            I => \N__20941\
        );

    \I__4915\ : Odrv4
    port map (
            O => \N__20944\,
            I => \b2v_inst.un8_dir_mem_3_ac0_9_0\
        );

    \I__4914\ : LocalMux
    port map (
            O => \N__20941\,
            I => \b2v_inst.un8_dir_mem_3_ac0_9_0\
        );

    \I__4913\ : InMux
    port map (
            O => \N__20936\,
            I => \N__20929\
        );

    \I__4912\ : InMux
    port map (
            O => \N__20935\,
            I => \N__20924\
        );

    \I__4911\ : InMux
    port map (
            O => \N__20934\,
            I => \N__20921\
        );

    \I__4910\ : InMux
    port map (
            O => \N__20933\,
            I => \N__20918\
        );

    \I__4909\ : InMux
    port map (
            O => \N__20932\,
            I => \N__20915\
        );

    \I__4908\ : LocalMux
    port map (
            O => \N__20929\,
            I => \N__20909\
        );

    \I__4907\ : InMux
    port map (
            O => \N__20928\,
            I => \N__20906\
        );

    \I__4906\ : InMux
    port map (
            O => \N__20927\,
            I => \N__20903\
        );

    \I__4905\ : LocalMux
    port map (
            O => \N__20924\,
            I => \N__20900\
        );

    \I__4904\ : LocalMux
    port map (
            O => \N__20921\,
            I => \N__20890\
        );

    \I__4903\ : LocalMux
    port map (
            O => \N__20918\,
            I => \N__20890\
        );

    \I__4902\ : LocalMux
    port map (
            O => \N__20915\,
            I => \N__20890\
        );

    \I__4901\ : InMux
    port map (
            O => \N__20914\,
            I => \N__20883\
        );

    \I__4900\ : InMux
    port map (
            O => \N__20913\,
            I => \N__20883\
        );

    \I__4899\ : InMux
    port map (
            O => \N__20912\,
            I => \N__20883\
        );

    \I__4898\ : Span4Mux_v
    port map (
            O => \N__20909\,
            I => \N__20878\
        );

    \I__4897\ : LocalMux
    port map (
            O => \N__20906\,
            I => \N__20878\
        );

    \I__4896\ : LocalMux
    port map (
            O => \N__20903\,
            I => \N__20873\
        );

    \I__4895\ : Span4Mux_h
    port map (
            O => \N__20900\,
            I => \N__20873\
        );

    \I__4894\ : CascadeMux
    port map (
            O => \N__20899\,
            I => \N__20869\
        );

    \I__4893\ : InMux
    port map (
            O => \N__20898\,
            I => \N__20862\
        );

    \I__4892\ : InMux
    port map (
            O => \N__20897\,
            I => \N__20862\
        );

    \I__4891\ : Span4Mux_v
    port map (
            O => \N__20890\,
            I => \N__20857\
        );

    \I__4890\ : LocalMux
    port map (
            O => \N__20883\,
            I => \N__20857\
        );

    \I__4889\ : Span4Mux_h
    port map (
            O => \N__20878\,
            I => \N__20852\
        );

    \I__4888\ : Span4Mux_v
    port map (
            O => \N__20873\,
            I => \N__20852\
        );

    \I__4887\ : InMux
    port map (
            O => \N__20872\,
            I => \N__20847\
        );

    \I__4886\ : InMux
    port map (
            O => \N__20869\,
            I => \N__20847\
        );

    \I__4885\ : InMux
    port map (
            O => \N__20868\,
            I => \N__20842\
        );

    \I__4884\ : InMux
    port map (
            O => \N__20867\,
            I => \N__20842\
        );

    \I__4883\ : LocalMux
    port map (
            O => \N__20862\,
            I => \b2v_inst.indiceZ0Z_7\
        );

    \I__4882\ : Odrv4
    port map (
            O => \N__20857\,
            I => \b2v_inst.indiceZ0Z_7\
        );

    \I__4881\ : Odrv4
    port map (
            O => \N__20852\,
            I => \b2v_inst.indiceZ0Z_7\
        );

    \I__4880\ : LocalMux
    port map (
            O => \N__20847\,
            I => \b2v_inst.indiceZ0Z_7\
        );

    \I__4879\ : LocalMux
    port map (
            O => \N__20842\,
            I => \b2v_inst.indiceZ0Z_7\
        );

    \I__4878\ : CascadeMux
    port map (
            O => \N__20831\,
            I => \N__20828\
        );

    \I__4877\ : InMux
    port map (
            O => \N__20828\,
            I => \N__20815\
        );

    \I__4876\ : InMux
    port map (
            O => \N__20827\,
            I => \N__20815\
        );

    \I__4875\ : InMux
    port map (
            O => \N__20826\,
            I => \N__20815\
        );

    \I__4874\ : InMux
    port map (
            O => \N__20825\,
            I => \N__20812\
        );

    \I__4873\ : InMux
    port map (
            O => \N__20824\,
            I => \N__20809\
        );

    \I__4872\ : InMux
    port map (
            O => \N__20823\,
            I => \N__20804\
        );

    \I__4871\ : InMux
    port map (
            O => \N__20822\,
            I => \N__20804\
        );

    \I__4870\ : LocalMux
    port map (
            O => \N__20815\,
            I => \N__20801\
        );

    \I__4869\ : LocalMux
    port map (
            O => \N__20812\,
            I => \N__20798\
        );

    \I__4868\ : LocalMux
    port map (
            O => \N__20809\,
            I => \N__20792\
        );

    \I__4867\ : LocalMux
    port map (
            O => \N__20804\,
            I => \N__20792\
        );

    \I__4866\ : Span4Mux_v
    port map (
            O => \N__20801\,
            I => \N__20789\
        );

    \I__4865\ : Span4Mux_h
    port map (
            O => \N__20798\,
            I => \N__20786\
        );

    \I__4864\ : InMux
    port map (
            O => \N__20797\,
            I => \N__20783\
        );

    \I__4863\ : Span4Mux_v
    port map (
            O => \N__20792\,
            I => \N__20780\
        );

    \I__4862\ : Span4Mux_h
    port map (
            O => \N__20789\,
            I => \N__20777\
        );

    \I__4861\ : Odrv4
    port map (
            O => \N__20786\,
            I => \b2v_inst.un8_dir_mem_3_c4\
        );

    \I__4860\ : LocalMux
    port map (
            O => \N__20783\,
            I => \b2v_inst.un8_dir_mem_3_c4\
        );

    \I__4859\ : Odrv4
    port map (
            O => \N__20780\,
            I => \b2v_inst.un8_dir_mem_3_c4\
        );

    \I__4858\ : Odrv4
    port map (
            O => \N__20777\,
            I => \b2v_inst.un8_dir_mem_3_c4\
        );

    \I__4857\ : CascadeMux
    port map (
            O => \N__20768\,
            I => \N__20765\
        );

    \I__4856\ : InMux
    port map (
            O => \N__20765\,
            I => \N__20760\
        );

    \I__4855\ : CascadeMux
    port map (
            O => \N__20764\,
            I => \N__20757\
        );

    \I__4854\ : CascadeMux
    port map (
            O => \N__20763\,
            I => \N__20751\
        );

    \I__4853\ : LocalMux
    port map (
            O => \N__20760\,
            I => \N__20748\
        );

    \I__4852\ : InMux
    port map (
            O => \N__20757\,
            I => \N__20745\
        );

    \I__4851\ : InMux
    port map (
            O => \N__20756\,
            I => \N__20742\
        );

    \I__4850\ : InMux
    port map (
            O => \N__20755\,
            I => \N__20737\
        );

    \I__4849\ : InMux
    port map (
            O => \N__20754\,
            I => \N__20737\
        );

    \I__4848\ : InMux
    port map (
            O => \N__20751\,
            I => \N__20734\
        );

    \I__4847\ : Odrv4
    port map (
            O => \N__20748\,
            I => \b2v_inst.indice_fastZ0Z_4\
        );

    \I__4846\ : LocalMux
    port map (
            O => \N__20745\,
            I => \b2v_inst.indice_fastZ0Z_4\
        );

    \I__4845\ : LocalMux
    port map (
            O => \N__20742\,
            I => \b2v_inst.indice_fastZ0Z_4\
        );

    \I__4844\ : LocalMux
    port map (
            O => \N__20737\,
            I => \b2v_inst.indice_fastZ0Z_4\
        );

    \I__4843\ : LocalMux
    port map (
            O => \N__20734\,
            I => \b2v_inst.indice_fastZ0Z_4\
        );

    \I__4842\ : InMux
    port map (
            O => \N__20723\,
            I => \N__20719\
        );

    \I__4841\ : InMux
    port map (
            O => \N__20722\,
            I => \N__20716\
        );

    \I__4840\ : LocalMux
    port map (
            O => \N__20719\,
            I => \N__20713\
        );

    \I__4839\ : LocalMux
    port map (
            O => \N__20716\,
            I => \N__20707\
        );

    \I__4838\ : Span4Mux_h
    port map (
            O => \N__20713\,
            I => \N__20704\
        );

    \I__4837\ : InMux
    port map (
            O => \N__20712\,
            I => \N__20699\
        );

    \I__4836\ : InMux
    port map (
            O => \N__20711\,
            I => \N__20699\
        );

    \I__4835\ : InMux
    port map (
            O => \N__20710\,
            I => \N__20696\
        );

    \I__4834\ : Odrv12
    port map (
            O => \N__20707\,
            I => \b2v_inst.indice_fastZ0Z_3\
        );

    \I__4833\ : Odrv4
    port map (
            O => \N__20704\,
            I => \b2v_inst.indice_fastZ0Z_3\
        );

    \I__4832\ : LocalMux
    port map (
            O => \N__20699\,
            I => \b2v_inst.indice_fastZ0Z_3\
        );

    \I__4831\ : LocalMux
    port map (
            O => \N__20696\,
            I => \b2v_inst.indice_fastZ0Z_3\
        );

    \I__4830\ : InMux
    port map (
            O => \N__20687\,
            I => \N__20682\
        );

    \I__4829\ : InMux
    port map (
            O => \N__20686\,
            I => \N__20677\
        );

    \I__4828\ : InMux
    port map (
            O => \N__20685\,
            I => \N__20677\
        );

    \I__4827\ : LocalMux
    port map (
            O => \N__20682\,
            I => \N__20674\
        );

    \I__4826\ : LocalMux
    port map (
            O => \N__20677\,
            I => \N__20671\
        );

    \I__4825\ : Odrv12
    port map (
            O => \N__20674\,
            I => \b2v_inst.un8_dir_mem_1_ac0_7_out\
        );

    \I__4824\ : Odrv4
    port map (
            O => \N__20671\,
            I => \b2v_inst.un8_dir_mem_1_ac0_7_out\
        );

    \I__4823\ : CascadeMux
    port map (
            O => \N__20666\,
            I => \N__20661\
        );

    \I__4822\ : InMux
    port map (
            O => \N__20665\,
            I => \N__20658\
        );

    \I__4821\ : InMux
    port map (
            O => \N__20664\,
            I => \N__20653\
        );

    \I__4820\ : InMux
    port map (
            O => \N__20661\,
            I => \N__20653\
        );

    \I__4819\ : LocalMux
    port map (
            O => \N__20658\,
            I => \N__20650\
        );

    \I__4818\ : LocalMux
    port map (
            O => \N__20653\,
            I => \N__20647\
        );

    \I__4817\ : Span4Mux_v
    port map (
            O => \N__20650\,
            I => \N__20642\
        );

    \I__4816\ : Span4Mux_v
    port map (
            O => \N__20647\,
            I => \N__20642\
        );

    \I__4815\ : Odrv4
    port map (
            O => \N__20642\,
            I => \b2v_inst.un8_dir_mem_2_c4\
        );

    \I__4814\ : InMux
    port map (
            O => \N__20639\,
            I => \N__20627\
        );

    \I__4813\ : InMux
    port map (
            O => \N__20638\,
            I => \N__20624\
        );

    \I__4812\ : InMux
    port map (
            O => \N__20637\,
            I => \N__20621\
        );

    \I__4811\ : InMux
    port map (
            O => \N__20636\,
            I => \N__20618\
        );

    \I__4810\ : InMux
    port map (
            O => \N__20635\,
            I => \N__20614\
        );

    \I__4809\ : InMux
    port map (
            O => \N__20634\,
            I => \N__20611\
        );

    \I__4808\ : InMux
    port map (
            O => \N__20633\,
            I => \N__20605\
        );

    \I__4807\ : InMux
    port map (
            O => \N__20632\,
            I => \N__20605\
        );

    \I__4806\ : InMux
    port map (
            O => \N__20631\,
            I => \N__20600\
        );

    \I__4805\ : InMux
    port map (
            O => \N__20630\,
            I => \N__20597\
        );

    \I__4804\ : LocalMux
    port map (
            O => \N__20627\,
            I => \N__20588\
        );

    \I__4803\ : LocalMux
    port map (
            O => \N__20624\,
            I => \N__20588\
        );

    \I__4802\ : LocalMux
    port map (
            O => \N__20621\,
            I => \N__20588\
        );

    \I__4801\ : LocalMux
    port map (
            O => \N__20618\,
            I => \N__20588\
        );

    \I__4800\ : InMux
    port map (
            O => \N__20617\,
            I => \N__20585\
        );

    \I__4799\ : LocalMux
    port map (
            O => \N__20614\,
            I => \N__20580\
        );

    \I__4798\ : LocalMux
    port map (
            O => \N__20611\,
            I => \N__20580\
        );

    \I__4797\ : InMux
    port map (
            O => \N__20610\,
            I => \N__20573\
        );

    \I__4796\ : LocalMux
    port map (
            O => \N__20605\,
            I => \N__20570\
        );

    \I__4795\ : InMux
    port map (
            O => \N__20604\,
            I => \N__20565\
        );

    \I__4794\ : InMux
    port map (
            O => \N__20603\,
            I => \N__20565\
        );

    \I__4793\ : LocalMux
    port map (
            O => \N__20600\,
            I => \N__20562\
        );

    \I__4792\ : LocalMux
    port map (
            O => \N__20597\,
            I => \N__20558\
        );

    \I__4791\ : Span4Mux_v
    port map (
            O => \N__20588\,
            I => \N__20550\
        );

    \I__4790\ : LocalMux
    port map (
            O => \N__20585\,
            I => \N__20550\
        );

    \I__4789\ : Span4Mux_v
    port map (
            O => \N__20580\,
            I => \N__20550\
        );

    \I__4788\ : InMux
    port map (
            O => \N__20579\,
            I => \N__20547\
        );

    \I__4787\ : InMux
    port map (
            O => \N__20578\,
            I => \N__20540\
        );

    \I__4786\ : InMux
    port map (
            O => \N__20577\,
            I => \N__20540\
        );

    \I__4785\ : InMux
    port map (
            O => \N__20576\,
            I => \N__20540\
        );

    \I__4784\ : LocalMux
    port map (
            O => \N__20573\,
            I => \N__20531\
        );

    \I__4783\ : Span12Mux_s11_v
    port map (
            O => \N__20570\,
            I => \N__20531\
        );

    \I__4782\ : LocalMux
    port map (
            O => \N__20565\,
            I => \N__20531\
        );

    \I__4781\ : Span12Mux_v
    port map (
            O => \N__20562\,
            I => \N__20531\
        );

    \I__4780\ : InMux
    port map (
            O => \N__20561\,
            I => \N__20528\
        );

    \I__4779\ : Span4Mux_v
    port map (
            O => \N__20558\,
            I => \N__20525\
        );

    \I__4778\ : InMux
    port map (
            O => \N__20557\,
            I => \N__20522\
        );

    \I__4777\ : Span4Mux_h
    port map (
            O => \N__20550\,
            I => \N__20519\
        );

    \I__4776\ : LocalMux
    port map (
            O => \N__20547\,
            I => \b2v_inst.indiceZ0Z_6\
        );

    \I__4775\ : LocalMux
    port map (
            O => \N__20540\,
            I => \b2v_inst.indiceZ0Z_6\
        );

    \I__4774\ : Odrv12
    port map (
            O => \N__20531\,
            I => \b2v_inst.indiceZ0Z_6\
        );

    \I__4773\ : LocalMux
    port map (
            O => \N__20528\,
            I => \b2v_inst.indiceZ0Z_6\
        );

    \I__4772\ : Odrv4
    port map (
            O => \N__20525\,
            I => \b2v_inst.indiceZ0Z_6\
        );

    \I__4771\ : LocalMux
    port map (
            O => \N__20522\,
            I => \b2v_inst.indiceZ0Z_6\
        );

    \I__4770\ : Odrv4
    port map (
            O => \N__20519\,
            I => \b2v_inst.indiceZ0Z_6\
        );

    \I__4769\ : InMux
    port map (
            O => \N__20504\,
            I => \N__20495\
        );

    \I__4768\ : InMux
    port map (
            O => \N__20503\,
            I => \N__20495\
        );

    \I__4767\ : InMux
    port map (
            O => \N__20502\,
            I => \N__20489\
        );

    \I__4766\ : InMux
    port map (
            O => \N__20501\,
            I => \N__20486\
        );

    \I__4765\ : CascadeMux
    port map (
            O => \N__20500\,
            I => \N__20479\
        );

    \I__4764\ : LocalMux
    port map (
            O => \N__20495\,
            I => \N__20473\
        );

    \I__4763\ : InMux
    port map (
            O => \N__20494\,
            I => \N__20468\
        );

    \I__4762\ : InMux
    port map (
            O => \N__20493\,
            I => \N__20468\
        );

    \I__4761\ : InMux
    port map (
            O => \N__20492\,
            I => \N__20465\
        );

    \I__4760\ : LocalMux
    port map (
            O => \N__20489\,
            I => \N__20462\
        );

    \I__4759\ : LocalMux
    port map (
            O => \N__20486\,
            I => \N__20459\
        );

    \I__4758\ : InMux
    port map (
            O => \N__20485\,
            I => \N__20454\
        );

    \I__4757\ : InMux
    port map (
            O => \N__20484\,
            I => \N__20454\
        );

    \I__4756\ : InMux
    port map (
            O => \N__20483\,
            I => \N__20448\
        );

    \I__4755\ : InMux
    port map (
            O => \N__20482\,
            I => \N__20448\
        );

    \I__4754\ : InMux
    port map (
            O => \N__20479\,
            I => \N__20445\
        );

    \I__4753\ : InMux
    port map (
            O => \N__20478\,
            I => \N__20442\
        );

    \I__4752\ : InMux
    port map (
            O => \N__20477\,
            I => \N__20436\
        );

    \I__4751\ : InMux
    port map (
            O => \N__20476\,
            I => \N__20436\
        );

    \I__4750\ : Span4Mux_h
    port map (
            O => \N__20473\,
            I => \N__20425\
        );

    \I__4749\ : LocalMux
    port map (
            O => \N__20468\,
            I => \N__20425\
        );

    \I__4748\ : LocalMux
    port map (
            O => \N__20465\,
            I => \N__20425\
        );

    \I__4747\ : Span4Mux_v
    port map (
            O => \N__20462\,
            I => \N__20425\
        );

    \I__4746\ : Span4Mux_v
    port map (
            O => \N__20459\,
            I => \N__20425\
        );

    \I__4745\ : LocalMux
    port map (
            O => \N__20454\,
            I => \N__20422\
        );

    \I__4744\ : InMux
    port map (
            O => \N__20453\,
            I => \N__20419\
        );

    \I__4743\ : LocalMux
    port map (
            O => \N__20448\,
            I => \N__20416\
        );

    \I__4742\ : LocalMux
    port map (
            O => \N__20445\,
            I => \N__20411\
        );

    \I__4741\ : LocalMux
    port map (
            O => \N__20442\,
            I => \N__20411\
        );

    \I__4740\ : InMux
    port map (
            O => \N__20441\,
            I => \N__20408\
        );

    \I__4739\ : LocalMux
    port map (
            O => \N__20436\,
            I => \N__20399\
        );

    \I__4738\ : Span4Mux_v
    port map (
            O => \N__20425\,
            I => \N__20394\
        );

    \I__4737\ : Span4Mux_v
    port map (
            O => \N__20422\,
            I => \N__20394\
        );

    \I__4736\ : LocalMux
    port map (
            O => \N__20419\,
            I => \N__20391\
        );

    \I__4735\ : Span4Mux_h
    port map (
            O => \N__20416\,
            I => \N__20384\
        );

    \I__4734\ : Span4Mux_h
    port map (
            O => \N__20411\,
            I => \N__20384\
        );

    \I__4733\ : LocalMux
    port map (
            O => \N__20408\,
            I => \N__20384\
        );

    \I__4732\ : InMux
    port map (
            O => \N__20407\,
            I => \N__20375\
        );

    \I__4731\ : InMux
    port map (
            O => \N__20406\,
            I => \N__20375\
        );

    \I__4730\ : InMux
    port map (
            O => \N__20405\,
            I => \N__20375\
        );

    \I__4729\ : InMux
    port map (
            O => \N__20404\,
            I => \N__20375\
        );

    \I__4728\ : InMux
    port map (
            O => \N__20403\,
            I => \N__20370\
        );

    \I__4727\ : InMux
    port map (
            O => \N__20402\,
            I => \N__20370\
        );

    \I__4726\ : Span4Mux_h
    port map (
            O => \N__20399\,
            I => \N__20367\
        );

    \I__4725\ : Odrv4
    port map (
            O => \N__20394\,
            I => \b2v_inst.indiceZ0Z_5\
        );

    \I__4724\ : Odrv4
    port map (
            O => \N__20391\,
            I => \b2v_inst.indiceZ0Z_5\
        );

    \I__4723\ : Odrv4
    port map (
            O => \N__20384\,
            I => \b2v_inst.indiceZ0Z_5\
        );

    \I__4722\ : LocalMux
    port map (
            O => \N__20375\,
            I => \b2v_inst.indiceZ0Z_5\
        );

    \I__4721\ : LocalMux
    port map (
            O => \N__20370\,
            I => \b2v_inst.indiceZ0Z_5\
        );

    \I__4720\ : Odrv4
    port map (
            O => \N__20367\,
            I => \b2v_inst.indiceZ0Z_5\
        );

    \I__4719\ : InMux
    port map (
            O => \N__20354\,
            I => \N__20351\
        );

    \I__4718\ : LocalMux
    port map (
            O => \N__20351\,
            I => \N__20348\
        );

    \I__4717\ : Span4Mux_h
    port map (
            O => \N__20348\,
            I => \N__20345\
        );

    \I__4716\ : Span4Mux_h
    port map (
            O => \N__20345\,
            I => \N__20342\
        );

    \I__4715\ : Odrv4
    port map (
            O => \N__20342\,
            I => \b2v_inst.dir_mem_2_RNO_1Z0Z_6\
        );

    \I__4714\ : InMux
    port map (
            O => \N__20339\,
            I => \N__20336\
        );

    \I__4713\ : LocalMux
    port map (
            O => \N__20336\,
            I => \b2v_inst1.g0_i_o5_0_2\
        );

    \I__4712\ : CascadeMux
    port map (
            O => \N__20333\,
            I => \N__20320\
        );

    \I__4711\ : InMux
    port map (
            O => \N__20332\,
            I => \N__20317\
        );

    \I__4710\ : InMux
    port map (
            O => \N__20331\,
            I => \N__20312\
        );

    \I__4709\ : InMux
    port map (
            O => \N__20330\,
            I => \N__20312\
        );

    \I__4708\ : CascadeMux
    port map (
            O => \N__20329\,
            I => \N__20309\
        );

    \I__4707\ : InMux
    port map (
            O => \N__20328\,
            I => \N__20304\
        );

    \I__4706\ : InMux
    port map (
            O => \N__20327\,
            I => \N__20304\
        );

    \I__4705\ : InMux
    port map (
            O => \N__20326\,
            I => \N__20299\
        );

    \I__4704\ : InMux
    port map (
            O => \N__20325\,
            I => \N__20299\
        );

    \I__4703\ : CascadeMux
    port map (
            O => \N__20324\,
            I => \N__20291\
        );

    \I__4702\ : InMux
    port map (
            O => \N__20323\,
            I => \N__20286\
        );

    \I__4701\ : InMux
    port map (
            O => \N__20320\,
            I => \N__20286\
        );

    \I__4700\ : LocalMux
    port map (
            O => \N__20317\,
            I => \N__20281\
        );

    \I__4699\ : LocalMux
    port map (
            O => \N__20312\,
            I => \N__20281\
        );

    \I__4698\ : InMux
    port map (
            O => \N__20309\,
            I => \N__20278\
        );

    \I__4697\ : LocalMux
    port map (
            O => \N__20304\,
            I => \N__20271\
        );

    \I__4696\ : LocalMux
    port map (
            O => \N__20299\,
            I => \N__20271\
        );

    \I__4695\ : InMux
    port map (
            O => \N__20298\,
            I => \N__20266\
        );

    \I__4694\ : InMux
    port map (
            O => \N__20297\,
            I => \N__20266\
        );

    \I__4693\ : InMux
    port map (
            O => \N__20296\,
            I => \N__20257\
        );

    \I__4692\ : InMux
    port map (
            O => \N__20295\,
            I => \N__20257\
        );

    \I__4691\ : InMux
    port map (
            O => \N__20294\,
            I => \N__20257\
        );

    \I__4690\ : InMux
    port map (
            O => \N__20291\,
            I => \N__20257\
        );

    \I__4689\ : LocalMux
    port map (
            O => \N__20286\,
            I => \N__20254\
        );

    \I__4688\ : Span4Mux_h
    port map (
            O => \N__20281\,
            I => \N__20249\
        );

    \I__4687\ : LocalMux
    port map (
            O => \N__20278\,
            I => \N__20249\
        );

    \I__4686\ : InMux
    port map (
            O => \N__20277\,
            I => \N__20246\
        );

    \I__4685\ : CascadeMux
    port map (
            O => \N__20276\,
            I => \N__20243\
        );

    \I__4684\ : Span4Mux_v
    port map (
            O => \N__20271\,
            I => \N__20239\
        );

    \I__4683\ : LocalMux
    port map (
            O => \N__20266\,
            I => \N__20234\
        );

    \I__4682\ : LocalMux
    port map (
            O => \N__20257\,
            I => \N__20234\
        );

    \I__4681\ : Span4Mux_v
    port map (
            O => \N__20254\,
            I => \N__20227\
        );

    \I__4680\ : Span4Mux_v
    port map (
            O => \N__20249\,
            I => \N__20227\
        );

    \I__4679\ : LocalMux
    port map (
            O => \N__20246\,
            I => \N__20227\
        );

    \I__4678\ : InMux
    port map (
            O => \N__20243\,
            I => \N__20222\
        );

    \I__4677\ : InMux
    port map (
            O => \N__20242\,
            I => \N__20222\
        );

    \I__4676\ : Odrv4
    port map (
            O => \N__20239\,
            I => \b2v_inst.indiceZ0Z_3\
        );

    \I__4675\ : Odrv12
    port map (
            O => \N__20234\,
            I => \b2v_inst.indiceZ0Z_3\
        );

    \I__4674\ : Odrv4
    port map (
            O => \N__20227\,
            I => \b2v_inst.indiceZ0Z_3\
        );

    \I__4673\ : LocalMux
    port map (
            O => \N__20222\,
            I => \b2v_inst.indiceZ0Z_3\
        );

    \I__4672\ : CascadeMux
    port map (
            O => \N__20213\,
            I => \b2v_inst.dir_mem_1_RNO_0Z0Z_3_cascade_\
        );

    \I__4671\ : CascadeMux
    port map (
            O => \N__20210\,
            I => \N__20207\
        );

    \I__4670\ : InMux
    port map (
            O => \N__20207\,
            I => \N__20204\
        );

    \I__4669\ : LocalMux
    port map (
            O => \N__20204\,
            I => \N__20201\
        );

    \I__4668\ : Odrv12
    port map (
            O => \N__20201\,
            I => \b2v_inst.dir_mem_1Z0Z_3\
        );

    \I__4667\ : InMux
    port map (
            O => \N__20198\,
            I => \N__20195\
        );

    \I__4666\ : LocalMux
    port map (
            O => \N__20195\,
            I => \b2v_inst.indice_fast_RNIF91EZ0Z_0\
        );

    \I__4665\ : InMux
    port map (
            O => \N__20192\,
            I => \N__20189\
        );

    \I__4664\ : LocalMux
    port map (
            O => \N__20189\,
            I => \b2v_inst.dir_mem_115lto8_1\
        );

    \I__4663\ : InMux
    port map (
            O => \N__20186\,
            I => \N__20183\
        );

    \I__4662\ : LocalMux
    port map (
            O => \N__20183\,
            I => \b2v_inst.dir_mem_115lto6_1\
        );

    \I__4661\ : InMux
    port map (
            O => \N__20180\,
            I => \N__20176\
        );

    \I__4660\ : InMux
    port map (
            O => \N__20179\,
            I => \N__20173\
        );

    \I__4659\ : LocalMux
    port map (
            O => \N__20176\,
            I => \b2v_inst.un8_dir_mem_1_c7\
        );

    \I__4658\ : LocalMux
    port map (
            O => \N__20173\,
            I => \b2v_inst.un8_dir_mem_1_c7\
        );

    \I__4657\ : CascadeMux
    port map (
            O => \N__20168\,
            I => \b2v_inst.dir_mem_115lto8_1_cascade_\
        );

    \I__4656\ : CascadeMux
    port map (
            O => \N__20165\,
            I => \b2v_inst.dir_mem_115_0_cascade_\
        );

    \I__4655\ : InMux
    port map (
            O => \N__20162\,
            I => \N__20159\
        );

    \I__4654\ : LocalMux
    port map (
            O => \N__20159\,
            I => \N__20156\
        );

    \I__4653\ : Span4Mux_v
    port map (
            O => \N__20156\,
            I => \N__20153\
        );

    \I__4652\ : Span4Mux_h
    port map (
            O => \N__20153\,
            I => \N__20150\
        );

    \I__4651\ : Odrv4
    port map (
            O => \N__20150\,
            I => \b2v_inst.dir_mem_1Z0Z_0\
        );

    \I__4650\ : InMux
    port map (
            O => \N__20147\,
            I => \N__20143\
        );

    \I__4649\ : CascadeMux
    port map (
            O => \N__20146\,
            I => \N__20136\
        );

    \I__4648\ : LocalMux
    port map (
            O => \N__20143\,
            I => \N__20133\
        );

    \I__4647\ : InMux
    port map (
            O => \N__20142\,
            I => \N__20128\
        );

    \I__4646\ : InMux
    port map (
            O => \N__20141\,
            I => \N__20128\
        );

    \I__4645\ : InMux
    port map (
            O => \N__20140\,
            I => \N__20125\
        );

    \I__4644\ : InMux
    port map (
            O => \N__20139\,
            I => \N__20118\
        );

    \I__4643\ : InMux
    port map (
            O => \N__20136\,
            I => \N__20118\
        );

    \I__4642\ : Span4Mux_v
    port map (
            O => \N__20133\,
            I => \N__20110\
        );

    \I__4641\ : LocalMux
    port map (
            O => \N__20128\,
            I => \N__20107\
        );

    \I__4640\ : LocalMux
    port map (
            O => \N__20125\,
            I => \N__20103\
        );

    \I__4639\ : InMux
    port map (
            O => \N__20124\,
            I => \N__20098\
        );

    \I__4638\ : InMux
    port map (
            O => \N__20123\,
            I => \N__20098\
        );

    \I__4637\ : LocalMux
    port map (
            O => \N__20118\,
            I => \N__20090\
        );

    \I__4636\ : InMux
    port map (
            O => \N__20117\,
            I => \N__20085\
        );

    \I__4635\ : InMux
    port map (
            O => \N__20116\,
            I => \N__20085\
        );

    \I__4634\ : InMux
    port map (
            O => \N__20115\,
            I => \N__20082\
        );

    \I__4633\ : InMux
    port map (
            O => \N__20114\,
            I => \N__20077\
        );

    \I__4632\ : InMux
    port map (
            O => \N__20113\,
            I => \N__20077\
        );

    \I__4631\ : Span4Mux_h
    port map (
            O => \N__20110\,
            I => \N__20072\
        );

    \I__4630\ : Span4Mux_v
    port map (
            O => \N__20107\,
            I => \N__20072\
        );

    \I__4629\ : InMux
    port map (
            O => \N__20106\,
            I => \N__20069\
        );

    \I__4628\ : Span4Mux_h
    port map (
            O => \N__20103\,
            I => \N__20064\
        );

    \I__4627\ : LocalMux
    port map (
            O => \N__20098\,
            I => \N__20064\
        );

    \I__4626\ : InMux
    port map (
            O => \N__20097\,
            I => \N__20059\
        );

    \I__4625\ : InMux
    port map (
            O => \N__20096\,
            I => \N__20059\
        );

    \I__4624\ : InMux
    port map (
            O => \N__20095\,
            I => \N__20054\
        );

    \I__4623\ : InMux
    port map (
            O => \N__20094\,
            I => \N__20054\
        );

    \I__4622\ : InMux
    port map (
            O => \N__20093\,
            I => \N__20051\
        );

    \I__4621\ : Span4Mux_h
    port map (
            O => \N__20090\,
            I => \N__20048\
        );

    \I__4620\ : LocalMux
    port map (
            O => \N__20085\,
            I => \b2v_inst.indiceZ0Z_2\
        );

    \I__4619\ : LocalMux
    port map (
            O => \N__20082\,
            I => \b2v_inst.indiceZ0Z_2\
        );

    \I__4618\ : LocalMux
    port map (
            O => \N__20077\,
            I => \b2v_inst.indiceZ0Z_2\
        );

    \I__4617\ : Odrv4
    port map (
            O => \N__20072\,
            I => \b2v_inst.indiceZ0Z_2\
        );

    \I__4616\ : LocalMux
    port map (
            O => \N__20069\,
            I => \b2v_inst.indiceZ0Z_2\
        );

    \I__4615\ : Odrv4
    port map (
            O => \N__20064\,
            I => \b2v_inst.indiceZ0Z_2\
        );

    \I__4614\ : LocalMux
    port map (
            O => \N__20059\,
            I => \b2v_inst.indiceZ0Z_2\
        );

    \I__4613\ : LocalMux
    port map (
            O => \N__20054\,
            I => \b2v_inst.indiceZ0Z_2\
        );

    \I__4612\ : LocalMux
    port map (
            O => \N__20051\,
            I => \b2v_inst.indiceZ0Z_2\
        );

    \I__4611\ : Odrv4
    port map (
            O => \N__20048\,
            I => \b2v_inst.indiceZ0Z_2\
        );

    \I__4610\ : CascadeMux
    port map (
            O => \N__20027\,
            I => \N__20024\
        );

    \I__4609\ : InMux
    port map (
            O => \N__20024\,
            I => \N__20021\
        );

    \I__4608\ : LocalMux
    port map (
            O => \N__20021\,
            I => \N__20016\
        );

    \I__4607\ : InMux
    port map (
            O => \N__20020\,
            I => \N__20013\
        );

    \I__4606\ : InMux
    port map (
            O => \N__20019\,
            I => \N__20010\
        );

    \I__4605\ : Span4Mux_v
    port map (
            O => \N__20016\,
            I => \N__20007\
        );

    \I__4604\ : LocalMux
    port map (
            O => \N__20013\,
            I => \b2v_inst.un2_dir_mem_2_c2\
        );

    \I__4603\ : LocalMux
    port map (
            O => \N__20010\,
            I => \b2v_inst.un2_dir_mem_2_c2\
        );

    \I__4602\ : Odrv4
    port map (
            O => \N__20007\,
            I => \b2v_inst.un2_dir_mem_2_c2\
        );

    \I__4601\ : InMux
    port map (
            O => \N__20000\,
            I => \N__19997\
        );

    \I__4600\ : LocalMux
    port map (
            O => \N__19997\,
            I => \N__19994\
        );

    \I__4599\ : Span4Mux_v
    port map (
            O => \N__19994\,
            I => \N__19991\
        );

    \I__4598\ : Span4Mux_h
    port map (
            O => \N__19991\,
            I => \N__19988\
        );

    \I__4597\ : Odrv4
    port map (
            O => \N__19988\,
            I => \b2v_inst.dir_mem_1Z0Z_2\
        );

    \I__4596\ : InMux
    port map (
            O => \N__19985\,
            I => \N__19982\
        );

    \I__4595\ : LocalMux
    port map (
            O => \N__19982\,
            I => \b2v_inst.dir_mem_1_RNO_0Z0Z_5\
        );

    \I__4594\ : InMux
    port map (
            O => \N__19979\,
            I => \N__19976\
        );

    \I__4593\ : LocalMux
    port map (
            O => \N__19976\,
            I => \N__19973\
        );

    \I__4592\ : Span4Mux_h
    port map (
            O => \N__19973\,
            I => \N__19970\
        );

    \I__4591\ : Span4Mux_h
    port map (
            O => \N__19970\,
            I => \N__19967\
        );

    \I__4590\ : Odrv4
    port map (
            O => \N__19967\,
            I => \b2v_inst.dir_mem_1Z0Z_5\
        );

    \I__4589\ : InMux
    port map (
            O => \N__19964\,
            I => \N__19952\
        );

    \I__4588\ : InMux
    port map (
            O => \N__19963\,
            I => \N__19952\
        );

    \I__4587\ : InMux
    port map (
            O => \N__19962\,
            I => \N__19952\
        );

    \I__4586\ : InMux
    port map (
            O => \N__19961\,
            I => \N__19952\
        );

    \I__4585\ : LocalMux
    port map (
            O => \N__19952\,
            I => \b2v_inst.dir_mem_115_0\
        );

    \I__4584\ : InMux
    port map (
            O => \N__19949\,
            I => \N__19946\
        );

    \I__4583\ : LocalMux
    port map (
            O => \N__19946\,
            I => \N__19943\
        );

    \I__4582\ : Span4Mux_h
    port map (
            O => \N__19943\,
            I => \N__19940\
        );

    \I__4581\ : Span4Mux_h
    port map (
            O => \N__19940\,
            I => \N__19937\
        );

    \I__4580\ : Odrv4
    port map (
            O => \N__19937\,
            I => \b2v_inst.dir_mem_1Z0Z_1\
        );

    \I__4579\ : CEMux
    port map (
            O => \N__19934\,
            I => \N__19930\
        );

    \I__4578\ : CEMux
    port map (
            O => \N__19933\,
            I => \N__19927\
        );

    \I__4577\ : LocalMux
    port map (
            O => \N__19930\,
            I => \N__19921\
        );

    \I__4576\ : LocalMux
    port map (
            O => \N__19927\,
            I => \N__19921\
        );

    \I__4575\ : CEMux
    port map (
            O => \N__19926\,
            I => \N__19917\
        );

    \I__4574\ : Span4Mux_v
    port map (
            O => \N__19921\,
            I => \N__19914\
        );

    \I__4573\ : CEMux
    port map (
            O => \N__19920\,
            I => \N__19911\
        );

    \I__4572\ : LocalMux
    port map (
            O => \N__19917\,
            I => \N__19908\
        );

    \I__4571\ : Sp12to4
    port map (
            O => \N__19914\,
            I => \N__19905\
        );

    \I__4570\ : LocalMux
    port map (
            O => \N__19911\,
            I => \N__19900\
        );

    \I__4569\ : Span4Mux_v
    port map (
            O => \N__19908\,
            I => \N__19900\
        );

    \I__4568\ : Odrv12
    port map (
            O => \N__19905\,
            I => \b2v_inst.N_134_i\
        );

    \I__4567\ : Odrv4
    port map (
            O => \N__19900\,
            I => \b2v_inst.N_134_i\
        );

    \I__4566\ : InMux
    port map (
            O => \N__19895\,
            I => \N__19891\
        );

    \I__4565\ : InMux
    port map (
            O => \N__19894\,
            I => \N__19886\
        );

    \I__4564\ : LocalMux
    port map (
            O => \N__19891\,
            I => \N__19883\
        );

    \I__4563\ : InMux
    port map (
            O => \N__19890\,
            I => \N__19880\
        );

    \I__4562\ : CascadeMux
    port map (
            O => \N__19889\,
            I => \N__19877\
        );

    \I__4561\ : LocalMux
    port map (
            O => \N__19886\,
            I => \N__19870\
        );

    \I__4560\ : Span4Mux_h
    port map (
            O => \N__19883\,
            I => \N__19866\
        );

    \I__4559\ : LocalMux
    port map (
            O => \N__19880\,
            I => \N__19863\
        );

    \I__4558\ : InMux
    port map (
            O => \N__19877\,
            I => \N__19857\
        );

    \I__4557\ : InMux
    port map (
            O => \N__19876\,
            I => \N__19857\
        );

    \I__4556\ : InMux
    port map (
            O => \N__19875\,
            I => \N__19852\
        );

    \I__4555\ : InMux
    port map (
            O => \N__19874\,
            I => \N__19852\
        );

    \I__4554\ : InMux
    port map (
            O => \N__19873\,
            I => \N__19849\
        );

    \I__4553\ : Span4Mux_h
    port map (
            O => \N__19870\,
            I => \N__19846\
        );

    \I__4552\ : InMux
    port map (
            O => \N__19869\,
            I => \N__19843\
        );

    \I__4551\ : Span4Mux_h
    port map (
            O => \N__19866\,
            I => \N__19838\
        );

    \I__4550\ : Span4Mux_h
    port map (
            O => \N__19863\,
            I => \N__19838\
        );

    \I__4549\ : InMux
    port map (
            O => \N__19862\,
            I => \N__19835\
        );

    \I__4548\ : LocalMux
    port map (
            O => \N__19857\,
            I => \N__19830\
        );

    \I__4547\ : LocalMux
    port map (
            O => \N__19852\,
            I => \N__19830\
        );

    \I__4546\ : LocalMux
    port map (
            O => \N__19849\,
            I => \b2v_inst.dir_memZ0Z_0\
        );

    \I__4545\ : Odrv4
    port map (
            O => \N__19846\,
            I => \b2v_inst.dir_memZ0Z_0\
        );

    \I__4544\ : LocalMux
    port map (
            O => \N__19843\,
            I => \b2v_inst.dir_memZ0Z_0\
        );

    \I__4543\ : Odrv4
    port map (
            O => \N__19838\,
            I => \b2v_inst.dir_memZ0Z_0\
        );

    \I__4542\ : LocalMux
    port map (
            O => \N__19835\,
            I => \b2v_inst.dir_memZ0Z_0\
        );

    \I__4541\ : Odrv4
    port map (
            O => \N__19830\,
            I => \b2v_inst.dir_memZ0Z_0\
        );

    \I__4540\ : InMux
    port map (
            O => \N__19817\,
            I => \N__19812\
        );

    \I__4539\ : InMux
    port map (
            O => \N__19816\,
            I => \N__19809\
        );

    \I__4538\ : InMux
    port map (
            O => \N__19815\,
            I => \N__19801\
        );

    \I__4537\ : LocalMux
    port map (
            O => \N__19812\,
            I => \N__19798\
        );

    \I__4536\ : LocalMux
    port map (
            O => \N__19809\,
            I => \N__19795\
        );

    \I__4535\ : InMux
    port map (
            O => \N__19808\,
            I => \N__19792\
        );

    \I__4534\ : InMux
    port map (
            O => \N__19807\,
            I => \N__19789\
        );

    \I__4533\ : InMux
    port map (
            O => \N__19806\,
            I => \N__19786\
        );

    \I__4532\ : InMux
    port map (
            O => \N__19805\,
            I => \N__19781\
        );

    \I__4531\ : InMux
    port map (
            O => \N__19804\,
            I => \N__19781\
        );

    \I__4530\ : LocalMux
    port map (
            O => \N__19801\,
            I => \N__19778\
        );

    \I__4529\ : Span4Mux_h
    port map (
            O => \N__19798\,
            I => \N__19773\
        );

    \I__4528\ : Span4Mux_h
    port map (
            O => \N__19795\,
            I => \N__19773\
        );

    \I__4527\ : LocalMux
    port map (
            O => \N__19792\,
            I => \b2v_inst.dir_memZ0Z_1\
        );

    \I__4526\ : LocalMux
    port map (
            O => \N__19789\,
            I => \b2v_inst.dir_memZ0Z_1\
        );

    \I__4525\ : LocalMux
    port map (
            O => \N__19786\,
            I => \b2v_inst.dir_memZ0Z_1\
        );

    \I__4524\ : LocalMux
    port map (
            O => \N__19781\,
            I => \b2v_inst.dir_memZ0Z_1\
        );

    \I__4523\ : Odrv4
    port map (
            O => \N__19778\,
            I => \b2v_inst.dir_memZ0Z_1\
        );

    \I__4522\ : Odrv4
    port map (
            O => \N__19773\,
            I => \b2v_inst.dir_memZ0Z_1\
        );

    \I__4521\ : InMux
    port map (
            O => \N__19760\,
            I => \N__19751\
        );

    \I__4520\ : InMux
    port map (
            O => \N__19759\,
            I => \N__19744\
        );

    \I__4519\ : InMux
    port map (
            O => \N__19758\,
            I => \N__19744\
        );

    \I__4518\ : InMux
    port map (
            O => \N__19757\,
            I => \N__19744\
        );

    \I__4517\ : InMux
    port map (
            O => \N__19756\,
            I => \N__19741\
        );

    \I__4516\ : InMux
    port map (
            O => \N__19755\,
            I => \N__19735\
        );

    \I__4515\ : InMux
    port map (
            O => \N__19754\,
            I => \N__19735\
        );

    \I__4514\ : LocalMux
    port map (
            O => \N__19751\,
            I => \N__19728\
        );

    \I__4513\ : LocalMux
    port map (
            O => \N__19744\,
            I => \N__19728\
        );

    \I__4512\ : LocalMux
    port map (
            O => \N__19741\,
            I => \N__19728\
        );

    \I__4511\ : InMux
    port map (
            O => \N__19740\,
            I => \N__19718\
        );

    \I__4510\ : LocalMux
    port map (
            O => \N__19735\,
            I => \N__19713\
        );

    \I__4509\ : Span4Mux_v
    port map (
            O => \N__19728\,
            I => \N__19713\
        );

    \I__4508\ : InMux
    port map (
            O => \N__19727\,
            I => \N__19708\
        );

    \I__4507\ : InMux
    port map (
            O => \N__19726\,
            I => \N__19708\
        );

    \I__4506\ : InMux
    port map (
            O => \N__19725\,
            I => \N__19703\
        );

    \I__4505\ : InMux
    port map (
            O => \N__19724\,
            I => \N__19703\
        );

    \I__4504\ : InMux
    port map (
            O => \N__19723\,
            I => \N__19696\
        );

    \I__4503\ : InMux
    port map (
            O => \N__19722\,
            I => \N__19696\
        );

    \I__4502\ : InMux
    port map (
            O => \N__19721\,
            I => \N__19696\
        );

    \I__4501\ : LocalMux
    port map (
            O => \N__19718\,
            I => \b2v_inst.N_253\
        );

    \I__4500\ : Odrv4
    port map (
            O => \N__19713\,
            I => \b2v_inst.N_253\
        );

    \I__4499\ : LocalMux
    port map (
            O => \N__19708\,
            I => \b2v_inst.N_253\
        );

    \I__4498\ : LocalMux
    port map (
            O => \N__19703\,
            I => \b2v_inst.N_253\
        );

    \I__4497\ : LocalMux
    port map (
            O => \N__19696\,
            I => \b2v_inst.N_253\
        );

    \I__4496\ : CascadeMux
    port map (
            O => \N__19685\,
            I => \N__19682\
        );

    \I__4495\ : InMux
    port map (
            O => \N__19682\,
            I => \N__19679\
        );

    \I__4494\ : LocalMux
    port map (
            O => \N__19679\,
            I => \N__19676\
        );

    \I__4493\ : Odrv4
    port map (
            O => \N__19676\,
            I => \b2v_inst.un2_indice_21_s1_1\
        );

    \I__4492\ : InMux
    port map (
            O => \N__19673\,
            I => \N__19668\
        );

    \I__4491\ : InMux
    port map (
            O => \N__19672\,
            I => \N__19660\
        );

    \I__4490\ : InMux
    port map (
            O => \N__19671\,
            I => \N__19660\
        );

    \I__4489\ : LocalMux
    port map (
            O => \N__19668\,
            I => \N__19657\
        );

    \I__4488\ : InMux
    port map (
            O => \N__19667\,
            I => \N__19652\
        );

    \I__4487\ : InMux
    port map (
            O => \N__19666\,
            I => \N__19649\
        );

    \I__4486\ : InMux
    port map (
            O => \N__19665\,
            I => \N__19646\
        );

    \I__4485\ : LocalMux
    port map (
            O => \N__19660\,
            I => \N__19643\
        );

    \I__4484\ : Span4Mux_h
    port map (
            O => \N__19657\,
            I => \N__19640\
        );

    \I__4483\ : InMux
    port map (
            O => \N__19656\,
            I => \N__19637\
        );

    \I__4482\ : InMux
    port map (
            O => \N__19655\,
            I => \N__19634\
        );

    \I__4481\ : LocalMux
    port map (
            O => \N__19652\,
            I => \N__19631\
        );

    \I__4480\ : LocalMux
    port map (
            O => \N__19649\,
            I => \b2v_inst.un10_indice_2\
        );

    \I__4479\ : LocalMux
    port map (
            O => \N__19646\,
            I => \b2v_inst.un10_indice_2\
        );

    \I__4478\ : Odrv4
    port map (
            O => \N__19643\,
            I => \b2v_inst.un10_indice_2\
        );

    \I__4477\ : Odrv4
    port map (
            O => \N__19640\,
            I => \b2v_inst.un10_indice_2\
        );

    \I__4476\ : LocalMux
    port map (
            O => \N__19637\,
            I => \b2v_inst.un10_indice_2\
        );

    \I__4475\ : LocalMux
    port map (
            O => \N__19634\,
            I => \b2v_inst.un10_indice_2\
        );

    \I__4474\ : Odrv4
    port map (
            O => \N__19631\,
            I => \b2v_inst.un10_indice_2\
        );

    \I__4473\ : CascadeMux
    port map (
            O => \N__19616\,
            I => \N__19610\
        );

    \I__4472\ : InMux
    port map (
            O => \N__19615\,
            I => \N__19607\
        );

    \I__4471\ : CascadeMux
    port map (
            O => \N__19614\,
            I => \N__19604\
        );

    \I__4470\ : InMux
    port map (
            O => \N__19613\,
            I => \N__19598\
        );

    \I__4469\ : InMux
    port map (
            O => \N__19610\,
            I => \N__19598\
        );

    \I__4468\ : LocalMux
    port map (
            O => \N__19607\,
            I => \N__19595\
        );

    \I__4467\ : InMux
    port map (
            O => \N__19604\,
            I => \N__19592\
        );

    \I__4466\ : InMux
    port map (
            O => \N__19603\,
            I => \N__19589\
        );

    \I__4465\ : LocalMux
    port map (
            O => \N__19598\,
            I => \N__19584\
        );

    \I__4464\ : Span4Mux_h
    port map (
            O => \N__19595\,
            I => \N__19581\
        );

    \I__4463\ : LocalMux
    port map (
            O => \N__19592\,
            I => \N__19576\
        );

    \I__4462\ : LocalMux
    port map (
            O => \N__19589\,
            I => \N__19576\
        );

    \I__4461\ : InMux
    port map (
            O => \N__19588\,
            I => \N__19573\
        );

    \I__4460\ : InMux
    port map (
            O => \N__19587\,
            I => \N__19570\
        );

    \I__4459\ : Span4Mux_v
    port map (
            O => \N__19584\,
            I => \N__19563\
        );

    \I__4458\ : Span4Mux_v
    port map (
            O => \N__19581\,
            I => \N__19563\
        );

    \I__4457\ : Span4Mux_v
    port map (
            O => \N__19576\,
            I => \N__19563\
        );

    \I__4456\ : LocalMux
    port map (
            O => \N__19573\,
            I => \b2v_inst.CO1\
        );

    \I__4455\ : LocalMux
    port map (
            O => \N__19570\,
            I => \b2v_inst.CO1\
        );

    \I__4454\ : Odrv4
    port map (
            O => \N__19563\,
            I => \b2v_inst.CO1\
        );

    \I__4453\ : CascadeMux
    port map (
            O => \N__19556\,
            I => \b2v_inst.CO1_cascade_\
        );

    \I__4452\ : CascadeMux
    port map (
            O => \N__19553\,
            I => \b2v_inst.un2_dir_mem_2_c2_cascade_\
        );

    \I__4451\ : InMux
    port map (
            O => \N__19550\,
            I => \N__19541\
        );

    \I__4450\ : InMux
    port map (
            O => \N__19549\,
            I => \N__19541\
        );

    \I__4449\ : InMux
    port map (
            O => \N__19548\,
            I => \N__19541\
        );

    \I__4448\ : LocalMux
    port map (
            O => \N__19541\,
            I => \b2v_inst.indice_fastZ0Z_0\
        );

    \I__4447\ : CascadeMux
    port map (
            O => \N__19538\,
            I => \N__19533\
        );

    \I__4446\ : CascadeMux
    port map (
            O => \N__19537\,
            I => \N__19530\
        );

    \I__4445\ : InMux
    port map (
            O => \N__19536\,
            I => \N__19523\
        );

    \I__4444\ : InMux
    port map (
            O => \N__19533\,
            I => \N__19523\
        );

    \I__4443\ : InMux
    port map (
            O => \N__19530\,
            I => \N__19523\
        );

    \I__4442\ : LocalMux
    port map (
            O => \N__19523\,
            I => \b2v_inst.indice_fastZ0Z_1\
        );

    \I__4441\ : CascadeMux
    port map (
            O => \N__19520\,
            I => \N__19511\
        );

    \I__4440\ : CascadeMux
    port map (
            O => \N__19519\,
            I => \N__19508\
        );

    \I__4439\ : CascadeMux
    port map (
            O => \N__19518\,
            I => \N__19505\
        );

    \I__4438\ : CascadeMux
    port map (
            O => \N__19517\,
            I => \N__19501\
        );

    \I__4437\ : CascadeMux
    port map (
            O => \N__19516\,
            I => \N__19498\
        );

    \I__4436\ : CascadeMux
    port map (
            O => \N__19515\,
            I => \N__19495\
        );

    \I__4435\ : InMux
    port map (
            O => \N__19514\,
            I => \N__19492\
        );

    \I__4434\ : InMux
    port map (
            O => \N__19511\,
            I => \N__19489\
        );

    \I__4433\ : InMux
    port map (
            O => \N__19508\,
            I => \N__19486\
        );

    \I__4432\ : InMux
    port map (
            O => \N__19505\,
            I => \N__19483\
        );

    \I__4431\ : InMux
    port map (
            O => \N__19504\,
            I => \N__19478\
        );

    \I__4430\ : InMux
    port map (
            O => \N__19501\,
            I => \N__19478\
        );

    \I__4429\ : InMux
    port map (
            O => \N__19498\,
            I => \N__19473\
        );

    \I__4428\ : InMux
    port map (
            O => \N__19495\,
            I => \N__19473\
        );

    \I__4427\ : LocalMux
    port map (
            O => \N__19492\,
            I => \N__19469\
        );

    \I__4426\ : LocalMux
    port map (
            O => \N__19489\,
            I => \N__19463\
        );

    \I__4425\ : LocalMux
    port map (
            O => \N__19486\,
            I => \N__19460\
        );

    \I__4424\ : LocalMux
    port map (
            O => \N__19483\,
            I => \N__19455\
        );

    \I__4423\ : LocalMux
    port map (
            O => \N__19478\,
            I => \N__19455\
        );

    \I__4422\ : LocalMux
    port map (
            O => \N__19473\,
            I => \N__19452\
        );

    \I__4421\ : InMux
    port map (
            O => \N__19472\,
            I => \N__19449\
        );

    \I__4420\ : Span4Mux_h
    port map (
            O => \N__19469\,
            I => \N__19446\
        );

    \I__4419\ : InMux
    port map (
            O => \N__19468\,
            I => \N__19439\
        );

    \I__4418\ : InMux
    port map (
            O => \N__19467\,
            I => \N__19439\
        );

    \I__4417\ : InMux
    port map (
            O => \N__19466\,
            I => \N__19439\
        );

    \I__4416\ : Span4Mux_v
    port map (
            O => \N__19463\,
            I => \N__19432\
        );

    \I__4415\ : Span4Mux_v
    port map (
            O => \N__19460\,
            I => \N__19432\
        );

    \I__4414\ : Span4Mux_h
    port map (
            O => \N__19455\,
            I => \N__19432\
        );

    \I__4413\ : Span4Mux_h
    port map (
            O => \N__19452\,
            I => \N__19429\
        );

    \I__4412\ : LocalMux
    port map (
            O => \N__19449\,
            I => \b2v_inst.indice_2_repZ0Z1\
        );

    \I__4411\ : Odrv4
    port map (
            O => \N__19446\,
            I => \b2v_inst.indice_2_repZ0Z1\
        );

    \I__4410\ : LocalMux
    port map (
            O => \N__19439\,
            I => \b2v_inst.indice_2_repZ0Z1\
        );

    \I__4409\ : Odrv4
    port map (
            O => \N__19432\,
            I => \b2v_inst.indice_2_repZ0Z1\
        );

    \I__4408\ : Odrv4
    port map (
            O => \N__19429\,
            I => \b2v_inst.indice_2_repZ0Z1\
        );

    \I__4407\ : InMux
    port map (
            O => \N__19418\,
            I => \N__19412\
        );

    \I__4406\ : InMux
    port map (
            O => \N__19417\,
            I => \N__19408\
        );

    \I__4405\ : InMux
    port map (
            O => \N__19416\,
            I => \N__19405\
        );

    \I__4404\ : InMux
    port map (
            O => \N__19415\,
            I => \N__19402\
        );

    \I__4403\ : LocalMux
    port map (
            O => \N__19412\,
            I => \N__19399\
        );

    \I__4402\ : InMux
    port map (
            O => \N__19411\,
            I => \N__19396\
        );

    \I__4401\ : LocalMux
    port map (
            O => \N__19408\,
            I => \b2v_inst1.m6_2\
        );

    \I__4400\ : LocalMux
    port map (
            O => \N__19405\,
            I => \b2v_inst1.m6_2\
        );

    \I__4399\ : LocalMux
    port map (
            O => \N__19402\,
            I => \b2v_inst1.m6_2\
        );

    \I__4398\ : Odrv4
    port map (
            O => \N__19399\,
            I => \b2v_inst1.m6_2\
        );

    \I__4397\ : LocalMux
    port map (
            O => \N__19396\,
            I => \b2v_inst1.m6_2\
        );

    \I__4396\ : CascadeMux
    port map (
            O => \N__19385\,
            I => \N__19382\
        );

    \I__4395\ : InMux
    port map (
            O => \N__19382\,
            I => \N__19379\
        );

    \I__4394\ : LocalMux
    port map (
            O => \N__19379\,
            I => \N__19376\
        );

    \I__4393\ : Odrv4
    port map (
            O => \N__19376\,
            I => \b2v_inst.un2_indice_0_d1_c5\
        );

    \I__4392\ : InMux
    port map (
            O => \N__19373\,
            I => \N__19369\
        );

    \I__4391\ : InMux
    port map (
            O => \N__19372\,
            I => \N__19366\
        );

    \I__4390\ : LocalMux
    port map (
            O => \N__19369\,
            I => \N__19363\
        );

    \I__4389\ : LocalMux
    port map (
            O => \N__19366\,
            I => \N__19358\
        );

    \I__4388\ : Span4Mux_v
    port map (
            O => \N__19363\,
            I => \N__19354\
        );

    \I__4387\ : InMux
    port map (
            O => \N__19362\,
            I => \N__19351\
        );

    \I__4386\ : InMux
    port map (
            O => \N__19361\,
            I => \N__19348\
        );

    \I__4385\ : Span4Mux_h
    port map (
            O => \N__19358\,
            I => \N__19345\
        );

    \I__4384\ : InMux
    port map (
            O => \N__19357\,
            I => \N__19342\
        );

    \I__4383\ : Odrv4
    port map (
            O => \N__19354\,
            I => \b2v_inst.dir_memZ0Z_4\
        );

    \I__4382\ : LocalMux
    port map (
            O => \N__19351\,
            I => \b2v_inst.dir_memZ0Z_4\
        );

    \I__4381\ : LocalMux
    port map (
            O => \N__19348\,
            I => \b2v_inst.dir_memZ0Z_4\
        );

    \I__4380\ : Odrv4
    port map (
            O => \N__19345\,
            I => \b2v_inst.dir_memZ0Z_4\
        );

    \I__4379\ : LocalMux
    port map (
            O => \N__19342\,
            I => \b2v_inst.dir_memZ0Z_4\
        );

    \I__4378\ : CascadeMux
    port map (
            O => \N__19331\,
            I => \N__19328\
        );

    \I__4377\ : InMux
    port map (
            O => \N__19328\,
            I => \N__19325\
        );

    \I__4376\ : LocalMux
    port map (
            O => \N__19325\,
            I => \b2v_inst.un2_indice_0_d1_ac0_7_s_0_0\
        );

    \I__4375\ : InMux
    port map (
            O => \N__19322\,
            I => \N__19316\
        );

    \I__4374\ : CascadeMux
    port map (
            O => \N__19321\,
            I => \N__19312\
        );

    \I__4373\ : InMux
    port map (
            O => \N__19320\,
            I => \N__19309\
        );

    \I__4372\ : InMux
    port map (
            O => \N__19319\,
            I => \N__19306\
        );

    \I__4371\ : LocalMux
    port map (
            O => \N__19316\,
            I => \N__19303\
        );

    \I__4370\ : InMux
    port map (
            O => \N__19315\,
            I => \N__19296\
        );

    \I__4369\ : InMux
    port map (
            O => \N__19312\,
            I => \N__19296\
        );

    \I__4368\ : LocalMux
    port map (
            O => \N__19309\,
            I => \N__19293\
        );

    \I__4367\ : LocalMux
    port map (
            O => \N__19306\,
            I => \N__19290\
        );

    \I__4366\ : Span4Mux_v
    port map (
            O => \N__19303\,
            I => \N__19287\
        );

    \I__4365\ : InMux
    port map (
            O => \N__19302\,
            I => \N__19282\
        );

    \I__4364\ : InMux
    port map (
            O => \N__19301\,
            I => \N__19282\
        );

    \I__4363\ : LocalMux
    port map (
            O => \N__19296\,
            I => \N__19277\
        );

    \I__4362\ : Span4Mux_v
    port map (
            O => \N__19293\,
            I => \N__19277\
        );

    \I__4361\ : Span4Mux_h
    port map (
            O => \N__19290\,
            I => \N__19274\
        );

    \I__4360\ : Odrv4
    port map (
            O => \N__19287\,
            I => \b2v_inst.dir_memZ0Z_3\
        );

    \I__4359\ : LocalMux
    port map (
            O => \N__19282\,
            I => \b2v_inst.dir_memZ0Z_3\
        );

    \I__4358\ : Odrv4
    port map (
            O => \N__19277\,
            I => \b2v_inst.dir_memZ0Z_3\
        );

    \I__4357\ : Odrv4
    port map (
            O => \N__19274\,
            I => \b2v_inst.dir_memZ0Z_3\
        );

    \I__4356\ : InMux
    port map (
            O => \N__19265\,
            I => \N__19261\
        );

    \I__4355\ : InMux
    port map (
            O => \N__19264\,
            I => \N__19257\
        );

    \I__4354\ : LocalMux
    port map (
            O => \N__19261\,
            I => \N__19252\
        );

    \I__4353\ : CascadeMux
    port map (
            O => \N__19260\,
            I => \N__19249\
        );

    \I__4352\ : LocalMux
    port map (
            O => \N__19257\,
            I => \N__19246\
        );

    \I__4351\ : InMux
    port map (
            O => \N__19256\,
            I => \N__19243\
        );

    \I__4350\ : InMux
    port map (
            O => \N__19255\,
            I => \N__19240\
        );

    \I__4349\ : Span4Mux_v
    port map (
            O => \N__19252\,
            I => \N__19237\
        );

    \I__4348\ : InMux
    port map (
            O => \N__19249\,
            I => \N__19234\
        );

    \I__4347\ : Span4Mux_h
    port map (
            O => \N__19246\,
            I => \N__19229\
        );

    \I__4346\ : LocalMux
    port map (
            O => \N__19243\,
            I => \N__19229\
        );

    \I__4345\ : LocalMux
    port map (
            O => \N__19240\,
            I => \b2v_inst.dir_memZ0Z_5\
        );

    \I__4344\ : Odrv4
    port map (
            O => \N__19237\,
            I => \b2v_inst.dir_memZ0Z_5\
        );

    \I__4343\ : LocalMux
    port map (
            O => \N__19234\,
            I => \b2v_inst.dir_memZ0Z_5\
        );

    \I__4342\ : Odrv4
    port map (
            O => \N__19229\,
            I => \b2v_inst.dir_memZ0Z_5\
        );

    \I__4341\ : CascadeMux
    port map (
            O => \N__19220\,
            I => \b2v_inst.un2_indice_0_d1_ac0_7_s_0_0_cascade_\
        );

    \I__4340\ : InMux
    port map (
            O => \N__19217\,
            I => \N__19214\
        );

    \I__4339\ : LocalMux
    port map (
            O => \N__19214\,
            I => \N__19209\
        );

    \I__4338\ : InMux
    port map (
            O => \N__19213\,
            I => \N__19206\
        );

    \I__4337\ : CascadeMux
    port map (
            O => \N__19212\,
            I => \N__19202\
        );

    \I__4336\ : Span4Mux_h
    port map (
            O => \N__19209\,
            I => \N__19195\
        );

    \I__4335\ : LocalMux
    port map (
            O => \N__19206\,
            I => \N__19192\
        );

    \I__4334\ : InMux
    port map (
            O => \N__19205\,
            I => \N__19189\
        );

    \I__4333\ : InMux
    port map (
            O => \N__19202\,
            I => \N__19186\
        );

    \I__4332\ : InMux
    port map (
            O => \N__19201\,
            I => \N__19181\
        );

    \I__4331\ : InMux
    port map (
            O => \N__19200\,
            I => \N__19181\
        );

    \I__4330\ : InMux
    port map (
            O => \N__19199\,
            I => \N__19176\
        );

    \I__4329\ : InMux
    port map (
            O => \N__19198\,
            I => \N__19176\
        );

    \I__4328\ : Span4Mux_v
    port map (
            O => \N__19195\,
            I => \N__19169\
        );

    \I__4327\ : Span4Mux_v
    port map (
            O => \N__19192\,
            I => \N__19169\
        );

    \I__4326\ : LocalMux
    port map (
            O => \N__19189\,
            I => \N__19169\
        );

    \I__4325\ : LocalMux
    port map (
            O => \N__19186\,
            I => \b2v_inst.dir_memZ0Z_2\
        );

    \I__4324\ : LocalMux
    port map (
            O => \N__19181\,
            I => \b2v_inst.dir_memZ0Z_2\
        );

    \I__4323\ : LocalMux
    port map (
            O => \N__19176\,
            I => \b2v_inst.dir_memZ0Z_2\
        );

    \I__4322\ : Odrv4
    port map (
            O => \N__19169\,
            I => \b2v_inst.dir_memZ0Z_2\
        );

    \I__4321\ : InMux
    port map (
            O => \N__19160\,
            I => \N__19156\
        );

    \I__4320\ : CascadeMux
    port map (
            O => \N__19159\,
            I => \N__19153\
        );

    \I__4319\ : LocalMux
    port map (
            O => \N__19156\,
            I => \N__19150\
        );

    \I__4318\ : InMux
    port map (
            O => \N__19153\,
            I => \N__19146\
        );

    \I__4317\ : Span4Mux_v
    port map (
            O => \N__19150\,
            I => \N__19143\
        );

    \I__4316\ : InMux
    port map (
            O => \N__19149\,
            I => \N__19140\
        );

    \I__4315\ : LocalMux
    port map (
            O => \N__19146\,
            I => \N__19137\
        );

    \I__4314\ : Odrv4
    port map (
            O => \N__19143\,
            I => \b2v_inst.dir_memZ0Z_7\
        );

    \I__4313\ : LocalMux
    port map (
            O => \N__19140\,
            I => \b2v_inst.dir_memZ0Z_7\
        );

    \I__4312\ : Odrv4
    port map (
            O => \N__19137\,
            I => \b2v_inst.dir_memZ0Z_7\
        );

    \I__4311\ : CascadeMux
    port map (
            O => \N__19130\,
            I => \b2v_inst.un2_indice_0_d1_ac0_9_0_cascade_\
        );

    \I__4310\ : InMux
    port map (
            O => \N__19127\,
            I => \N__19123\
        );

    \I__4309\ : InMux
    port map (
            O => \N__19126\,
            I => \N__19120\
        );

    \I__4308\ : LocalMux
    port map (
            O => \N__19123\,
            I => \N__19116\
        );

    \I__4307\ : LocalMux
    port map (
            O => \N__19120\,
            I => \N__19113\
        );

    \I__4306\ : CascadeMux
    port map (
            O => \N__19119\,
            I => \N__19109\
        );

    \I__4305\ : Span4Mux_v
    port map (
            O => \N__19116\,
            I => \N__19106\
        );

    \I__4304\ : Span4Mux_h
    port map (
            O => \N__19113\,
            I => \N__19103\
        );

    \I__4303\ : InMux
    port map (
            O => \N__19112\,
            I => \N__19098\
        );

    \I__4302\ : InMux
    port map (
            O => \N__19109\,
            I => \N__19098\
        );

    \I__4301\ : Odrv4
    port map (
            O => \N__19106\,
            I => \b2v_inst.dir_memZ0Z_6\
        );

    \I__4300\ : Odrv4
    port map (
            O => \N__19103\,
            I => \b2v_inst.dir_memZ0Z_6\
        );

    \I__4299\ : LocalMux
    port map (
            O => \N__19098\,
            I => \b2v_inst.dir_memZ0Z_6\
        );

    \I__4298\ : InMux
    port map (
            O => \N__19091\,
            I => \N__19088\
        );

    \I__4297\ : LocalMux
    port map (
            O => \N__19088\,
            I => \N__19085\
        );

    \I__4296\ : Odrv4
    port map (
            O => \N__19085\,
            I => \b2v_inst.un2_indice_21_s1_7\
        );

    \I__4295\ : InMux
    port map (
            O => \N__19082\,
            I => \N__19077\
        );

    \I__4294\ : InMux
    port map (
            O => \N__19081\,
            I => \N__19072\
        );

    \I__4293\ : InMux
    port map (
            O => \N__19080\,
            I => \N__19067\
        );

    \I__4292\ : LocalMux
    port map (
            O => \N__19077\,
            I => \N__19063\
        );

    \I__4291\ : InMux
    port map (
            O => \N__19076\,
            I => \N__19059\
        );

    \I__4290\ : InMux
    port map (
            O => \N__19075\,
            I => \N__19056\
        );

    \I__4289\ : LocalMux
    port map (
            O => \N__19072\,
            I => \N__19053\
        );

    \I__4288\ : InMux
    port map (
            O => \N__19071\,
            I => \N__19049\
        );

    \I__4287\ : InMux
    port map (
            O => \N__19070\,
            I => \N__19045\
        );

    \I__4286\ : LocalMux
    port map (
            O => \N__19067\,
            I => \N__19042\
        );

    \I__4285\ : InMux
    port map (
            O => \N__19066\,
            I => \N__19039\
        );

    \I__4284\ : Span4Mux_h
    port map (
            O => \N__19063\,
            I => \N__19036\
        );

    \I__4283\ : InMux
    port map (
            O => \N__19062\,
            I => \N__19033\
        );

    \I__4282\ : LocalMux
    port map (
            O => \N__19059\,
            I => \N__19026\
        );

    \I__4281\ : LocalMux
    port map (
            O => \N__19056\,
            I => \N__19026\
        );

    \I__4280\ : Span4Mux_v
    port map (
            O => \N__19053\,
            I => \N__19026\
        );

    \I__4279\ : InMux
    port map (
            O => \N__19052\,
            I => \N__19023\
        );

    \I__4278\ : LocalMux
    port map (
            O => \N__19049\,
            I => \N__19020\
        );

    \I__4277\ : InMux
    port map (
            O => \N__19048\,
            I => \N__19017\
        );

    \I__4276\ : LocalMux
    port map (
            O => \N__19045\,
            I => \b2v_inst.state_17_repZ0Z1\
        );

    \I__4275\ : Odrv4
    port map (
            O => \N__19042\,
            I => \b2v_inst.state_17_repZ0Z1\
        );

    \I__4274\ : LocalMux
    port map (
            O => \N__19039\,
            I => \b2v_inst.state_17_repZ0Z1\
        );

    \I__4273\ : Odrv4
    port map (
            O => \N__19036\,
            I => \b2v_inst.state_17_repZ0Z1\
        );

    \I__4272\ : LocalMux
    port map (
            O => \N__19033\,
            I => \b2v_inst.state_17_repZ0Z1\
        );

    \I__4271\ : Odrv4
    port map (
            O => \N__19026\,
            I => \b2v_inst.state_17_repZ0Z1\
        );

    \I__4270\ : LocalMux
    port map (
            O => \N__19023\,
            I => \b2v_inst.state_17_repZ0Z1\
        );

    \I__4269\ : Odrv12
    port map (
            O => \N__19020\,
            I => \b2v_inst.state_17_repZ0Z1\
        );

    \I__4268\ : LocalMux
    port map (
            O => \N__19017\,
            I => \b2v_inst.state_17_repZ0Z1\
        );

    \I__4267\ : InMux
    port map (
            O => \N__18998\,
            I => \N__18994\
        );

    \I__4266\ : InMux
    port map (
            O => \N__18997\,
            I => \N__18991\
        );

    \I__4265\ : LocalMux
    port map (
            O => \N__18994\,
            I => \N__18987\
        );

    \I__4264\ : LocalMux
    port map (
            O => \N__18991\,
            I => \N__18978\
        );

    \I__4263\ : InMux
    port map (
            O => \N__18990\,
            I => \N__18975\
        );

    \I__4262\ : Span4Mux_v
    port map (
            O => \N__18987\,
            I => \N__18972\
        );

    \I__4261\ : InMux
    port map (
            O => \N__18986\,
            I => \N__18969\
        );

    \I__4260\ : InMux
    port map (
            O => \N__18985\,
            I => \N__18962\
        );

    \I__4259\ : InMux
    port map (
            O => \N__18984\,
            I => \N__18962\
        );

    \I__4258\ : InMux
    port map (
            O => \N__18983\,
            I => \N__18962\
        );

    \I__4257\ : InMux
    port map (
            O => \N__18982\,
            I => \N__18957\
        );

    \I__4256\ : InMux
    port map (
            O => \N__18981\,
            I => \N__18957\
        );

    \I__4255\ : Span4Mux_v
    port map (
            O => \N__18978\,
            I => \N__18952\
        );

    \I__4254\ : LocalMux
    port map (
            O => \N__18975\,
            I => \N__18952\
        );

    \I__4253\ : Odrv4
    port map (
            O => \N__18972\,
            I => \b2v_inst.stateZ0Z_15\
        );

    \I__4252\ : LocalMux
    port map (
            O => \N__18969\,
            I => \b2v_inst.stateZ0Z_15\
        );

    \I__4251\ : LocalMux
    port map (
            O => \N__18962\,
            I => \b2v_inst.stateZ0Z_15\
        );

    \I__4250\ : LocalMux
    port map (
            O => \N__18957\,
            I => \b2v_inst.stateZ0Z_15\
        );

    \I__4249\ : Odrv4
    port map (
            O => \N__18952\,
            I => \b2v_inst.stateZ0Z_15\
        );

    \I__4248\ : CascadeMux
    port map (
            O => \N__18941\,
            I => \N__18934\
        );

    \I__4247\ : CascadeMux
    port map (
            O => \N__18940\,
            I => \N__18928\
        );

    \I__4246\ : CascadeMux
    port map (
            O => \N__18939\,
            I => \N__18924\
        );

    \I__4245\ : InMux
    port map (
            O => \N__18938\,
            I => \N__18919\
        );

    \I__4244\ : InMux
    port map (
            O => \N__18937\,
            I => \N__18911\
        );

    \I__4243\ : InMux
    port map (
            O => \N__18934\,
            I => \N__18908\
        );

    \I__4242\ : InMux
    port map (
            O => \N__18933\,
            I => \N__18905\
        );

    \I__4241\ : InMux
    port map (
            O => \N__18932\,
            I => \N__18900\
        );

    \I__4240\ : InMux
    port map (
            O => \N__18931\,
            I => \N__18900\
        );

    \I__4239\ : InMux
    port map (
            O => \N__18928\,
            I => \N__18897\
        );

    \I__4238\ : InMux
    port map (
            O => \N__18927\,
            I => \N__18892\
        );

    \I__4237\ : InMux
    port map (
            O => \N__18924\,
            I => \N__18892\
        );

    \I__4236\ : InMux
    port map (
            O => \N__18923\,
            I => \N__18887\
        );

    \I__4235\ : InMux
    port map (
            O => \N__18922\,
            I => \N__18887\
        );

    \I__4234\ : LocalMux
    port map (
            O => \N__18919\,
            I => \N__18884\
        );

    \I__4233\ : InMux
    port map (
            O => \N__18918\,
            I => \N__18881\
        );

    \I__4232\ : InMux
    port map (
            O => \N__18917\,
            I => \N__18876\
        );

    \I__4231\ : InMux
    port map (
            O => \N__18916\,
            I => \N__18876\
        );

    \I__4230\ : InMux
    port map (
            O => \N__18915\,
            I => \N__18873\
        );

    \I__4229\ : InMux
    port map (
            O => \N__18914\,
            I => \N__18870\
        );

    \I__4228\ : LocalMux
    port map (
            O => \N__18911\,
            I => \N__18867\
        );

    \I__4227\ : LocalMux
    port map (
            O => \N__18908\,
            I => \N__18864\
        );

    \I__4226\ : LocalMux
    port map (
            O => \N__18905\,
            I => \N__18860\
        );

    \I__4225\ : LocalMux
    port map (
            O => \N__18900\,
            I => \N__18857\
        );

    \I__4224\ : LocalMux
    port map (
            O => \N__18897\,
            I => \N__18854\
        );

    \I__4223\ : LocalMux
    port map (
            O => \N__18892\,
            I => \N__18849\
        );

    \I__4222\ : LocalMux
    port map (
            O => \N__18887\,
            I => \N__18849\
        );

    \I__4221\ : Span4Mux_v
    port map (
            O => \N__18884\,
            I => \N__18842\
        );

    \I__4220\ : LocalMux
    port map (
            O => \N__18881\,
            I => \N__18842\
        );

    \I__4219\ : LocalMux
    port map (
            O => \N__18876\,
            I => \N__18842\
        );

    \I__4218\ : LocalMux
    port map (
            O => \N__18873\,
            I => \N__18836\
        );

    \I__4217\ : LocalMux
    port map (
            O => \N__18870\,
            I => \N__18836\
        );

    \I__4216\ : Span4Mux_h
    port map (
            O => \N__18867\,
            I => \N__18831\
        );

    \I__4215\ : Span4Mux_v
    port map (
            O => \N__18864\,
            I => \N__18831\
        );

    \I__4214\ : InMux
    port map (
            O => \N__18863\,
            I => \N__18828\
        );

    \I__4213\ : Span4Mux_h
    port map (
            O => \N__18860\,
            I => \N__18825\
        );

    \I__4212\ : Span4Mux_v
    port map (
            O => \N__18857\,
            I => \N__18822\
        );

    \I__4211\ : Span4Mux_v
    port map (
            O => \N__18854\,
            I => \N__18817\
        );

    \I__4210\ : Span4Mux_v
    port map (
            O => \N__18849\,
            I => \N__18817\
        );

    \I__4209\ : Span4Mux_v
    port map (
            O => \N__18842\,
            I => \N__18814\
        );

    \I__4208\ : InMux
    port map (
            O => \N__18841\,
            I => \N__18811\
        );

    \I__4207\ : Span4Mux_v
    port map (
            O => \N__18836\,
            I => \N__18808\
        );

    \I__4206\ : Span4Mux_v
    port map (
            O => \N__18831\,
            I => \N__18803\
        );

    \I__4205\ : LocalMux
    port map (
            O => \N__18828\,
            I => \N__18803\
        );

    \I__4204\ : Sp12to4
    port map (
            O => \N__18825\,
            I => \N__18800\
        );

    \I__4203\ : Sp12to4
    port map (
            O => \N__18822\,
            I => \N__18787\
        );

    \I__4202\ : Sp12to4
    port map (
            O => \N__18817\,
            I => \N__18787\
        );

    \I__4201\ : Sp12to4
    port map (
            O => \N__18814\,
            I => \N__18787\
        );

    \I__4200\ : LocalMux
    port map (
            O => \N__18811\,
            I => \N__18787\
        );

    \I__4199\ : Sp12to4
    port map (
            O => \N__18808\,
            I => \N__18787\
        );

    \I__4198\ : Sp12to4
    port map (
            O => \N__18803\,
            I => \N__18787\
        );

    \I__4197\ : Span12Mux_v
    port map (
            O => \N__18800\,
            I => \N__18782\
        );

    \I__4196\ : Span12Mux_h
    port map (
            O => \N__18787\,
            I => \N__18782\
        );

    \I__4195\ : Span12Mux_v
    port map (
            O => \N__18782\,
            I => \N__18779\
        );

    \I__4194\ : Odrv12
    port map (
            O => \N__18779\,
            I => reset
        );

    \I__4193\ : InMux
    port map (
            O => \N__18776\,
            I => \N__18759\
        );

    \I__4192\ : InMux
    port map (
            O => \N__18775\,
            I => \N__18756\
        );

    \I__4191\ : InMux
    port map (
            O => \N__18774\,
            I => \N__18753\
        );

    \I__4190\ : InMux
    port map (
            O => \N__18773\,
            I => \N__18750\
        );

    \I__4189\ : InMux
    port map (
            O => \N__18772\,
            I => \N__18746\
        );

    \I__4188\ : InMux
    port map (
            O => \N__18771\,
            I => \N__18742\
        );

    \I__4187\ : InMux
    port map (
            O => \N__18770\,
            I => \N__18735\
        );

    \I__4186\ : InMux
    port map (
            O => \N__18769\,
            I => \N__18735\
        );

    \I__4185\ : InMux
    port map (
            O => \N__18768\,
            I => \N__18735\
        );

    \I__4184\ : InMux
    port map (
            O => \N__18767\,
            I => \N__18730\
        );

    \I__4183\ : InMux
    port map (
            O => \N__18766\,
            I => \N__18730\
        );

    \I__4182\ : InMux
    port map (
            O => \N__18765\,
            I => \N__18727\
        );

    \I__4181\ : InMux
    port map (
            O => \N__18764\,
            I => \N__18724\
        );

    \I__4180\ : InMux
    port map (
            O => \N__18763\,
            I => \N__18719\
        );

    \I__4179\ : InMux
    port map (
            O => \N__18762\,
            I => \N__18719\
        );

    \I__4178\ : LocalMux
    port map (
            O => \N__18759\,
            I => \N__18716\
        );

    \I__4177\ : LocalMux
    port map (
            O => \N__18756\,
            I => \N__18713\
        );

    \I__4176\ : LocalMux
    port map (
            O => \N__18753\,
            I => \N__18710\
        );

    \I__4175\ : LocalMux
    port map (
            O => \N__18750\,
            I => \N__18704\
        );

    \I__4174\ : InMux
    port map (
            O => \N__18749\,
            I => \N__18700\
        );

    \I__4173\ : LocalMux
    port map (
            O => \N__18746\,
            I => \N__18696\
        );

    \I__4172\ : InMux
    port map (
            O => \N__18745\,
            I => \N__18693\
        );

    \I__4171\ : LocalMux
    port map (
            O => \N__18742\,
            I => \N__18686\
        );

    \I__4170\ : LocalMux
    port map (
            O => \N__18735\,
            I => \N__18686\
        );

    \I__4169\ : LocalMux
    port map (
            O => \N__18730\,
            I => \N__18686\
        );

    \I__4168\ : LocalMux
    port map (
            O => \N__18727\,
            I => \N__18683\
        );

    \I__4167\ : LocalMux
    port map (
            O => \N__18724\,
            I => \N__18678\
        );

    \I__4166\ : LocalMux
    port map (
            O => \N__18719\,
            I => \N__18678\
        );

    \I__4165\ : Span4Mux_h
    port map (
            O => \N__18716\,
            I => \N__18675\
        );

    \I__4164\ : Span4Mux_v
    port map (
            O => \N__18713\,
            I => \N__18670\
        );

    \I__4163\ : Span4Mux_v
    port map (
            O => \N__18710\,
            I => \N__18670\
        );

    \I__4162\ : InMux
    port map (
            O => \N__18709\,
            I => \N__18667\
        );

    \I__4161\ : InMux
    port map (
            O => \N__18708\,
            I => \N__18662\
        );

    \I__4160\ : InMux
    port map (
            O => \N__18707\,
            I => \N__18662\
        );

    \I__4159\ : Span4Mux_h
    port map (
            O => \N__18704\,
            I => \N__18659\
        );

    \I__4158\ : InMux
    port map (
            O => \N__18703\,
            I => \N__18656\
        );

    \I__4157\ : LocalMux
    port map (
            O => \N__18700\,
            I => \N__18653\
        );

    \I__4156\ : InMux
    port map (
            O => \N__18699\,
            I => \N__18650\
        );

    \I__4155\ : Span4Mux_h
    port map (
            O => \N__18696\,
            I => \N__18639\
        );

    \I__4154\ : LocalMux
    port map (
            O => \N__18693\,
            I => \N__18639\
        );

    \I__4153\ : Span4Mux_v
    port map (
            O => \N__18686\,
            I => \N__18639\
        );

    \I__4152\ : Span4Mux_h
    port map (
            O => \N__18683\,
            I => \N__18639\
        );

    \I__4151\ : Span4Mux_v
    port map (
            O => \N__18678\,
            I => \N__18639\
        );

    \I__4150\ : Odrv4
    port map (
            O => \N__18675\,
            I => \b2v_inst.N_351_0\
        );

    \I__4149\ : Odrv4
    port map (
            O => \N__18670\,
            I => \b2v_inst.N_351_0\
        );

    \I__4148\ : LocalMux
    port map (
            O => \N__18667\,
            I => \b2v_inst.N_351_0\
        );

    \I__4147\ : LocalMux
    port map (
            O => \N__18662\,
            I => \b2v_inst.N_351_0\
        );

    \I__4146\ : Odrv4
    port map (
            O => \N__18659\,
            I => \b2v_inst.N_351_0\
        );

    \I__4145\ : LocalMux
    port map (
            O => \N__18656\,
            I => \b2v_inst.N_351_0\
        );

    \I__4144\ : Odrv4
    port map (
            O => \N__18653\,
            I => \b2v_inst.N_351_0\
        );

    \I__4143\ : LocalMux
    port map (
            O => \N__18650\,
            I => \b2v_inst.N_351_0\
        );

    \I__4142\ : Odrv4
    port map (
            O => \N__18639\,
            I => \b2v_inst.N_351_0\
        );

    \I__4141\ : SRMux
    port map (
            O => \N__18620\,
            I => \N__18617\
        );

    \I__4140\ : LocalMux
    port map (
            O => \N__18617\,
            I => \N__18614\
        );

    \I__4139\ : Span4Mux_v
    port map (
            O => \N__18614\,
            I => \N__18610\
        );

    \I__4138\ : SRMux
    port map (
            O => \N__18613\,
            I => \N__18607\
        );

    \I__4137\ : Span4Mux_v
    port map (
            O => \N__18610\,
            I => \N__18596\
        );

    \I__4136\ : LocalMux
    port map (
            O => \N__18607\,
            I => \N__18596\
        );

    \I__4135\ : CascadeMux
    port map (
            O => \N__18606\,
            I => \N__18593\
        );

    \I__4134\ : CascadeMux
    port map (
            O => \N__18605\,
            I => \N__18590\
        );

    \I__4133\ : CascadeMux
    port map (
            O => \N__18604\,
            I => \N__18587\
        );

    \I__4132\ : CascadeMux
    port map (
            O => \N__18603\,
            I => \N__18584\
        );

    \I__4131\ : CascadeMux
    port map (
            O => \N__18602\,
            I => \N__18581\
        );

    \I__4130\ : CascadeMux
    port map (
            O => \N__18601\,
            I => \N__18578\
        );

    \I__4129\ : Span4Mux_h
    port map (
            O => \N__18596\,
            I => \N__18575\
        );

    \I__4128\ : InMux
    port map (
            O => \N__18593\,
            I => \N__18568\
        );

    \I__4127\ : InMux
    port map (
            O => \N__18590\,
            I => \N__18568\
        );

    \I__4126\ : InMux
    port map (
            O => \N__18587\,
            I => \N__18568\
        );

    \I__4125\ : InMux
    port map (
            O => \N__18584\,
            I => \N__18561\
        );

    \I__4124\ : InMux
    port map (
            O => \N__18581\,
            I => \N__18561\
        );

    \I__4123\ : InMux
    port map (
            O => \N__18578\,
            I => \N__18561\
        );

    \I__4122\ : Sp12to4
    port map (
            O => \N__18575\,
            I => \N__18558\
        );

    \I__4121\ : LocalMux
    port map (
            O => \N__18568\,
            I => \N__18553\
        );

    \I__4120\ : LocalMux
    port map (
            O => \N__18561\,
            I => \N__18553\
        );

    \I__4119\ : Span12Mux_v
    port map (
            O => \N__18558\,
            I => \N__18547\
        );

    \I__4118\ : Span12Mux_s11_h
    port map (
            O => \N__18553\,
            I => \N__18547\
        );

    \I__4117\ : InMux
    port map (
            O => \N__18552\,
            I => \N__18544\
        );

    \I__4116\ : Odrv12
    port map (
            O => \N__18547\,
            I => \CONSTANT_ONE_NET\
        );

    \I__4115\ : LocalMux
    port map (
            O => \N__18544\,
            I => \CONSTANT_ONE_NET\
        );

    \I__4114\ : CascadeMux
    port map (
            O => \N__18539\,
            I => \b2v_inst.N_384_cascade_\
        );

    \I__4113\ : InMux
    port map (
            O => \N__18536\,
            I => \N__18533\
        );

    \I__4112\ : LocalMux
    port map (
            O => \N__18533\,
            I => \b2v_inst.state_17_rep1_RNIN75CZ0Z3\
        );

    \I__4111\ : InMux
    port map (
            O => \N__18530\,
            I => \N__18520\
        );

    \I__4110\ : InMux
    port map (
            O => \N__18529\,
            I => \N__18520\
        );

    \I__4109\ : InMux
    port map (
            O => \N__18528\,
            I => \N__18520\
        );

    \I__4108\ : InMux
    port map (
            O => \N__18527\,
            I => \N__18517\
        );

    \I__4107\ : LocalMux
    port map (
            O => \N__18520\,
            I => \b2v_inst.un2_indice_3_0_iv_0_0_2\
        );

    \I__4106\ : LocalMux
    port map (
            O => \N__18517\,
            I => \b2v_inst.un2_indice_3_0_iv_0_0_2\
        );

    \I__4105\ : CascadeMux
    port map (
            O => \N__18512\,
            I => \b2v_inst1.m6_2_cascade_\
        );

    \I__4104\ : InMux
    port map (
            O => \N__18509\,
            I => \N__18506\
        );

    \I__4103\ : LocalMux
    port map (
            O => \N__18506\,
            I => \N__18503\
        );

    \I__4102\ : Odrv4
    port map (
            O => \N__18503\,
            I => \b2v_inst1.N_10_0\
        );

    \I__4101\ : InMux
    port map (
            O => \N__18500\,
            I => \N__18497\
        );

    \I__4100\ : LocalMux
    port map (
            O => \N__18497\,
            I => \N__18494\
        );

    \I__4099\ : Span4Mux_h
    port map (
            O => \N__18494\,
            I => \N__18491\
        );

    \I__4098\ : Odrv4
    port map (
            O => \N__18491\,
            I => \b2v_inst1.g0_7_1\
        );

    \I__4097\ : CascadeMux
    port map (
            O => \N__18488\,
            I => \b2v_inst1.g0_i_1_cascade_\
        );

    \I__4096\ : InMux
    port map (
            O => \N__18485\,
            I => \N__18482\
        );

    \I__4095\ : LocalMux
    port map (
            O => \N__18482\,
            I => \N__18479\
        );

    \I__4094\ : Odrv4
    port map (
            O => \N__18479\,
            I => \b2v_inst1.N_11_0\
        );

    \I__4093\ : InMux
    port map (
            O => \N__18476\,
            I => \N__18473\
        );

    \I__4092\ : LocalMux
    port map (
            O => \N__18473\,
            I => \N__18470\
        );

    \I__4091\ : Odrv4
    port map (
            O => \N__18470\,
            I => \b2v_inst1.N_32_mux\
        );

    \I__4090\ : CascadeMux
    port map (
            O => \N__18467\,
            I => \b2v_inst1.N_10_cascade_\
        );

    \I__4089\ : CascadeMux
    port map (
            O => \N__18464\,
            I => \b2v_inst1.g2_1_cascade_\
        );

    \I__4088\ : InMux
    port map (
            O => \N__18461\,
            I => \N__18458\
        );

    \I__4087\ : LocalMux
    port map (
            O => \N__18458\,
            I => \b2v_inst1.g2_0\
        );

    \I__4086\ : InMux
    port map (
            O => \N__18455\,
            I => \N__18452\
        );

    \I__4085\ : LocalMux
    port map (
            O => \N__18452\,
            I => \b2v_inst1.N_11_0_0\
        );

    \I__4084\ : InMux
    port map (
            O => \N__18449\,
            I => \N__18445\
        );

    \I__4083\ : InMux
    port map (
            O => \N__18448\,
            I => \N__18442\
        );

    \I__4082\ : LocalMux
    port map (
            O => \N__18445\,
            I => \b2v_inst1.N_9\
        );

    \I__4081\ : LocalMux
    port map (
            O => \N__18442\,
            I => \b2v_inst1.N_9\
        );

    \I__4080\ : CascadeMux
    port map (
            O => \N__18437\,
            I => \b2v_inst1.un1_r_Clk_Count_ac0_1_out_cascade_\
        );

    \I__4079\ : InMux
    port map (
            O => \N__18434\,
            I => \N__18431\
        );

    \I__4078\ : LocalMux
    port map (
            O => \N__18431\,
            I => \b2v_inst1.m22_ns_1\
        );

    \I__4077\ : CascadeMux
    port map (
            O => \N__18428\,
            I => \b2v_inst1.N_29_mux_cascade_\
        );

    \I__4076\ : CascadeMux
    port map (
            O => \N__18425\,
            I => \b2v_inst1.N_11_cascade_\
        );

    \I__4075\ : InMux
    port map (
            O => \N__18422\,
            I => \N__18419\
        );

    \I__4074\ : LocalMux
    port map (
            O => \N__18419\,
            I => \N__18416\
        );

    \I__4073\ : Odrv4
    port map (
            O => \N__18416\,
            I => \b2v_inst1.g0_0_i_1\
        );

    \I__4072\ : InMux
    port map (
            O => \N__18413\,
            I => \N__18410\
        );

    \I__4071\ : LocalMux
    port map (
            O => \N__18410\,
            I => \b2v_inst1.N_14_0\
        );

    \I__4070\ : CascadeMux
    port map (
            O => \N__18407\,
            I => \N__18404\
        );

    \I__4069\ : InMux
    port map (
            O => \N__18404\,
            I => \N__18401\
        );

    \I__4068\ : LocalMux
    port map (
            O => \N__18401\,
            I => \N__18398\
        );

    \I__4067\ : Odrv4
    port map (
            O => \N__18398\,
            I => \b2v_inst1.g0_0_i_0\
        );

    \I__4066\ : CascadeMux
    port map (
            O => \N__18395\,
            I => \N__18386\
        );

    \I__4065\ : CascadeMux
    port map (
            O => \N__18394\,
            I => \N__18383\
        );

    \I__4064\ : CascadeMux
    port map (
            O => \N__18393\,
            I => \N__18378\
        );

    \I__4063\ : InMux
    port map (
            O => \N__18392\,
            I => \N__18375\
        );

    \I__4062\ : InMux
    port map (
            O => \N__18391\,
            I => \N__18372\
        );

    \I__4061\ : InMux
    port map (
            O => \N__18390\,
            I => \N__18367\
        );

    \I__4060\ : InMux
    port map (
            O => \N__18389\,
            I => \N__18367\
        );

    \I__4059\ : InMux
    port map (
            O => \N__18386\,
            I => \N__18364\
        );

    \I__4058\ : InMux
    port map (
            O => \N__18383\,
            I => \N__18361\
        );

    \I__4057\ : InMux
    port map (
            O => \N__18382\,
            I => \N__18356\
        );

    \I__4056\ : InMux
    port map (
            O => \N__18381\,
            I => \N__18356\
        );

    \I__4055\ : InMux
    port map (
            O => \N__18378\,
            I => \N__18353\
        );

    \I__4054\ : LocalMux
    port map (
            O => \N__18375\,
            I => \b2v_inst.indice_1_repZ0Z1\
        );

    \I__4053\ : LocalMux
    port map (
            O => \N__18372\,
            I => \b2v_inst.indice_1_repZ0Z1\
        );

    \I__4052\ : LocalMux
    port map (
            O => \N__18367\,
            I => \b2v_inst.indice_1_repZ0Z1\
        );

    \I__4051\ : LocalMux
    port map (
            O => \N__18364\,
            I => \b2v_inst.indice_1_repZ0Z1\
        );

    \I__4050\ : LocalMux
    port map (
            O => \N__18361\,
            I => \b2v_inst.indice_1_repZ0Z1\
        );

    \I__4049\ : LocalMux
    port map (
            O => \N__18356\,
            I => \b2v_inst.indice_1_repZ0Z1\
        );

    \I__4048\ : LocalMux
    port map (
            O => \N__18353\,
            I => \b2v_inst.indice_1_repZ0Z1\
        );

    \I__4047\ : InMux
    port map (
            O => \N__18338\,
            I => \N__18333\
        );

    \I__4046\ : InMux
    port map (
            O => \N__18337\,
            I => \N__18327\
        );

    \I__4045\ : InMux
    port map (
            O => \N__18336\,
            I => \N__18324\
        );

    \I__4044\ : LocalMux
    port map (
            O => \N__18333\,
            I => \N__18321\
        );

    \I__4043\ : InMux
    port map (
            O => \N__18332\,
            I => \N__18316\
        );

    \I__4042\ : InMux
    port map (
            O => \N__18331\,
            I => \N__18316\
        );

    \I__4041\ : InMux
    port map (
            O => \N__18330\,
            I => \N__18313\
        );

    \I__4040\ : LocalMux
    port map (
            O => \N__18327\,
            I => \b2v_inst.indice_fastZ0Z_2\
        );

    \I__4039\ : LocalMux
    port map (
            O => \N__18324\,
            I => \b2v_inst.indice_fastZ0Z_2\
        );

    \I__4038\ : Odrv4
    port map (
            O => \N__18321\,
            I => \b2v_inst.indice_fastZ0Z_2\
        );

    \I__4037\ : LocalMux
    port map (
            O => \N__18316\,
            I => \b2v_inst.indice_fastZ0Z_2\
        );

    \I__4036\ : LocalMux
    port map (
            O => \N__18313\,
            I => \b2v_inst.indice_fastZ0Z_2\
        );

    \I__4035\ : CascadeMux
    port map (
            O => \N__18302\,
            I => \b2v_inst.dir_mem_215lt6_0_cascade_\
        );

    \I__4034\ : InMux
    port map (
            O => \N__18299\,
            I => \N__18296\
        );

    \I__4033\ : LocalMux
    port map (
            O => \N__18296\,
            I => \N__18293\
        );

    \I__4032\ : Span4Mux_h
    port map (
            O => \N__18293\,
            I => \N__18290\
        );

    \I__4031\ : Odrv4
    port map (
            O => \N__18290\,
            I => \b2v_inst.dir_mem_215lt8\
        );

    \I__4030\ : InMux
    port map (
            O => \N__18287\,
            I => \N__18284\
        );

    \I__4029\ : LocalMux
    port map (
            O => \N__18284\,
            I => \N__18281\
        );

    \I__4028\ : Odrv4
    port map (
            O => \N__18281\,
            I => \b2v_inst1.g0_0_i_a6_3_4\
        );

    \I__4027\ : InMux
    port map (
            O => \N__18278\,
            I => \N__18275\
        );

    \I__4026\ : LocalMux
    port map (
            O => \N__18275\,
            I => \N__18272\
        );

    \I__4025\ : Span4Mux_v
    port map (
            O => \N__18272\,
            I => \N__18269\
        );

    \I__4024\ : Span4Mux_h
    port map (
            O => \N__18269\,
            I => \N__18266\
        );

    \I__4023\ : Odrv4
    port map (
            O => \N__18266\,
            I => \b2v_inst1.r_rx_byteZ0Z_7\
        );

    \I__4022\ : CascadeMux
    port map (
            O => \N__18263\,
            I => \b2v_inst1.r_rx_byteZ0Z_7_cascade_\
        );

    \I__4021\ : InMux
    port map (
            O => \N__18260\,
            I => \N__18256\
        );

    \I__4020\ : CascadeMux
    port map (
            O => \N__18259\,
            I => \N__18252\
        );

    \I__4019\ : LocalMux
    port map (
            O => \N__18256\,
            I => \N__18248\
        );

    \I__4018\ : InMux
    port map (
            O => \N__18255\,
            I => \N__18245\
        );

    \I__4017\ : InMux
    port map (
            O => \N__18252\,
            I => \N__18240\
        );

    \I__4016\ : InMux
    port map (
            O => \N__18251\,
            I => \N__18240\
        );

    \I__4015\ : Span4Mux_h
    port map (
            O => \N__18248\,
            I => \N__18236\
        );

    \I__4014\ : LocalMux
    port map (
            O => \N__18245\,
            I => \N__18231\
        );

    \I__4013\ : LocalMux
    port map (
            O => \N__18240\,
            I => \N__18231\
        );

    \I__4012\ : InMux
    port map (
            O => \N__18239\,
            I => \N__18228\
        );

    \I__4011\ : Span4Mux_h
    port map (
            O => \N__18236\,
            I => \N__18221\
        );

    \I__4010\ : Span4Mux_v
    port map (
            O => \N__18231\,
            I => \N__18218\
        );

    \I__4009\ : LocalMux
    port map (
            O => \N__18228\,
            I => \N__18215\
        );

    \I__4008\ : InMux
    port map (
            O => \N__18227\,
            I => \N__18210\
        );

    \I__4007\ : InMux
    port map (
            O => \N__18226\,
            I => \N__18210\
        );

    \I__4006\ : InMux
    port map (
            O => \N__18225\,
            I => \N__18205\
        );

    \I__4005\ : InMux
    port map (
            O => \N__18224\,
            I => \N__18205\
        );

    \I__4004\ : Odrv4
    port map (
            O => \N__18221\,
            I => \b2v_inst1.r_Bit_IndexZ0Z_2\
        );

    \I__4003\ : Odrv4
    port map (
            O => \N__18218\,
            I => \b2v_inst1.r_Bit_IndexZ0Z_2\
        );

    \I__4002\ : Odrv12
    port map (
            O => \N__18215\,
            I => \b2v_inst1.r_Bit_IndexZ0Z_2\
        );

    \I__4001\ : LocalMux
    port map (
            O => \N__18210\,
            I => \b2v_inst1.r_Bit_IndexZ0Z_2\
        );

    \I__4000\ : LocalMux
    port map (
            O => \N__18205\,
            I => \b2v_inst1.r_Bit_IndexZ0Z_2\
        );

    \I__3999\ : CascadeMux
    port map (
            O => \N__18194\,
            I => \N__18188\
        );

    \I__3998\ : InMux
    port map (
            O => \N__18193\,
            I => \N__18179\
        );

    \I__3997\ : InMux
    port map (
            O => \N__18192\,
            I => \N__18179\
        );

    \I__3996\ : InMux
    port map (
            O => \N__18191\,
            I => \N__18176\
        );

    \I__3995\ : InMux
    port map (
            O => \N__18188\,
            I => \N__18169\
        );

    \I__3994\ : InMux
    port map (
            O => \N__18187\,
            I => \N__18169\
        );

    \I__3993\ : InMux
    port map (
            O => \N__18186\,
            I => \N__18169\
        );

    \I__3992\ : CascadeMux
    port map (
            O => \N__18185\,
            I => \N__18166\
        );

    \I__3991\ : InMux
    port map (
            O => \N__18184\,
            I => \N__18160\
        );

    \I__3990\ : LocalMux
    port map (
            O => \N__18179\,
            I => \N__18153\
        );

    \I__3989\ : LocalMux
    port map (
            O => \N__18176\,
            I => \N__18153\
        );

    \I__3988\ : LocalMux
    port map (
            O => \N__18169\,
            I => \N__18153\
        );

    \I__3987\ : InMux
    port map (
            O => \N__18166\,
            I => \N__18150\
        );

    \I__3986\ : InMux
    port map (
            O => \N__18165\,
            I => \N__18147\
        );

    \I__3985\ : InMux
    port map (
            O => \N__18164\,
            I => \N__18142\
        );

    \I__3984\ : InMux
    port map (
            O => \N__18163\,
            I => \N__18142\
        );

    \I__3983\ : LocalMux
    port map (
            O => \N__18160\,
            I => \N__18139\
        );

    \I__3982\ : Span4Mux_h
    port map (
            O => \N__18153\,
            I => \N__18136\
        );

    \I__3981\ : LocalMux
    port map (
            O => \N__18150\,
            I => \b2v_inst1.r_Bit_IndexZ0Z_0\
        );

    \I__3980\ : LocalMux
    port map (
            O => \N__18147\,
            I => \b2v_inst1.r_Bit_IndexZ0Z_0\
        );

    \I__3979\ : LocalMux
    port map (
            O => \N__18142\,
            I => \b2v_inst1.r_Bit_IndexZ0Z_0\
        );

    \I__3978\ : Odrv4
    port map (
            O => \N__18139\,
            I => \b2v_inst1.r_Bit_IndexZ0Z_0\
        );

    \I__3977\ : Odrv4
    port map (
            O => \N__18136\,
            I => \b2v_inst1.r_Bit_IndexZ0Z_0\
        );

    \I__3976\ : InMux
    port map (
            O => \N__18125\,
            I => \N__18120\
        );

    \I__3975\ : InMux
    port map (
            O => \N__18124\,
            I => \N__18114\
        );

    \I__3974\ : InMux
    port map (
            O => \N__18123\,
            I => \N__18114\
        );

    \I__3973\ : LocalMux
    port map (
            O => \N__18120\,
            I => \N__18111\
        );

    \I__3972\ : InMux
    port map (
            O => \N__18119\,
            I => \N__18108\
        );

    \I__3971\ : LocalMux
    port map (
            O => \N__18114\,
            I => \N__18105\
        );

    \I__3970\ : Span4Mux_h
    port map (
            O => \N__18111\,
            I => \N__18099\
        );

    \I__3969\ : LocalMux
    port map (
            O => \N__18108\,
            I => \N__18094\
        );

    \I__3968\ : Sp12to4
    port map (
            O => \N__18105\,
            I => \N__18094\
        );

    \I__3967\ : InMux
    port map (
            O => \N__18104\,
            I => \N__18091\
        );

    \I__3966\ : InMux
    port map (
            O => \N__18103\,
            I => \N__18083\
        );

    \I__3965\ : InMux
    port map (
            O => \N__18102\,
            I => \N__18083\
        );

    \I__3964\ : Span4Mux_h
    port map (
            O => \N__18099\,
            I => \N__18080\
        );

    \I__3963\ : Span12Mux_s10_v
    port map (
            O => \N__18094\,
            I => \N__18075\
        );

    \I__3962\ : LocalMux
    port map (
            O => \N__18091\,
            I => \N__18075\
        );

    \I__3961\ : InMux
    port map (
            O => \N__18090\,
            I => \N__18070\
        );

    \I__3960\ : InMux
    port map (
            O => \N__18089\,
            I => \N__18070\
        );

    \I__3959\ : InMux
    port map (
            O => \N__18088\,
            I => \N__18067\
        );

    \I__3958\ : LocalMux
    port map (
            O => \N__18083\,
            I => \b2v_inst1.r_Bit_IndexZ0Z_1\
        );

    \I__3957\ : Odrv4
    port map (
            O => \N__18080\,
            I => \b2v_inst1.r_Bit_IndexZ0Z_1\
        );

    \I__3956\ : Odrv12
    port map (
            O => \N__18075\,
            I => \b2v_inst1.r_Bit_IndexZ0Z_1\
        );

    \I__3955\ : LocalMux
    port map (
            O => \N__18070\,
            I => \b2v_inst1.r_Bit_IndexZ0Z_1\
        );

    \I__3954\ : LocalMux
    port map (
            O => \N__18067\,
            I => \b2v_inst1.r_Bit_IndexZ0Z_1\
        );

    \I__3953\ : CascadeMux
    port map (
            O => \N__18056\,
            I => \b2v_inst.un10_indice_2_cascade_\
        );

    \I__3952\ : InMux
    port map (
            O => \N__18053\,
            I => \N__18050\
        );

    \I__3951\ : LocalMux
    port map (
            O => \N__18050\,
            I => \b2v_inst.indice_fast_RNIDAJGZ0Z_2\
        );

    \I__3950\ : CascadeMux
    port map (
            O => \N__18047\,
            I => \b2v_inst.dir_mem_115lto6_1_cascade_\
        );

    \I__3949\ : CascadeMux
    port map (
            O => \N__18044\,
            I => \b2v_inst.un1_dir_mem_1_mb_1_7_cascade_\
        );

    \I__3948\ : InMux
    port map (
            O => \N__18041\,
            I => \N__18038\
        );

    \I__3947\ : LocalMux
    port map (
            O => \N__18038\,
            I => \N__18035\
        );

    \I__3946\ : Span4Mux_h
    port map (
            O => \N__18035\,
            I => \N__18032\
        );

    \I__3945\ : Odrv4
    port map (
            O => \N__18032\,
            I => \b2v_inst.dir_mem_1Z0Z_7\
        );

    \I__3944\ : InMux
    port map (
            O => \N__18029\,
            I => \N__18023\
        );

    \I__3943\ : InMux
    port map (
            O => \N__18028\,
            I => \N__18020\
        );

    \I__3942\ : InMux
    port map (
            O => \N__18027\,
            I => \N__18013\
        );

    \I__3941\ : InMux
    port map (
            O => \N__18026\,
            I => \N__18013\
        );

    \I__3940\ : LocalMux
    port map (
            O => \N__18023\,
            I => \N__18008\
        );

    \I__3939\ : LocalMux
    port map (
            O => \N__18020\,
            I => \N__18008\
        );

    \I__3938\ : CascadeMux
    port map (
            O => \N__18019\,
            I => \N__17999\
        );

    \I__3937\ : InMux
    port map (
            O => \N__18018\,
            I => \N__17996\
        );

    \I__3936\ : LocalMux
    port map (
            O => \N__18013\,
            I => \N__17991\
        );

    \I__3935\ : Span4Mux_v
    port map (
            O => \N__18008\,
            I => \N__17991\
        );

    \I__3934\ : InMux
    port map (
            O => \N__18007\,
            I => \N__17984\
        );

    \I__3933\ : InMux
    port map (
            O => \N__18006\,
            I => \N__17984\
        );

    \I__3932\ : InMux
    port map (
            O => \N__18005\,
            I => \N__17984\
        );

    \I__3931\ : InMux
    port map (
            O => \N__18004\,
            I => \N__17975\
        );

    \I__3930\ : InMux
    port map (
            O => \N__18003\,
            I => \N__17975\
        );

    \I__3929\ : InMux
    port map (
            O => \N__18002\,
            I => \N__17975\
        );

    \I__3928\ : InMux
    port map (
            O => \N__17999\,
            I => \N__17975\
        );

    \I__3927\ : LocalMux
    port map (
            O => \N__17996\,
            I => \N__17970\
        );

    \I__3926\ : Span4Mux_h
    port map (
            O => \N__17991\,
            I => \N__17963\
        );

    \I__3925\ : LocalMux
    port map (
            O => \N__17984\,
            I => \N__17963\
        );

    \I__3924\ : LocalMux
    port map (
            O => \N__17975\,
            I => \N__17963\
        );

    \I__3923\ : CascadeMux
    port map (
            O => \N__17974\,
            I => \N__17959\
        );

    \I__3922\ : CascadeMux
    port map (
            O => \N__17973\,
            I => \N__17955\
        );

    \I__3921\ : Span4Mux_v
    port map (
            O => \N__17970\,
            I => \N__17952\
        );

    \I__3920\ : Span4Mux_v
    port map (
            O => \N__17963\,
            I => \N__17949\
        );

    \I__3919\ : InMux
    port map (
            O => \N__17962\,
            I => \N__17946\
        );

    \I__3918\ : InMux
    port map (
            O => \N__17959\,
            I => \N__17939\
        );

    \I__3917\ : InMux
    port map (
            O => \N__17958\,
            I => \N__17939\
        );

    \I__3916\ : InMux
    port map (
            O => \N__17955\,
            I => \N__17939\
        );

    \I__3915\ : Odrv4
    port map (
            O => \N__17952\,
            I => \b2v_inst.indiceZ0Z_4\
        );

    \I__3914\ : Odrv4
    port map (
            O => \N__17949\,
            I => \b2v_inst.indiceZ0Z_4\
        );

    \I__3913\ : LocalMux
    port map (
            O => \N__17946\,
            I => \b2v_inst.indiceZ0Z_4\
        );

    \I__3912\ : LocalMux
    port map (
            O => \N__17939\,
            I => \b2v_inst.indiceZ0Z_4\
        );

    \I__3911\ : CascadeMux
    port map (
            O => \N__17930\,
            I => \N__17927\
        );

    \I__3910\ : InMux
    port map (
            O => \N__17927\,
            I => \N__17924\
        );

    \I__3909\ : LocalMux
    port map (
            O => \N__17924\,
            I => \N__17921\
        );

    \I__3908\ : Span4Mux_h
    port map (
            O => \N__17921\,
            I => \N__17918\
        );

    \I__3907\ : Odrv4
    port map (
            O => \N__17918\,
            I => \b2v_inst.un2_dir_mem_2_c5\
        );

    \I__3906\ : CascadeMux
    port map (
            O => \N__17915\,
            I => \b2v_inst.N_4_0_0_cascade_\
        );

    \I__3905\ : InMux
    port map (
            O => \N__17912\,
            I => \N__17909\
        );

    \I__3904\ : LocalMux
    port map (
            O => \N__17909\,
            I => \N__17906\
        );

    \I__3903\ : Odrv4
    port map (
            O => \N__17906\,
            I => \b2v_inst.N_8_0\
        );

    \I__3902\ : CascadeMux
    port map (
            O => \N__17903\,
            I => \b2v_inst.dir_mem_315lto8_a0_1_cascade_\
        );

    \I__3901\ : CascadeMux
    port map (
            O => \N__17900\,
            I => \N__17897\
        );

    \I__3900\ : InMux
    port map (
            O => \N__17897\,
            I => \N__17894\
        );

    \I__3899\ : LocalMux
    port map (
            O => \N__17894\,
            I => \N__17891\
        );

    \I__3898\ : Span4Mux_v
    port map (
            O => \N__17891\,
            I => \N__17888\
        );

    \I__3897\ : Span4Mux_h
    port map (
            O => \N__17888\,
            I => \N__17885\
        );

    \I__3896\ : Odrv4
    port map (
            O => \N__17885\,
            I => \b2v_inst.indice_fast_RNIRFV61Z0Z_3\
        );

    \I__3895\ : InMux
    port map (
            O => \N__17882\,
            I => \N__17879\
        );

    \I__3894\ : LocalMux
    port map (
            O => \N__17879\,
            I => \N__17876\
        );

    \I__3893\ : Span4Mux_h
    port map (
            O => \N__17876\,
            I => \N__17865\
        );

    \I__3892\ : InMux
    port map (
            O => \N__17875\,
            I => \N__17858\
        );

    \I__3891\ : InMux
    port map (
            O => \N__17874\,
            I => \N__17858\
        );

    \I__3890\ : InMux
    port map (
            O => \N__17873\,
            I => \N__17858\
        );

    \I__3889\ : InMux
    port map (
            O => \N__17872\,
            I => \N__17853\
        );

    \I__3888\ : InMux
    port map (
            O => \N__17871\,
            I => \N__17853\
        );

    \I__3887\ : InMux
    port map (
            O => \N__17870\,
            I => \N__17848\
        );

    \I__3886\ : InMux
    port map (
            O => \N__17869\,
            I => \N__17848\
        );

    \I__3885\ : InMux
    port map (
            O => \N__17868\,
            I => \N__17845\
        );

    \I__3884\ : Odrv4
    port map (
            O => \N__17865\,
            I => \b2v_inst.indice_0_repZ0Z1\
        );

    \I__3883\ : LocalMux
    port map (
            O => \N__17858\,
            I => \b2v_inst.indice_0_repZ0Z1\
        );

    \I__3882\ : LocalMux
    port map (
            O => \N__17853\,
            I => \b2v_inst.indice_0_repZ0Z1\
        );

    \I__3881\ : LocalMux
    port map (
            O => \N__17848\,
            I => \b2v_inst.indice_0_repZ0Z1\
        );

    \I__3880\ : LocalMux
    port map (
            O => \N__17845\,
            I => \b2v_inst.indice_0_repZ0Z1\
        );

    \I__3879\ : InMux
    port map (
            O => \N__17834\,
            I => \N__17831\
        );

    \I__3878\ : LocalMux
    port map (
            O => \N__17831\,
            I => \b2v_inst.indice_0_rep1_RNIFJJGZ0\
        );

    \I__3877\ : InMux
    port map (
            O => \N__17828\,
            I => \N__17825\
        );

    \I__3876\ : LocalMux
    port map (
            O => \N__17825\,
            I => \N__17820\
        );

    \I__3875\ : InMux
    port map (
            O => \N__17824\,
            I => \N__17815\
        );

    \I__3874\ : InMux
    port map (
            O => \N__17823\,
            I => \N__17815\
        );

    \I__3873\ : Span4Mux_v
    port map (
            O => \N__17820\,
            I => \N__17810\
        );

    \I__3872\ : LocalMux
    port map (
            O => \N__17815\,
            I => \N__17810\
        );

    \I__3871\ : Span4Mux_h
    port map (
            O => \N__17810\,
            I => \N__17807\
        );

    \I__3870\ : Odrv4
    port map (
            O => \N__17807\,
            I => \b2v_inst.N_410\
        );

    \I__3869\ : InMux
    port map (
            O => \N__17804\,
            I => \N__17801\
        );

    \I__3868\ : LocalMux
    port map (
            O => \N__17801\,
            I => \b2v_inst.un2_indice_3_iv_0_0_1\
        );

    \I__3867\ : InMux
    port map (
            O => \N__17798\,
            I => \N__17795\
        );

    \I__3866\ : LocalMux
    port map (
            O => \N__17795\,
            I => \N__17787\
        );

    \I__3865\ : CascadeMux
    port map (
            O => \N__17794\,
            I => \N__17783\
        );

    \I__3864\ : CascadeMux
    port map (
            O => \N__17793\,
            I => \N__17777\
        );

    \I__3863\ : CascadeMux
    port map (
            O => \N__17792\,
            I => \N__17774\
        );

    \I__3862\ : CascadeMux
    port map (
            O => \N__17791\,
            I => \N__17770\
        );

    \I__3861\ : CascadeMux
    port map (
            O => \N__17790\,
            I => \N__17765\
        );

    \I__3860\ : Span4Mux_h
    port map (
            O => \N__17787\,
            I => \N__17761\
        );

    \I__3859\ : InMux
    port map (
            O => \N__17786\,
            I => \N__17756\
        );

    \I__3858\ : InMux
    port map (
            O => \N__17783\,
            I => \N__17756\
        );

    \I__3857\ : InMux
    port map (
            O => \N__17782\,
            I => \N__17753\
        );

    \I__3856\ : InMux
    port map (
            O => \N__17781\,
            I => \N__17742\
        );

    \I__3855\ : InMux
    port map (
            O => \N__17780\,
            I => \N__17742\
        );

    \I__3854\ : InMux
    port map (
            O => \N__17777\,
            I => \N__17742\
        );

    \I__3853\ : InMux
    port map (
            O => \N__17774\,
            I => \N__17742\
        );

    \I__3852\ : InMux
    port map (
            O => \N__17773\,
            I => \N__17742\
        );

    \I__3851\ : InMux
    port map (
            O => \N__17770\,
            I => \N__17737\
        );

    \I__3850\ : InMux
    port map (
            O => \N__17769\,
            I => \N__17737\
        );

    \I__3849\ : InMux
    port map (
            O => \N__17768\,
            I => \N__17730\
        );

    \I__3848\ : InMux
    port map (
            O => \N__17765\,
            I => \N__17730\
        );

    \I__3847\ : InMux
    port map (
            O => \N__17764\,
            I => \N__17730\
        );

    \I__3846\ : Odrv4
    port map (
            O => \N__17761\,
            I => \b2v_inst.N_253_i\
        );

    \I__3845\ : LocalMux
    port map (
            O => \N__17756\,
            I => \b2v_inst.N_253_i\
        );

    \I__3844\ : LocalMux
    port map (
            O => \N__17753\,
            I => \b2v_inst.N_253_i\
        );

    \I__3843\ : LocalMux
    port map (
            O => \N__17742\,
            I => \b2v_inst.N_253_i\
        );

    \I__3842\ : LocalMux
    port map (
            O => \N__17737\,
            I => \b2v_inst.N_253_i\
        );

    \I__3841\ : LocalMux
    port map (
            O => \N__17730\,
            I => \b2v_inst.N_253_i\
        );

    \I__3840\ : InMux
    port map (
            O => \N__17717\,
            I => \N__17707\
        );

    \I__3839\ : InMux
    port map (
            O => \N__17716\,
            I => \N__17707\
        );

    \I__3838\ : InMux
    port map (
            O => \N__17715\,
            I => \N__17707\
        );

    \I__3837\ : InMux
    port map (
            O => \N__17714\,
            I => \N__17704\
        );

    \I__3836\ : LocalMux
    port map (
            O => \N__17707\,
            I => \N__17693\
        );

    \I__3835\ : LocalMux
    port map (
            O => \N__17704\,
            I => \N__17693\
        );

    \I__3834\ : InMux
    port map (
            O => \N__17703\,
            I => \N__17687\
        );

    \I__3833\ : InMux
    port map (
            O => \N__17702\,
            I => \N__17687\
        );

    \I__3832\ : CascadeMux
    port map (
            O => \N__17701\,
            I => \N__17684\
        );

    \I__3831\ : CascadeMux
    port map (
            O => \N__17700\,
            I => \N__17680\
        );

    \I__3830\ : InMux
    port map (
            O => \N__17699\,
            I => \N__17676\
        );

    \I__3829\ : InMux
    port map (
            O => \N__17698\,
            I => \N__17673\
        );

    \I__3828\ : Span4Mux_v
    port map (
            O => \N__17693\,
            I => \N__17670\
        );

    \I__3827\ : CascadeMux
    port map (
            O => \N__17692\,
            I => \N__17663\
        );

    \I__3826\ : LocalMux
    port map (
            O => \N__17687\,
            I => \N__17660\
        );

    \I__3825\ : InMux
    port map (
            O => \N__17684\,
            I => \N__17657\
        );

    \I__3824\ : InMux
    port map (
            O => \N__17683\,
            I => \N__17654\
        );

    \I__3823\ : InMux
    port map (
            O => \N__17680\,
            I => \N__17651\
        );

    \I__3822\ : InMux
    port map (
            O => \N__17679\,
            I => \N__17648\
        );

    \I__3821\ : LocalMux
    port map (
            O => \N__17676\,
            I => \N__17645\
        );

    \I__3820\ : LocalMux
    port map (
            O => \N__17673\,
            I => \N__17640\
        );

    \I__3819\ : Span4Mux_h
    port map (
            O => \N__17670\,
            I => \N__17640\
        );

    \I__3818\ : InMux
    port map (
            O => \N__17669\,
            I => \N__17636\
        );

    \I__3817\ : InMux
    port map (
            O => \N__17668\,
            I => \N__17633\
        );

    \I__3816\ : InMux
    port map (
            O => \N__17667\,
            I => \N__17628\
        );

    \I__3815\ : InMux
    port map (
            O => \N__17666\,
            I => \N__17628\
        );

    \I__3814\ : InMux
    port map (
            O => \N__17663\,
            I => \N__17625\
        );

    \I__3813\ : Span4Mux_h
    port map (
            O => \N__17660\,
            I => \N__17622\
        );

    \I__3812\ : LocalMux
    port map (
            O => \N__17657\,
            I => \N__17613\
        );

    \I__3811\ : LocalMux
    port map (
            O => \N__17654\,
            I => \N__17613\
        );

    \I__3810\ : LocalMux
    port map (
            O => \N__17651\,
            I => \N__17613\
        );

    \I__3809\ : LocalMux
    port map (
            O => \N__17648\,
            I => \N__17613\
        );

    \I__3808\ : Span4Mux_h
    port map (
            O => \N__17645\,
            I => \N__17608\
        );

    \I__3807\ : Span4Mux_v
    port map (
            O => \N__17640\,
            I => \N__17608\
        );

    \I__3806\ : InMux
    port map (
            O => \N__17639\,
            I => \N__17605\
        );

    \I__3805\ : LocalMux
    port map (
            O => \N__17636\,
            I => \b2v_inst.stateZ0Z_17\
        );

    \I__3804\ : LocalMux
    port map (
            O => \N__17633\,
            I => \b2v_inst.stateZ0Z_17\
        );

    \I__3803\ : LocalMux
    port map (
            O => \N__17628\,
            I => \b2v_inst.stateZ0Z_17\
        );

    \I__3802\ : LocalMux
    port map (
            O => \N__17625\,
            I => \b2v_inst.stateZ0Z_17\
        );

    \I__3801\ : Odrv4
    port map (
            O => \N__17622\,
            I => \b2v_inst.stateZ0Z_17\
        );

    \I__3800\ : Odrv12
    port map (
            O => \N__17613\,
            I => \b2v_inst.stateZ0Z_17\
        );

    \I__3799\ : Odrv4
    port map (
            O => \N__17608\,
            I => \b2v_inst.stateZ0Z_17\
        );

    \I__3798\ : LocalMux
    port map (
            O => \N__17605\,
            I => \b2v_inst.stateZ0Z_17\
        );

    \I__3797\ : CascadeMux
    port map (
            O => \N__17588\,
            I => \b2v_inst.un2_indice_20_0_cascade_\
        );

    \I__3796\ : InMux
    port map (
            O => \N__17585\,
            I => \N__17582\
        );

    \I__3795\ : LocalMux
    port map (
            O => \N__17582\,
            I => \N__17579\
        );

    \I__3794\ : Span4Mux_v
    port map (
            O => \N__17579\,
            I => \N__17576\
        );

    \I__3793\ : Odrv4
    port map (
            O => \N__17576\,
            I => \b2v_inst.N_4_0\
        );

    \I__3792\ : InMux
    port map (
            O => \N__17573\,
            I => \N__17569\
        );

    \I__3791\ : CascadeMux
    port map (
            O => \N__17572\,
            I => \N__17566\
        );

    \I__3790\ : LocalMux
    port map (
            O => \N__17569\,
            I => \N__17563\
        );

    \I__3789\ : InMux
    port map (
            O => \N__17566\,
            I => \N__17560\
        );

    \I__3788\ : Span4Mux_h
    port map (
            O => \N__17563\,
            I => \N__17557\
        );

    \I__3787\ : LocalMux
    port map (
            O => \N__17560\,
            I => \b2v_inst.un2_cuentalto7_3\
        );

    \I__3786\ : Odrv4
    port map (
            O => \N__17557\,
            I => \b2v_inst.un2_cuentalto7_3\
        );

    \I__3785\ : CascadeMux
    port map (
            O => \N__17552\,
            I => \b2v_inst.N_228_cascade_\
        );

    \I__3784\ : InMux
    port map (
            O => \N__17549\,
            I => \N__17546\
        );

    \I__3783\ : LocalMux
    port map (
            O => \N__17546\,
            I => \N__17543\
        );

    \I__3782\ : Span4Mux_h
    port map (
            O => \N__17543\,
            I => \N__17540\
        );

    \I__3781\ : Odrv4
    port map (
            O => \N__17540\,
            I => \b2v_inst.cuenta_RNI925FZ0Z_7\
        );

    \I__3780\ : InMux
    port map (
            O => \N__17537\,
            I => \N__17527\
        );

    \I__3779\ : InMux
    port map (
            O => \N__17536\,
            I => \N__17527\
        );

    \I__3778\ : InMux
    port map (
            O => \N__17535\,
            I => \N__17527\
        );

    \I__3777\ : InMux
    port map (
            O => \N__17534\,
            I => \N__17522\
        );

    \I__3776\ : LocalMux
    port map (
            O => \N__17527\,
            I => \N__17519\
        );

    \I__3775\ : InMux
    port map (
            O => \N__17526\,
            I => \N__17514\
        );

    \I__3774\ : InMux
    port map (
            O => \N__17525\,
            I => \N__17514\
        );

    \I__3773\ : LocalMux
    port map (
            O => \N__17522\,
            I => \b2v_inst.N_234\
        );

    \I__3772\ : Odrv4
    port map (
            O => \N__17519\,
            I => \b2v_inst.N_234\
        );

    \I__3771\ : LocalMux
    port map (
            O => \N__17514\,
            I => \b2v_inst.N_234\
        );

    \I__3770\ : InMux
    port map (
            O => \N__17507\,
            I => \N__17503\
        );

    \I__3769\ : InMux
    port map (
            O => \N__17506\,
            I => \N__17500\
        );

    \I__3768\ : LocalMux
    port map (
            O => \N__17503\,
            I => \b2v_inst.un2_indice_3_0_iv_0_a2_0_8_2_2\
        );

    \I__3767\ : LocalMux
    port map (
            O => \N__17500\,
            I => \b2v_inst.un2_indice_3_0_iv_0_a2_0_8_2_2\
        );

    \I__3766\ : InMux
    port map (
            O => \N__17495\,
            I => \N__17492\
        );

    \I__3765\ : LocalMux
    port map (
            O => \N__17492\,
            I => \b2v_inst.N_228\
        );

    \I__3764\ : CascadeMux
    port map (
            O => \N__17489\,
            I => \b2v_inst.N_383_8_cascade_\
        );

    \I__3763\ : InMux
    port map (
            O => \N__17486\,
            I => \N__17483\
        );

    \I__3762\ : LocalMux
    port map (
            O => \N__17483\,
            I => \N__17479\
        );

    \I__3761\ : InMux
    port map (
            O => \N__17482\,
            I => \N__17476\
        );

    \I__3760\ : Odrv4
    port map (
            O => \N__17479\,
            I => \b2v_inst.un2_indice_3_0_iv_0_a2_0_8_3_2\
        );

    \I__3759\ : LocalMux
    port map (
            O => \N__17476\,
            I => \b2v_inst.un2_indice_3_0_iv_0_a2_0_8_3_2\
        );

    \I__3758\ : CascadeMux
    port map (
            O => \N__17471\,
            I => \N__17468\
        );

    \I__3757\ : InMux
    port map (
            O => \N__17468\,
            I => \N__17464\
        );

    \I__3756\ : CascadeMux
    port map (
            O => \N__17467\,
            I => \N__17461\
        );

    \I__3755\ : LocalMux
    port map (
            O => \N__17464\,
            I => \N__17458\
        );

    \I__3754\ : InMux
    port map (
            O => \N__17461\,
            I => \N__17455\
        );

    \I__3753\ : Span4Mux_v
    port map (
            O => \N__17458\,
            I => \N__17452\
        );

    \I__3752\ : LocalMux
    port map (
            O => \N__17455\,
            I => \N__17449\
        );

    \I__3751\ : Odrv4
    port map (
            O => \N__17452\,
            I => \b2v_inst.un2_indice_21_s0_2\
        );

    \I__3750\ : Odrv4
    port map (
            O => \N__17449\,
            I => \b2v_inst.un2_indice_21_s0_2\
        );

    \I__3749\ : InMux
    port map (
            O => \N__17444\,
            I => \N__17441\
        );

    \I__3748\ : LocalMux
    port map (
            O => \N__17441\,
            I => \b2v_inst.un2_indice_20_2\
        );

    \I__3747\ : InMux
    port map (
            O => \N__17438\,
            I => \N__17435\
        );

    \I__3746\ : LocalMux
    port map (
            O => \N__17435\,
            I => \b2v_inst.un2_indice_21_s1_2\
        );

    \I__3745\ : CascadeMux
    port map (
            O => \N__17432\,
            I => \b2v_inst.un2_indice_3_0_iv_0_1_2_cascade_\
        );

    \I__3744\ : CascadeMux
    port map (
            O => \N__17429\,
            I => \N__17426\
        );

    \I__3743\ : InMux
    port map (
            O => \N__17426\,
            I => \N__17423\
        );

    \I__3742\ : LocalMux
    port map (
            O => \N__17423\,
            I => \N__17420\
        );

    \I__3741\ : Odrv4
    port map (
            O => \N__17420\,
            I => \b2v_inst.dir_mem_RNO_3Z0Z_4\
        );

    \I__3740\ : InMux
    port map (
            O => \N__17417\,
            I => \N__17414\
        );

    \I__3739\ : LocalMux
    port map (
            O => \N__17414\,
            I => \b2v_inst.un2_indice_0_d1_c2\
        );

    \I__3738\ : InMux
    port map (
            O => \N__17411\,
            I => \N__17404\
        );

    \I__3737\ : InMux
    port map (
            O => \N__17410\,
            I => \N__17404\
        );

    \I__3736\ : InMux
    port map (
            O => \N__17409\,
            I => \N__17401\
        );

    \I__3735\ : LocalMux
    port map (
            O => \N__17404\,
            I => \N__17395\
        );

    \I__3734\ : LocalMux
    port map (
            O => \N__17401\,
            I => \N__17392\
        );

    \I__3733\ : InMux
    port map (
            O => \N__17400\,
            I => \N__17387\
        );

    \I__3732\ : InMux
    port map (
            O => \N__17399\,
            I => \N__17384\
        );

    \I__3731\ : CascadeMux
    port map (
            O => \N__17398\,
            I => \N__17381\
        );

    \I__3730\ : Span4Mux_v
    port map (
            O => \N__17395\,
            I => \N__17377\
        );

    \I__3729\ : Span12Mux_h
    port map (
            O => \N__17392\,
            I => \N__17374\
        );

    \I__3728\ : InMux
    port map (
            O => \N__17391\,
            I => \N__17371\
        );

    \I__3727\ : InMux
    port map (
            O => \N__17390\,
            I => \N__17368\
        );

    \I__3726\ : LocalMux
    port map (
            O => \N__17387\,
            I => \N__17363\
        );

    \I__3725\ : LocalMux
    port map (
            O => \N__17384\,
            I => \N__17363\
        );

    \I__3724\ : InMux
    port map (
            O => \N__17381\,
            I => \N__17360\
        );

    \I__3723\ : InMux
    port map (
            O => \N__17380\,
            I => \N__17357\
        );

    \I__3722\ : Odrv4
    port map (
            O => \N__17377\,
            I => \b2v_inst.N_451\
        );

    \I__3721\ : Odrv12
    port map (
            O => \N__17374\,
            I => \b2v_inst.N_451\
        );

    \I__3720\ : LocalMux
    port map (
            O => \N__17371\,
            I => \b2v_inst.N_451\
        );

    \I__3719\ : LocalMux
    port map (
            O => \N__17368\,
            I => \b2v_inst.N_451\
        );

    \I__3718\ : Odrv4
    port map (
            O => \N__17363\,
            I => \b2v_inst.N_451\
        );

    \I__3717\ : LocalMux
    port map (
            O => \N__17360\,
            I => \b2v_inst.N_451\
        );

    \I__3716\ : LocalMux
    port map (
            O => \N__17357\,
            I => \b2v_inst.N_451\
        );

    \I__3715\ : CascadeMux
    port map (
            O => \N__17342\,
            I => \N__17338\
        );

    \I__3714\ : InMux
    port map (
            O => \N__17341\,
            I => \N__17335\
        );

    \I__3713\ : InMux
    port map (
            O => \N__17338\,
            I => \N__17332\
        );

    \I__3712\ : LocalMux
    port map (
            O => \N__17335\,
            I => \b2v_inst.un2_indice_21_s0_3\
        );

    \I__3711\ : LocalMux
    port map (
            O => \N__17332\,
            I => \b2v_inst.un2_indice_21_s0_3\
        );

    \I__3710\ : InMux
    port map (
            O => \N__17327\,
            I => \N__17324\
        );

    \I__3709\ : LocalMux
    port map (
            O => \N__17324\,
            I => \N__17321\
        );

    \I__3708\ : Odrv4
    port map (
            O => \N__17321\,
            I => \b2v_inst.un2_indice_20_3\
        );

    \I__3707\ : InMux
    port map (
            O => \N__17318\,
            I => \N__17315\
        );

    \I__3706\ : LocalMux
    port map (
            O => \N__17315\,
            I => \b2v_inst.un2_indice_21_s1_3\
        );

    \I__3705\ : CascadeMux
    port map (
            O => \N__17312\,
            I => \b2v_inst.un2_indice_3_0_iv_0_0_3_cascade_\
        );

    \I__3704\ : InMux
    port map (
            O => \N__17309\,
            I => \N__17306\
        );

    \I__3703\ : LocalMux
    port map (
            O => \N__17306\,
            I => \b2v_inst.dir_mem_RNO_5Z0Z_4\
        );

    \I__3702\ : InMux
    port map (
            O => \N__17303\,
            I => \N__17300\
        );

    \I__3701\ : LocalMux
    port map (
            O => \N__17300\,
            I => \b2v_inst.un2_indice_3_iv_0_1_0_5\
        );

    \I__3700\ : CascadeMux
    port map (
            O => \N__17297\,
            I => \b2v_inst1.g0_0_i_a6_2_2_cascade_\
        );

    \I__3699\ : InMux
    port map (
            O => \N__17294\,
            I => \N__17291\
        );

    \I__3698\ : LocalMux
    port map (
            O => \N__17291\,
            I => \b2v_inst1.g0_0_i_a6_2_1\
        );

    \I__3697\ : InMux
    port map (
            O => \N__17288\,
            I => \N__17285\
        );

    \I__3696\ : LocalMux
    port map (
            O => \N__17285\,
            I => \b2v_inst1.N_18\
        );

    \I__3695\ : InMux
    port map (
            O => \N__17282\,
            I => \N__17279\
        );

    \I__3694\ : LocalMux
    port map (
            O => \N__17279\,
            I => \N__17276\
        );

    \I__3693\ : Span4Mux_v
    port map (
            O => \N__17276\,
            I => \N__17273\
        );

    \I__3692\ : Odrv4
    port map (
            O => \N__17273\,
            I => \b2v_inst.dir_mem_RNO_2Z0Z_4\
        );

    \I__3691\ : CascadeMux
    port map (
            O => \N__17270\,
            I => \b2v_inst.un2_indice_3_0_i_1_4_cascade_\
        );

    \I__3690\ : InMux
    port map (
            O => \N__17267\,
            I => \N__17264\
        );

    \I__3689\ : LocalMux
    port map (
            O => \N__17264\,
            I => \N__17261\
        );

    \I__3688\ : Odrv4
    port map (
            O => \N__17261\,
            I => \b2v_inst.un2_indice_20_4\
        );

    \I__3687\ : CascadeMux
    port map (
            O => \N__17258\,
            I => \N__17255\
        );

    \I__3686\ : InMux
    port map (
            O => \N__17255\,
            I => \N__17252\
        );

    \I__3685\ : LocalMux
    port map (
            O => \N__17252\,
            I => \N__17249\
        );

    \I__3684\ : Odrv4
    port map (
            O => \N__17249\,
            I => \b2v_inst.dir_mem_RNO_2Z0Z_7\
        );

    \I__3683\ : InMux
    port map (
            O => \N__17246\,
            I => \N__17243\
        );

    \I__3682\ : LocalMux
    port map (
            O => \N__17243\,
            I => \b2v_inst.un2_indice_20_7\
        );

    \I__3681\ : CascadeMux
    port map (
            O => \N__17240\,
            I => \b2v_inst.un2_indice_3_0_iv_0_0_7_cascade_\
        );

    \I__3680\ : CascadeMux
    port map (
            O => \N__17237\,
            I => \b2v_inst1.N_7_cascade_\
        );

    \I__3679\ : InMux
    port map (
            O => \N__17234\,
            I => \N__17231\
        );

    \I__3678\ : LocalMux
    port map (
            O => \N__17231\,
            I => \b2v_inst1.g0_0_i_a6_1_2\
        );

    \I__3677\ : CascadeMux
    port map (
            O => \N__17228\,
            I => \b2v_inst1.N_9_cascade_\
        );

    \I__3676\ : InMux
    port map (
            O => \N__17225\,
            I => \N__17222\
        );

    \I__3675\ : LocalMux
    port map (
            O => \N__17222\,
            I => \N__17219\
        );

    \I__3674\ : Odrv12
    port map (
            O => \N__17219\,
            I => \b2v_inst1.g0_0_i_a6_3_5\
        );

    \I__3673\ : CascadeMux
    port map (
            O => \N__17216\,
            I => \b2v_inst1.N_19_cascade_\
        );

    \I__3672\ : InMux
    port map (
            O => \N__17213\,
            I => \N__17210\
        );

    \I__3671\ : LocalMux
    port map (
            O => \N__17210\,
            I => \N__17207\
        );

    \I__3670\ : Odrv4
    port map (
            O => \N__17207\,
            I => \b2v_inst1.N_6\
        );

    \I__3669\ : InMux
    port map (
            O => \N__17204\,
            I => \N__17201\
        );

    \I__3668\ : LocalMux
    port map (
            O => \N__17201\,
            I => \b2v_inst1.r_SM_Main_1_sqmuxa_1_0\
        );

    \I__3667\ : CascadeMux
    port map (
            O => \N__17198\,
            I => \N__17195\
        );

    \I__3666\ : InMux
    port map (
            O => \N__17195\,
            I => \N__17192\
        );

    \I__3665\ : LocalMux
    port map (
            O => \N__17192\,
            I => \b2v_inst1.g0_3_4\
        );

    \I__3664\ : InMux
    port map (
            O => \N__17189\,
            I => \N__17186\
        );

    \I__3663\ : LocalMux
    port map (
            O => \N__17186\,
            I => \N__17183\
        );

    \I__3662\ : Span4Mux_h
    port map (
            O => \N__17183\,
            I => \N__17180\
        );

    \I__3661\ : Odrv4
    port map (
            O => \N__17180\,
            I => \b2v_inst1.r_RX_Bytece_0_2\
        );

    \I__3660\ : InMux
    port map (
            O => \N__17177\,
            I => \N__17167\
        );

    \I__3659\ : InMux
    port map (
            O => \N__17176\,
            I => \N__17154\
        );

    \I__3658\ : InMux
    port map (
            O => \N__17175\,
            I => \N__17154\
        );

    \I__3657\ : InMux
    port map (
            O => \N__17174\,
            I => \N__17154\
        );

    \I__3656\ : InMux
    port map (
            O => \N__17173\,
            I => \N__17154\
        );

    \I__3655\ : InMux
    port map (
            O => \N__17172\,
            I => \N__17154\
        );

    \I__3654\ : InMux
    port map (
            O => \N__17171\,
            I => \N__17154\
        );

    \I__3653\ : InMux
    port map (
            O => \N__17170\,
            I => \N__17151\
        );

    \I__3652\ : LocalMux
    port map (
            O => \N__17167\,
            I => \N__17148\
        );

    \I__3651\ : LocalMux
    port map (
            O => \N__17154\,
            I => \N__17145\
        );

    \I__3650\ : LocalMux
    port map (
            O => \N__17151\,
            I => \N__17142\
        );

    \I__3649\ : Span4Mux_h
    port map (
            O => \N__17148\,
            I => \N__17139\
        );

    \I__3648\ : Span4Mux_h
    port map (
            O => \N__17145\,
            I => \N__17136\
        );

    \I__3647\ : Span4Mux_v
    port map (
            O => \N__17142\,
            I => \N__17133\
        );

    \I__3646\ : Odrv4
    port map (
            O => \N__17139\,
            I => \b2v_inst1.r_RX_Byte_1_sqmuxa\
        );

    \I__3645\ : Odrv4
    port map (
            O => \N__17136\,
            I => \b2v_inst1.r_RX_Byte_1_sqmuxa\
        );

    \I__3644\ : Odrv4
    port map (
            O => \N__17133\,
            I => \b2v_inst1.r_RX_Byte_1_sqmuxa\
        );

    \I__3643\ : InMux
    port map (
            O => \N__17126\,
            I => \N__17123\
        );

    \I__3642\ : LocalMux
    port map (
            O => \N__17123\,
            I => \N__17120\
        );

    \I__3641\ : Odrv12
    port map (
            O => \N__17120\,
            I => \b2v_inst1.r_RX_Bytece_0_0_0\
        );

    \I__3640\ : CascadeMux
    port map (
            O => \N__17117\,
            I => \N__17109\
        );

    \I__3639\ : InMux
    port map (
            O => \N__17116\,
            I => \N__17105\
        );

    \I__3638\ : InMux
    port map (
            O => \N__17115\,
            I => \N__17102\
        );

    \I__3637\ : InMux
    port map (
            O => \N__17114\,
            I => \N__17099\
        );

    \I__3636\ : InMux
    port map (
            O => \N__17113\,
            I => \N__17094\
        );

    \I__3635\ : InMux
    port map (
            O => \N__17112\,
            I => \N__17094\
        );

    \I__3634\ : InMux
    port map (
            O => \N__17109\,
            I => \N__17089\
        );

    \I__3633\ : InMux
    port map (
            O => \N__17108\,
            I => \N__17089\
        );

    \I__3632\ : LocalMux
    port map (
            O => \N__17105\,
            I => \N__17084\
        );

    \I__3631\ : LocalMux
    port map (
            O => \N__17102\,
            I => \N__17081\
        );

    \I__3630\ : LocalMux
    port map (
            O => \N__17099\,
            I => \N__17074\
        );

    \I__3629\ : LocalMux
    port map (
            O => \N__17094\,
            I => \N__17074\
        );

    \I__3628\ : LocalMux
    port map (
            O => \N__17089\,
            I => \N__17074\
        );

    \I__3627\ : InMux
    port map (
            O => \N__17088\,
            I => \N__17069\
        );

    \I__3626\ : InMux
    port map (
            O => \N__17087\,
            I => \N__17069\
        );

    \I__3625\ : Odrv4
    port map (
            O => \N__17084\,
            I => \b2v_inst.indice_3_repZ0Z1\
        );

    \I__3624\ : Odrv4
    port map (
            O => \N__17081\,
            I => \b2v_inst.indice_3_repZ0Z1\
        );

    \I__3623\ : Odrv12
    port map (
            O => \N__17074\,
            I => \b2v_inst.indice_3_repZ0Z1\
        );

    \I__3622\ : LocalMux
    port map (
            O => \N__17069\,
            I => \b2v_inst.indice_3_repZ0Z1\
        );

    \I__3621\ : CascadeMux
    port map (
            O => \N__17060\,
            I => \N__17057\
        );

    \I__3620\ : InMux
    port map (
            O => \N__17057\,
            I => \N__17054\
        );

    \I__3619\ : LocalMux
    port map (
            O => \N__17054\,
            I => \N__17051\
        );

    \I__3618\ : Odrv4
    port map (
            O => \N__17051\,
            I => \b2v_inst.un2_dir_mem_2_c4_d\
        );

    \I__3617\ : CascadeMux
    port map (
            O => \N__17048\,
            I => \b2v_inst.dir_mem_RNO_4Z0Z_4_cascade_\
        );

    \I__3616\ : InMux
    port map (
            O => \N__17045\,
            I => \N__17042\
        );

    \I__3615\ : LocalMux
    port map (
            O => \N__17042\,
            I => \N__17039\
        );

    \I__3614\ : Span4Mux_h
    port map (
            O => \N__17039\,
            I => \N__17036\
        );

    \I__3613\ : Odrv4
    port map (
            O => \N__17036\,
            I => \b2v_inst.indice_RNIA33NZ0Z_1\
        );

    \I__3612\ : InMux
    port map (
            O => \N__17033\,
            I => \N__17021\
        );

    \I__3611\ : InMux
    port map (
            O => \N__17032\,
            I => \N__17021\
        );

    \I__3610\ : InMux
    port map (
            O => \N__17031\,
            I => \N__17021\
        );

    \I__3609\ : InMux
    port map (
            O => \N__17030\,
            I => \N__17021\
        );

    \I__3608\ : LocalMux
    port map (
            O => \N__17021\,
            I => \N__17014\
        );

    \I__3607\ : InMux
    port map (
            O => \N__17020\,
            I => \N__17004\
        );

    \I__3606\ : InMux
    port map (
            O => \N__17019\,
            I => \N__17004\
        );

    \I__3605\ : InMux
    port map (
            O => \N__17018\,
            I => \N__17004\
        );

    \I__3604\ : InMux
    port map (
            O => \N__17017\,
            I => \N__17001\
        );

    \I__3603\ : Span4Mux_v
    port map (
            O => \N__17014\,
            I => \N__16997\
        );

    \I__3602\ : InMux
    port map (
            O => \N__17013\,
            I => \N__16994\
        );

    \I__3601\ : InMux
    port map (
            O => \N__17012\,
            I => \N__16991\
        );

    \I__3600\ : InMux
    port map (
            O => \N__17011\,
            I => \N__16988\
        );

    \I__3599\ : LocalMux
    port map (
            O => \N__17004\,
            I => \N__16985\
        );

    \I__3598\ : LocalMux
    port map (
            O => \N__17001\,
            I => \N__16982\
        );

    \I__3597\ : InMux
    port map (
            O => \N__17000\,
            I => \N__16979\
        );

    \I__3596\ : Span4Mux_h
    port map (
            O => \N__16997\,
            I => \N__16976\
        );

    \I__3595\ : LocalMux
    port map (
            O => \N__16994\,
            I => \N__16969\
        );

    \I__3594\ : LocalMux
    port map (
            O => \N__16991\,
            I => \N__16969\
        );

    \I__3593\ : LocalMux
    port map (
            O => \N__16988\,
            I => \N__16969\
        );

    \I__3592\ : Odrv4
    port map (
            O => \N__16985\,
            I => \b2v_inst.N_238\
        );

    \I__3591\ : Odrv4
    port map (
            O => \N__16982\,
            I => \b2v_inst.N_238\
        );

    \I__3590\ : LocalMux
    port map (
            O => \N__16979\,
            I => \b2v_inst.N_238\
        );

    \I__3589\ : Odrv4
    port map (
            O => \N__16976\,
            I => \b2v_inst.N_238\
        );

    \I__3588\ : Odrv12
    port map (
            O => \N__16969\,
            I => \b2v_inst.N_238\
        );

    \I__3587\ : InMux
    port map (
            O => \N__16958\,
            I => \N__16954\
        );

    \I__3586\ : InMux
    port map (
            O => \N__16957\,
            I => \N__16947\
        );

    \I__3585\ : LocalMux
    port map (
            O => \N__16954\,
            I => \N__16943\
        );

    \I__3584\ : InMux
    port map (
            O => \N__16953\,
            I => \N__16940\
        );

    \I__3583\ : InMux
    port map (
            O => \N__16952\,
            I => \N__16937\
        );

    \I__3582\ : InMux
    port map (
            O => \N__16951\,
            I => \N__16930\
        );

    \I__3581\ : InMux
    port map (
            O => \N__16950\,
            I => \N__16930\
        );

    \I__3580\ : LocalMux
    port map (
            O => \N__16947\,
            I => \N__16927\
        );

    \I__3579\ : InMux
    port map (
            O => \N__16946\,
            I => \N__16924\
        );

    \I__3578\ : Span4Mux_v
    port map (
            O => \N__16943\,
            I => \N__16921\
        );

    \I__3577\ : LocalMux
    port map (
            O => \N__16940\,
            I => \N__16916\
        );

    \I__3576\ : LocalMux
    port map (
            O => \N__16937\,
            I => \N__16916\
        );

    \I__3575\ : InMux
    port map (
            O => \N__16936\,
            I => \N__16911\
        );

    \I__3574\ : InMux
    port map (
            O => \N__16935\,
            I => \N__16911\
        );

    \I__3573\ : LocalMux
    port map (
            O => \N__16930\,
            I => \N__16906\
        );

    \I__3572\ : Span4Mux_h
    port map (
            O => \N__16927\,
            I => \N__16906\
        );

    \I__3571\ : LocalMux
    port map (
            O => \N__16924\,
            I => \b2v_inst.N_236\
        );

    \I__3570\ : Odrv4
    port map (
            O => \N__16921\,
            I => \b2v_inst.N_236\
        );

    \I__3569\ : Odrv4
    port map (
            O => \N__16916\,
            I => \b2v_inst.N_236\
        );

    \I__3568\ : LocalMux
    port map (
            O => \N__16911\,
            I => \b2v_inst.N_236\
        );

    \I__3567\ : Odrv4
    port map (
            O => \N__16906\,
            I => \b2v_inst.N_236\
        );

    \I__3566\ : CascadeMux
    port map (
            O => \N__16895\,
            I => \N__16892\
        );

    \I__3565\ : InMux
    port map (
            O => \N__16892\,
            I => \N__16889\
        );

    \I__3564\ : LocalMux
    port map (
            O => \N__16889\,
            I => \N__16886\
        );

    \I__3563\ : Span4Mux_h
    port map (
            O => \N__16886\,
            I => \N__16883\
        );

    \I__3562\ : Odrv4
    port map (
            O => \N__16883\,
            I => \b2v_inst.dir_mem_3Z0Z_2\
        );

    \I__3561\ : InMux
    port map (
            O => \N__16880\,
            I => \N__16877\
        );

    \I__3560\ : LocalMux
    port map (
            O => \N__16877\,
            I => \N__16874\
        );

    \I__3559\ : Odrv12
    port map (
            O => \N__16874\,
            I => \b2v_inst.addr_ram_1_0_iv_i_1_2\
        );

    \I__3558\ : CascadeMux
    port map (
            O => \N__16871\,
            I => \b2v_inst.un10_indice_cascade_\
        );

    \I__3557\ : InMux
    port map (
            O => \N__16868\,
            I => \N__16865\
        );

    \I__3556\ : LocalMux
    port map (
            O => \N__16865\,
            I => \b2v_inst.un2_indice_3_iv_0_a2_2_sx_5\
        );

    \I__3555\ : CascadeMux
    port map (
            O => \N__16862\,
            I => \N__16859\
        );

    \I__3554\ : InMux
    port map (
            O => \N__16859\,
            I => \N__16856\
        );

    \I__3553\ : LocalMux
    port map (
            O => \N__16856\,
            I => \N__16852\
        );

    \I__3552\ : InMux
    port map (
            O => \N__16855\,
            I => \N__16849\
        );

    \I__3551\ : Odrv4
    port map (
            O => \N__16852\,
            I => \b2v_inst.un2_indice_0_d0_c4_d\
        );

    \I__3550\ : LocalMux
    port map (
            O => \N__16849\,
            I => \b2v_inst.un2_indice_0_d0_c4_d\
        );

    \I__3549\ : CascadeMux
    port map (
            O => \N__16844\,
            I => \b2v_inst.un2_m1_e_0_cascade_\
        );

    \I__3548\ : CascadeMux
    port map (
            O => \N__16841\,
            I => \N__16838\
        );

    \I__3547\ : InMux
    port map (
            O => \N__16838\,
            I => \N__16835\
        );

    \I__3546\ : LocalMux
    port map (
            O => \N__16835\,
            I => \N__16832\
        );

    \I__3545\ : Odrv4
    port map (
            O => \N__16832\,
            I => \b2v_inst.dir_mem_RNIR93H1Z0Z_5\
        );

    \I__3544\ : CascadeMux
    port map (
            O => \N__16829\,
            I => \N__16826\
        );

    \I__3543\ : InMux
    port map (
            O => \N__16826\,
            I => \N__16823\
        );

    \I__3542\ : LocalMux
    port map (
            O => \N__16823\,
            I => \N__16820\
        );

    \I__3541\ : Span4Mux_h
    port map (
            O => \N__16820\,
            I => \N__16817\
        );

    \I__3540\ : Odrv4
    port map (
            O => \N__16817\,
            I => \b2v_inst.g1_0_3\
        );

    \I__3539\ : InMux
    port map (
            O => \N__16814\,
            I => \N__16811\
        );

    \I__3538\ : LocalMux
    port map (
            O => \N__16811\,
            I => \b2v_inst.g0_2_7\
        );

    \I__3537\ : InMux
    port map (
            O => \N__16808\,
            I => \N__16805\
        );

    \I__3536\ : LocalMux
    port map (
            O => \N__16805\,
            I => \N__16800\
        );

    \I__3535\ : InMux
    port map (
            O => \N__16804\,
            I => \N__16797\
        );

    \I__3534\ : InMux
    port map (
            O => \N__16803\,
            I => \N__16794\
        );

    \I__3533\ : Odrv4
    port map (
            O => \N__16800\,
            I => \b2v_inst.N_467\
        );

    \I__3532\ : LocalMux
    port map (
            O => \N__16797\,
            I => \b2v_inst.N_467\
        );

    \I__3531\ : LocalMux
    port map (
            O => \N__16794\,
            I => \b2v_inst.N_467\
        );

    \I__3530\ : CascadeMux
    port map (
            O => \N__16787\,
            I => \b2v_inst.N_411_cascade_\
        );

    \I__3529\ : InMux
    port map (
            O => \N__16784\,
            I => \N__16781\
        );

    \I__3528\ : LocalMux
    port map (
            O => \N__16781\,
            I => \N__16778\
        );

    \I__3527\ : Odrv4
    port map (
            O => \N__16778\,
            I => \b2v_inst.un2_indice_20_5\
        );

    \I__3526\ : InMux
    port map (
            O => \N__16775\,
            I => \b2v_inst.un2_indice_cry_6\
        );

    \I__3525\ : CascadeMux
    port map (
            O => \N__16772\,
            I => \b2v_inst.un2_indice_21_s0_1_cascade_\
        );

    \I__3524\ : CascadeMux
    port map (
            O => \N__16769\,
            I => \N__16766\
        );

    \I__3523\ : InMux
    port map (
            O => \N__16766\,
            I => \N__16763\
        );

    \I__3522\ : LocalMux
    port map (
            O => \N__16763\,
            I => \b2v_inst.un2_indice_21_s0_1\
        );

    \I__3521\ : InMux
    port map (
            O => \N__16760\,
            I => \N__16757\
        );

    \I__3520\ : LocalMux
    port map (
            O => \N__16757\,
            I => \b2v_inst.un2_indice_20_1\
        );

    \I__3519\ : InMux
    port map (
            O => \N__16754\,
            I => \N__16751\
        );

    \I__3518\ : LocalMux
    port map (
            O => \N__16751\,
            I => \b2v_inst.dir_mem_RNO_2Z0Z_1\
        );

    \I__3517\ : CascadeMux
    port map (
            O => \N__16748\,
            I => \b2v_inst.dir_mem_RNO_3Z0Z_1_cascade_\
        );

    \I__3516\ : CascadeMux
    port map (
            O => \N__16745\,
            I => \N__16742\
        );

    \I__3515\ : InMux
    port map (
            O => \N__16742\,
            I => \N__16739\
        );

    \I__3514\ : LocalMux
    port map (
            O => \N__16739\,
            I => \N__16736\
        );

    \I__3513\ : Odrv4
    port map (
            O => \N__16736\,
            I => \b2v_inst.dir_mem_RNIP73H1Z0Z_4\
        );

    \I__3512\ : InMux
    port map (
            O => \N__16733\,
            I => \N__16729\
        );

    \I__3511\ : InMux
    port map (
            O => \N__16732\,
            I => \N__16726\
        );

    \I__3510\ : LocalMux
    port map (
            O => \N__16729\,
            I => \N__16719\
        );

    \I__3509\ : LocalMux
    port map (
            O => \N__16726\,
            I => \N__16716\
        );

    \I__3508\ : InMux
    port map (
            O => \N__16725\,
            I => \N__16713\
        );

    \I__3507\ : InMux
    port map (
            O => \N__16724\,
            I => \N__16706\
        );

    \I__3506\ : InMux
    port map (
            O => \N__16723\,
            I => \N__16706\
        );

    \I__3505\ : InMux
    port map (
            O => \N__16722\,
            I => \N__16706\
        );

    \I__3504\ : Odrv4
    port map (
            O => \N__16719\,
            I => \b2v_inst.dir_mem_215_0\
        );

    \I__3503\ : Odrv4
    port map (
            O => \N__16716\,
            I => \b2v_inst.dir_mem_215_0\
        );

    \I__3502\ : LocalMux
    port map (
            O => \N__16713\,
            I => \b2v_inst.dir_mem_215_0\
        );

    \I__3501\ : LocalMux
    port map (
            O => \N__16706\,
            I => \b2v_inst.dir_mem_215_0\
        );

    \I__3500\ : CascadeMux
    port map (
            O => \N__16697\,
            I => \N__16694\
        );

    \I__3499\ : InMux
    port map (
            O => \N__16694\,
            I => \N__16691\
        );

    \I__3498\ : LocalMux
    port map (
            O => \N__16691\,
            I => \N__16688\
        );

    \I__3497\ : Span4Mux_v
    port map (
            O => \N__16688\,
            I => \N__16685\
        );

    \I__3496\ : Odrv4
    port map (
            O => \N__16685\,
            I => \b2v_inst.dir_mem_2Z0Z_5\
        );

    \I__3495\ : CEMux
    port map (
            O => \N__16682\,
            I => \N__16679\
        );

    \I__3494\ : LocalMux
    port map (
            O => \N__16679\,
            I => \N__16674\
        );

    \I__3493\ : CEMux
    port map (
            O => \N__16678\,
            I => \N__16670\
        );

    \I__3492\ : CEMux
    port map (
            O => \N__16677\,
            I => \N__16667\
        );

    \I__3491\ : Span4Mux_v
    port map (
            O => \N__16674\,
            I => \N__16664\
        );

    \I__3490\ : CEMux
    port map (
            O => \N__16673\,
            I => \N__16661\
        );

    \I__3489\ : LocalMux
    port map (
            O => \N__16670\,
            I => \N__16656\
        );

    \I__3488\ : LocalMux
    port map (
            O => \N__16667\,
            I => \N__16656\
        );

    \I__3487\ : Span4Mux_h
    port map (
            O => \N__16664\,
            I => \N__16651\
        );

    \I__3486\ : LocalMux
    port map (
            O => \N__16661\,
            I => \N__16651\
        );

    \I__3485\ : Span4Mux_v
    port map (
            O => \N__16656\,
            I => \N__16648\
        );

    \I__3484\ : Span4Mux_h
    port map (
            O => \N__16651\,
            I => \N__16645\
        );

    \I__3483\ : Span4Mux_h
    port map (
            O => \N__16648\,
            I => \N__16642\
        );

    \I__3482\ : Span4Mux_h
    port map (
            O => \N__16645\,
            I => \N__16639\
        );

    \I__3481\ : Odrv4
    port map (
            O => \N__16642\,
            I => \b2v_inst.N_136_i\
        );

    \I__3480\ : Odrv4
    port map (
            O => \N__16639\,
            I => \b2v_inst.N_136_i\
        );

    \I__3479\ : InMux
    port map (
            O => \N__16634\,
            I => \N__16628\
        );

    \I__3478\ : InMux
    port map (
            O => \N__16633\,
            I => \N__16628\
        );

    \I__3477\ : LocalMux
    port map (
            O => \N__16628\,
            I => \b2v_inst1.N_14\
        );

    \I__3476\ : CascadeMux
    port map (
            O => \N__16625\,
            I => \N__16622\
        );

    \I__3475\ : InMux
    port map (
            O => \N__16622\,
            I => \N__16619\
        );

    \I__3474\ : LocalMux
    port map (
            O => \N__16619\,
            I => \b2v_inst.dir_mem_RNIGVEE1Z0Z_0\
        );

    \I__3473\ : InMux
    port map (
            O => \N__16616\,
            I => \N__16613\
        );

    \I__3472\ : LocalMux
    port map (
            O => \N__16613\,
            I => \b2v_inst.dir_mem_RNII5PO1Z0Z_1\
        );

    \I__3471\ : InMux
    port map (
            O => \N__16610\,
            I => \b2v_inst.un2_indice_cry_0\
        );

    \I__3470\ : InMux
    port map (
            O => \N__16607\,
            I => \N__16604\
        );

    \I__3469\ : LocalMux
    port map (
            O => \N__16604\,
            I => \b2v_inst.dir_mem_RNIL33H1Z0Z_2\
        );

    \I__3468\ : InMux
    port map (
            O => \N__16601\,
            I => \b2v_inst.un2_indice_cry_1\
        );

    \I__3467\ : InMux
    port map (
            O => \N__16598\,
            I => \N__16595\
        );

    \I__3466\ : LocalMux
    port map (
            O => \N__16595\,
            I => \b2v_inst.dir_mem_RNIN53H1Z0Z_3\
        );

    \I__3465\ : InMux
    port map (
            O => \N__16592\,
            I => \b2v_inst.un2_indice_cry_2\
        );

    \I__3464\ : InMux
    port map (
            O => \N__16589\,
            I => \b2v_inst.un2_indice_cry_3\
        );

    \I__3463\ : InMux
    port map (
            O => \N__16586\,
            I => \b2v_inst.un2_indice_cry_4\
        );

    \I__3462\ : CascadeMux
    port map (
            O => \N__16583\,
            I => \N__16580\
        );

    \I__3461\ : InMux
    port map (
            O => \N__16580\,
            I => \N__16577\
        );

    \I__3460\ : LocalMux
    port map (
            O => \N__16577\,
            I => \b2v_inst.dir_mem_RNITB3H1Z0Z_6\
        );

    \I__3459\ : InMux
    port map (
            O => \N__16574\,
            I => \N__16571\
        );

    \I__3458\ : LocalMux
    port map (
            O => \N__16571\,
            I => \b2v_inst.un2_indice_20_6\
        );

    \I__3457\ : InMux
    port map (
            O => \N__16568\,
            I => \b2v_inst.un2_indice_cry_5\
        );

    \I__3456\ : CascadeMux
    port map (
            O => \N__16565\,
            I => \N__16562\
        );

    \I__3455\ : InMux
    port map (
            O => \N__16562\,
            I => \N__16559\
        );

    \I__3454\ : LocalMux
    port map (
            O => \N__16559\,
            I => \b2v_inst.m7_1\
        );

    \I__3453\ : CascadeMux
    port map (
            O => \N__16556\,
            I => \b2v_inst.un8_dir_mem_3_c4_cascade_\
        );

    \I__3452\ : InMux
    port map (
            O => \N__16553\,
            I => \N__16550\
        );

    \I__3451\ : LocalMux
    port map (
            O => \N__16550\,
            I => \N__16547\
        );

    \I__3450\ : Odrv4
    port map (
            O => \N__16547\,
            I => \b2v_inst.un8_dir_mem_3_c6\
        );

    \I__3449\ : CascadeMux
    port map (
            O => \N__16544\,
            I => \b2v_inst.un2_indice_1_1_4_cascade_\
        );

    \I__3448\ : CascadeMux
    port map (
            O => \N__16541\,
            I => \N__16538\
        );

    \I__3447\ : InMux
    port map (
            O => \N__16538\,
            I => \N__16535\
        );

    \I__3446\ : LocalMux
    port map (
            O => \N__16535\,
            I => \N__16532\
        );

    \I__3445\ : Span4Mux_h
    port map (
            O => \N__16532\,
            I => \N__16529\
        );

    \I__3444\ : Odrv4
    port map (
            O => \N__16529\,
            I => \b2v_inst.dir_mem_2Z0Z_4\
        );

    \I__3443\ : CascadeMux
    port map (
            O => \N__16526\,
            I => \N__16523\
        );

    \I__3442\ : InMux
    port map (
            O => \N__16523\,
            I => \N__16520\
        );

    \I__3441\ : LocalMux
    port map (
            O => \N__16520\,
            I => \N__16517\
        );

    \I__3440\ : Span4Mux_h
    port map (
            O => \N__16517\,
            I => \N__16514\
        );

    \I__3439\ : Sp12to4
    port map (
            O => \N__16514\,
            I => \N__16511\
        );

    \I__3438\ : Odrv12
    port map (
            O => \N__16511\,
            I => \b2v_inst.dir_mem_2Z0Z_1\
        );

    \I__3437\ : InMux
    port map (
            O => \N__16508\,
            I => \N__16505\
        );

    \I__3436\ : LocalMux
    port map (
            O => \N__16505\,
            I => \N__16502\
        );

    \I__3435\ : Span4Mux_v
    port map (
            O => \N__16502\,
            I => \N__16499\
        );

    \I__3434\ : Odrv4
    port map (
            O => \N__16499\,
            I => \b2v_inst.dir_mem_2Z0Z_2\
        );

    \I__3433\ : CascadeMux
    port map (
            O => \N__16496\,
            I => \b2v_inst.dir_mem_215_0_cascade_\
        );

    \I__3432\ : InMux
    port map (
            O => \N__16493\,
            I => \N__16490\
        );

    \I__3431\ : LocalMux
    port map (
            O => \N__16490\,
            I => \N__16487\
        );

    \I__3430\ : Span4Mux_v
    port map (
            O => \N__16487\,
            I => \N__16484\
        );

    \I__3429\ : Odrv4
    port map (
            O => \N__16484\,
            I => \b2v_inst.dir_mem_2Z0Z_0\
        );

    \I__3428\ : InMux
    port map (
            O => \N__16481\,
            I => \N__16475\
        );

    \I__3427\ : CascadeMux
    port map (
            O => \N__16480\,
            I => \N__16470\
        );

    \I__3426\ : CascadeMux
    port map (
            O => \N__16479\,
            I => \N__16467\
        );

    \I__3425\ : InMux
    port map (
            O => \N__16478\,
            I => \N__16462\
        );

    \I__3424\ : LocalMux
    port map (
            O => \N__16475\,
            I => \N__16459\
        );

    \I__3423\ : InMux
    port map (
            O => \N__16474\,
            I => \N__16455\
        );

    \I__3422\ : InMux
    port map (
            O => \N__16473\,
            I => \N__16452\
        );

    \I__3421\ : InMux
    port map (
            O => \N__16470\,
            I => \N__16445\
        );

    \I__3420\ : InMux
    port map (
            O => \N__16467\,
            I => \N__16445\
        );

    \I__3419\ : InMux
    port map (
            O => \N__16466\,
            I => \N__16445\
        );

    \I__3418\ : InMux
    port map (
            O => \N__16465\,
            I => \N__16442\
        );

    \I__3417\ : LocalMux
    port map (
            O => \N__16462\,
            I => \N__16437\
        );

    \I__3416\ : Span4Mux_v
    port map (
            O => \N__16459\,
            I => \N__16437\
        );

    \I__3415\ : InMux
    port map (
            O => \N__16458\,
            I => \N__16434\
        );

    \I__3414\ : LocalMux
    port map (
            O => \N__16455\,
            I => \N__16431\
        );

    \I__3413\ : LocalMux
    port map (
            O => \N__16452\,
            I => \b2v_inst.N_237\
        );

    \I__3412\ : LocalMux
    port map (
            O => \N__16445\,
            I => \b2v_inst.N_237\
        );

    \I__3411\ : LocalMux
    port map (
            O => \N__16442\,
            I => \b2v_inst.N_237\
        );

    \I__3410\ : Odrv4
    port map (
            O => \N__16437\,
            I => \b2v_inst.N_237\
        );

    \I__3409\ : LocalMux
    port map (
            O => \N__16434\,
            I => \b2v_inst.N_237\
        );

    \I__3408\ : Odrv4
    port map (
            O => \N__16431\,
            I => \b2v_inst.N_237\
        );

    \I__3407\ : CascadeMux
    port map (
            O => \N__16418\,
            I => \N__16415\
        );

    \I__3406\ : InMux
    port map (
            O => \N__16415\,
            I => \N__16412\
        );

    \I__3405\ : LocalMux
    port map (
            O => \N__16412\,
            I => \b2v_inst.dir_mem_2Z0Z_7\
        );

    \I__3404\ : InMux
    port map (
            O => \N__16409\,
            I => \N__16406\
        );

    \I__3403\ : LocalMux
    port map (
            O => \N__16406\,
            I => \N__16402\
        );

    \I__3402\ : CascadeMux
    port map (
            O => \N__16405\,
            I => \N__16397\
        );

    \I__3401\ : Span4Mux_h
    port map (
            O => \N__16402\,
            I => \N__16391\
        );

    \I__3400\ : InMux
    port map (
            O => \N__16401\,
            I => \N__16388\
        );

    \I__3399\ : InMux
    port map (
            O => \N__16400\,
            I => \N__16381\
        );

    \I__3398\ : InMux
    port map (
            O => \N__16397\,
            I => \N__16381\
        );

    \I__3397\ : InMux
    port map (
            O => \N__16396\,
            I => \N__16381\
        );

    \I__3396\ : InMux
    port map (
            O => \N__16395\,
            I => \N__16378\
        );

    \I__3395\ : InMux
    port map (
            O => \N__16394\,
            I => \N__16375\
        );

    \I__3394\ : Span4Mux_v
    port map (
            O => \N__16391\,
            I => \N__16371\
        );

    \I__3393\ : LocalMux
    port map (
            O => \N__16388\,
            I => \N__16368\
        );

    \I__3392\ : LocalMux
    port map (
            O => \N__16381\,
            I => \N__16361\
        );

    \I__3391\ : LocalMux
    port map (
            O => \N__16378\,
            I => \N__16361\
        );

    \I__3390\ : LocalMux
    port map (
            O => \N__16375\,
            I => \N__16361\
        );

    \I__3389\ : InMux
    port map (
            O => \N__16374\,
            I => \N__16358\
        );

    \I__3388\ : Odrv4
    port map (
            O => \N__16371\,
            I => \b2v_inst.N_239\
        );

    \I__3387\ : Odrv4
    port map (
            O => \N__16368\,
            I => \b2v_inst.N_239\
        );

    \I__3386\ : Odrv4
    port map (
            O => \N__16361\,
            I => \b2v_inst.N_239\
        );

    \I__3385\ : LocalMux
    port map (
            O => \N__16358\,
            I => \b2v_inst.N_239\
        );

    \I__3384\ : CascadeMux
    port map (
            O => \N__16349\,
            I => \b2v_inst.addr_ram_1_0_iv_i_1_7_cascade_\
        );

    \I__3383\ : InMux
    port map (
            O => \N__16346\,
            I => \N__16343\
        );

    \I__3382\ : LocalMux
    port map (
            O => \N__16343\,
            I => \N__16340\
        );

    \I__3381\ : Span4Mux_h
    port map (
            O => \N__16340\,
            I => \N__16337\
        );

    \I__3380\ : Odrv4
    port map (
            O => \N__16337\,
            I => \b2v_inst.addr_ram_1_0_iv_i_0_7\
        );

    \I__3379\ : CascadeMux
    port map (
            O => \N__16334\,
            I => \N__16331\
        );

    \I__3378\ : InMux
    port map (
            O => \N__16331\,
            I => \N__16327\
        );

    \I__3377\ : CascadeMux
    port map (
            O => \N__16330\,
            I => \N__16324\
        );

    \I__3376\ : LocalMux
    port map (
            O => \N__16327\,
            I => \N__16321\
        );

    \I__3375\ : InMux
    port map (
            O => \N__16324\,
            I => \N__16318\
        );

    \I__3374\ : Span4Mux_h
    port map (
            O => \N__16321\,
            I => \N__16315\
        );

    \I__3373\ : LocalMux
    port map (
            O => \N__16318\,
            I => \N__16312\
        );

    \I__3372\ : Span4Mux_h
    port map (
            O => \N__16315\,
            I => \N__16309\
        );

    \I__3371\ : Odrv12
    port map (
            O => \N__16312\,
            I => \N_50\
        );

    \I__3370\ : Odrv4
    port map (
            O => \N__16309\,
            I => \N_50\
        );

    \I__3369\ : CascadeMux
    port map (
            O => \N__16304\,
            I => \b2v_inst.g0_2_6_cascade_\
        );

    \I__3368\ : InMux
    port map (
            O => \N__16301\,
            I => \N__16298\
        );

    \I__3367\ : LocalMux
    port map (
            O => \N__16298\,
            I => \N__16295\
        );

    \I__3366\ : Span4Mux_h
    port map (
            O => \N__16295\,
            I => \N__16292\
        );

    \I__3365\ : Odrv4
    port map (
            O => \N__16292\,
            I => \b2v_inst.g0_2_8\
        );

    \I__3364\ : CascadeMux
    port map (
            O => \N__16289\,
            I => \b2v_inst.i4_mux_cascade_\
        );

    \I__3363\ : InMux
    port map (
            O => \N__16286\,
            I => \N__16283\
        );

    \I__3362\ : LocalMux
    port map (
            O => \N__16283\,
            I => \N__16280\
        );

    \I__3361\ : Span4Mux_h
    port map (
            O => \N__16280\,
            I => \N__16277\
        );

    \I__3360\ : Odrv4
    port map (
            O => \N__16277\,
            I => \b2v_inst.dir_mem_1Z0Z_6\
        );

    \I__3359\ : InMux
    port map (
            O => \N__16274\,
            I => \N__16271\
        );

    \I__3358\ : LocalMux
    port map (
            O => \N__16271\,
            I => \N__16267\
        );

    \I__3357\ : InMux
    port map (
            O => \N__16270\,
            I => \N__16264\
        );

    \I__3356\ : Odrv4
    port map (
            O => \N__16267\,
            I => \b2v_inst.un2_dir_mem_3_c5\
        );

    \I__3355\ : LocalMux
    port map (
            O => \N__16264\,
            I => \b2v_inst.un2_dir_mem_3_c5\
        );

    \I__3354\ : CascadeMux
    port map (
            O => \N__16259\,
            I => \N__16256\
        );

    \I__3353\ : InMux
    port map (
            O => \N__16256\,
            I => \N__16253\
        );

    \I__3352\ : LocalMux
    port map (
            O => \N__16253\,
            I => \b2v_inst.un2_dir_mem_3_ac0_3\
        );

    \I__3351\ : CascadeMux
    port map (
            O => \N__16250\,
            I => \b2v_inst.un2_dir_mem_3_ac0_3_cascade_\
        );

    \I__3350\ : InMux
    port map (
            O => \N__16247\,
            I => \N__16244\
        );

    \I__3349\ : LocalMux
    port map (
            O => \N__16244\,
            I => \N__16241\
        );

    \I__3348\ : Odrv4
    port map (
            O => \N__16241\,
            I => \b2v_inst.un1_dir_mem_3_ns_1_5\
        );

    \I__3347\ : CascadeMux
    port map (
            O => \N__16238\,
            I => \b2v_inst.g4_0_cascade_\
        );

    \I__3346\ : InMux
    port map (
            O => \N__16235\,
            I => \N__16232\
        );

    \I__3345\ : LocalMux
    port map (
            O => \N__16232\,
            I => \b2v_inst.g0_0\
        );

    \I__3344\ : CascadeMux
    port map (
            O => \N__16229\,
            I => \N__16225\
        );

    \I__3343\ : InMux
    port map (
            O => \N__16228\,
            I => \N__16218\
        );

    \I__3342\ : InMux
    port map (
            O => \N__16225\,
            I => \N__16214\
        );

    \I__3341\ : InMux
    port map (
            O => \N__16224\,
            I => \N__16211\
        );

    \I__3340\ : InMux
    port map (
            O => \N__16223\,
            I => \N__16206\
        );

    \I__3339\ : InMux
    port map (
            O => \N__16222\,
            I => \N__16206\
        );

    \I__3338\ : InMux
    port map (
            O => \N__16221\,
            I => \N__16203\
        );

    \I__3337\ : LocalMux
    port map (
            O => \N__16218\,
            I => \N__16199\
        );

    \I__3336\ : InMux
    port map (
            O => \N__16217\,
            I => \N__16196\
        );

    \I__3335\ : LocalMux
    port map (
            O => \N__16214\,
            I => \N__16187\
        );

    \I__3334\ : LocalMux
    port map (
            O => \N__16211\,
            I => \N__16187\
        );

    \I__3333\ : LocalMux
    port map (
            O => \N__16206\,
            I => \N__16187\
        );

    \I__3332\ : LocalMux
    port map (
            O => \N__16203\,
            I => \N__16187\
        );

    \I__3331\ : InMux
    port map (
            O => \N__16202\,
            I => \N__16184\
        );

    \I__3330\ : Odrv4
    port map (
            O => \N__16199\,
            I => \b2v_inst.state_ns_a2_0_o2_1_0_2\
        );

    \I__3329\ : LocalMux
    port map (
            O => \N__16196\,
            I => \b2v_inst.state_ns_a2_0_o2_1_0_2\
        );

    \I__3328\ : Odrv4
    port map (
            O => \N__16187\,
            I => \b2v_inst.state_ns_a2_0_o2_1_0_2\
        );

    \I__3327\ : LocalMux
    port map (
            O => \N__16184\,
            I => \b2v_inst.state_ns_a2_0_o2_1_0_2\
        );

    \I__3326\ : InMux
    port map (
            O => \N__16175\,
            I => \N__16165\
        );

    \I__3325\ : InMux
    port map (
            O => \N__16174\,
            I => \N__16162\
        );

    \I__3324\ : InMux
    port map (
            O => \N__16173\,
            I => \N__16159\
        );

    \I__3323\ : InMux
    port map (
            O => \N__16172\,
            I => \N__16152\
        );

    \I__3322\ : InMux
    port map (
            O => \N__16171\,
            I => \N__16152\
        );

    \I__3321\ : InMux
    port map (
            O => \N__16170\,
            I => \N__16152\
        );

    \I__3320\ : InMux
    port map (
            O => \N__16169\,
            I => \N__16147\
        );

    \I__3319\ : InMux
    port map (
            O => \N__16168\,
            I => \N__16144\
        );

    \I__3318\ : LocalMux
    port map (
            O => \N__16165\,
            I => \N__16141\
        );

    \I__3317\ : LocalMux
    port map (
            O => \N__16162\,
            I => \N__16138\
        );

    \I__3316\ : LocalMux
    port map (
            O => \N__16159\,
            I => \N__16133\
        );

    \I__3315\ : LocalMux
    port map (
            O => \N__16152\,
            I => \N__16133\
        );

    \I__3314\ : InMux
    port map (
            O => \N__16151\,
            I => \N__16128\
        );

    \I__3313\ : InMux
    port map (
            O => \N__16150\,
            I => \N__16128\
        );

    \I__3312\ : LocalMux
    port map (
            O => \N__16147\,
            I => \b2v_inst.cuenta_RNI4SC81Z0Z_7\
        );

    \I__3311\ : LocalMux
    port map (
            O => \N__16144\,
            I => \b2v_inst.cuenta_RNI4SC81Z0Z_7\
        );

    \I__3310\ : Odrv4
    port map (
            O => \N__16141\,
            I => \b2v_inst.cuenta_RNI4SC81Z0Z_7\
        );

    \I__3309\ : Odrv12
    port map (
            O => \N__16138\,
            I => \b2v_inst.cuenta_RNI4SC81Z0Z_7\
        );

    \I__3308\ : Odrv4
    port map (
            O => \N__16133\,
            I => \b2v_inst.cuenta_RNI4SC81Z0Z_7\
        );

    \I__3307\ : LocalMux
    port map (
            O => \N__16128\,
            I => \b2v_inst.cuenta_RNI4SC81Z0Z_7\
        );

    \I__3306\ : CascadeMux
    port map (
            O => \N__16115\,
            I => \N__16108\
        );

    \I__3305\ : CascadeMux
    port map (
            O => \N__16114\,
            I => \N__16105\
        );

    \I__3304\ : CascadeMux
    port map (
            O => \N__16113\,
            I => \N__16102\
        );

    \I__3303\ : CascadeMux
    port map (
            O => \N__16112\,
            I => \N__16097\
        );

    \I__3302\ : InMux
    port map (
            O => \N__16111\,
            I => \N__16094\
        );

    \I__3301\ : InMux
    port map (
            O => \N__16108\,
            I => \N__16091\
        );

    \I__3300\ : InMux
    port map (
            O => \N__16105\,
            I => \N__16088\
        );

    \I__3299\ : InMux
    port map (
            O => \N__16102\,
            I => \N__16085\
        );

    \I__3298\ : InMux
    port map (
            O => \N__16101\,
            I => \N__16078\
        );

    \I__3297\ : InMux
    port map (
            O => \N__16100\,
            I => \N__16078\
        );

    \I__3296\ : InMux
    port map (
            O => \N__16097\,
            I => \N__16078\
        );

    \I__3295\ : LocalMux
    port map (
            O => \N__16094\,
            I => \N__16069\
        );

    \I__3294\ : LocalMux
    port map (
            O => \N__16091\,
            I => \N__16069\
        );

    \I__3293\ : LocalMux
    port map (
            O => \N__16088\,
            I => \N__16069\
        );

    \I__3292\ : LocalMux
    port map (
            O => \N__16085\,
            I => \N__16064\
        );

    \I__3291\ : LocalMux
    port map (
            O => \N__16078\,
            I => \N__16064\
        );

    \I__3290\ : InMux
    port map (
            O => \N__16077\,
            I => \N__16059\
        );

    \I__3289\ : InMux
    port map (
            O => \N__16076\,
            I => \N__16059\
        );

    \I__3288\ : Span4Mux_v
    port map (
            O => \N__16069\,
            I => \N__16056\
        );

    \I__3287\ : Span4Mux_h
    port map (
            O => \N__16064\,
            I => \N__16051\
        );

    \I__3286\ : LocalMux
    port map (
            O => \N__16059\,
            I => \N__16051\
        );

    \I__3285\ : Odrv4
    port map (
            O => \N__16056\,
            I => \b2v_inst.state_ns_a2_0_o2_0_2\
        );

    \I__3284\ : Odrv4
    port map (
            O => \N__16051\,
            I => \b2v_inst.state_ns_a2_0_o2_0_2\
        );

    \I__3283\ : CEMux
    port map (
            O => \N__16046\,
            I => \N__16041\
        );

    \I__3282\ : CEMux
    port map (
            O => \N__16045\,
            I => \N__16038\
        );

    \I__3281\ : CascadeMux
    port map (
            O => \N__16044\,
            I => \N__16034\
        );

    \I__3280\ : LocalMux
    port map (
            O => \N__16041\,
            I => \N__16031\
        );

    \I__3279\ : LocalMux
    port map (
            O => \N__16038\,
            I => \N__16028\
        );

    \I__3278\ : InMux
    port map (
            O => \N__16037\,
            I => \N__16025\
        );

    \I__3277\ : InMux
    port map (
            O => \N__16034\,
            I => \N__16020\
        );

    \I__3276\ : Span4Mux_h
    port map (
            O => \N__16031\,
            I => \N__16017\
        );

    \I__3275\ : Span4Mux_h
    port map (
            O => \N__16028\,
            I => \N__16014\
        );

    \I__3274\ : LocalMux
    port map (
            O => \N__16025\,
            I => \N__16011\
        );

    \I__3273\ : InMux
    port map (
            O => \N__16024\,
            I => \N__16008\
        );

    \I__3272\ : InMux
    port map (
            O => \N__16023\,
            I => \N__16005\
        );

    \I__3271\ : LocalMux
    port map (
            O => \N__16020\,
            I => \b2v_inst.stateZ0Z_8\
        );

    \I__3270\ : Odrv4
    port map (
            O => \N__16017\,
            I => \b2v_inst.stateZ0Z_8\
        );

    \I__3269\ : Odrv4
    port map (
            O => \N__16014\,
            I => \b2v_inst.stateZ0Z_8\
        );

    \I__3268\ : Odrv4
    port map (
            O => \N__16011\,
            I => \b2v_inst.stateZ0Z_8\
        );

    \I__3267\ : LocalMux
    port map (
            O => \N__16008\,
            I => \b2v_inst.stateZ0Z_8\
        );

    \I__3266\ : LocalMux
    port map (
            O => \N__16005\,
            I => \b2v_inst.stateZ0Z_8\
        );

    \I__3265\ : CascadeMux
    port map (
            O => \N__15992\,
            I => \b2v_inst.dir_mem_2_RNO_0Z0Z_3_cascade_\
        );

    \I__3264\ : InMux
    port map (
            O => \N__15989\,
            I => \N__15986\
        );

    \I__3263\ : LocalMux
    port map (
            O => \N__15986\,
            I => \N__15983\
        );

    \I__3262\ : Odrv4
    port map (
            O => \N__15983\,
            I => \b2v_inst.dir_mem_2Z0Z_3\
        );

    \I__3261\ : CascadeMux
    port map (
            O => \N__15980\,
            I => \N__15977\
        );

    \I__3260\ : InMux
    port map (
            O => \N__15977\,
            I => \N__15974\
        );

    \I__3259\ : LocalMux
    port map (
            O => \N__15974\,
            I => \N__15971\
        );

    \I__3258\ : Span4Mux_h
    port map (
            O => \N__15971\,
            I => \N__15968\
        );

    \I__3257\ : Odrv4
    port map (
            O => \N__15968\,
            I => \b2v_inst.un1_dir_mem_3_ns_1_4\
        );

    \I__3256\ : InMux
    port map (
            O => \N__15965\,
            I => \N__15962\
        );

    \I__3255\ : LocalMux
    port map (
            O => \N__15962\,
            I => \b2v_inst.dir_mem_2_RNO_0Z0Z_7\
        );

    \I__3254\ : InMux
    port map (
            O => \N__15959\,
            I => \N__15956\
        );

    \I__3253\ : LocalMux
    port map (
            O => \N__15956\,
            I => \b2v_inst.un2_indice_3_0_iv_0_a2_5_sx_2\
        );

    \I__3252\ : CascadeMux
    port map (
            O => \N__15953\,
            I => \b2v_inst.N_452_cascade_\
        );

    \I__3251\ : InMux
    port map (
            O => \N__15950\,
            I => \N__15947\
        );

    \I__3250\ : LocalMux
    port map (
            O => \N__15947\,
            I => \N__15942\
        );

    \I__3249\ : InMux
    port map (
            O => \N__15946\,
            I => \N__15937\
        );

    \I__3248\ : InMux
    port map (
            O => \N__15945\,
            I => \N__15937\
        );

    \I__3247\ : Span4Mux_h
    port map (
            O => \N__15942\,
            I => \N__15934\
        );

    \I__3246\ : LocalMux
    port map (
            O => \N__15937\,
            I => \N__15931\
        );

    \I__3245\ : Odrv4
    port map (
            O => \N__15934\,
            I => \b2v_inst.stateZ0Z_13\
        );

    \I__3244\ : Odrv4
    port map (
            O => \N__15931\,
            I => \b2v_inst.stateZ0Z_13\
        );

    \I__3243\ : InMux
    port map (
            O => \N__15926\,
            I => \N__15923\
        );

    \I__3242\ : LocalMux
    port map (
            O => \N__15923\,
            I => \N__15920\
        );

    \I__3241\ : Span4Mux_h
    port map (
            O => \N__15920\,
            I => \N__15917\
        );

    \I__3240\ : Odrv4
    port map (
            O => \N__15917\,
            I => \b2v_inst.g2_3\
        );

    \I__3239\ : InMux
    port map (
            O => \N__15914\,
            I => \N__15911\
        );

    \I__3238\ : LocalMux
    port map (
            O => \N__15911\,
            I => \N__15907\
        );

    \I__3237\ : InMux
    port map (
            O => \N__15910\,
            I => \N__15904\
        );

    \I__3236\ : Span4Mux_h
    port map (
            O => \N__15907\,
            I => \N__15896\
        );

    \I__3235\ : LocalMux
    port map (
            O => \N__15904\,
            I => \N__15896\
        );

    \I__3234\ : InMux
    port map (
            O => \N__15903\,
            I => \N__15893\
        );

    \I__3233\ : InMux
    port map (
            O => \N__15902\,
            I => \N__15890\
        );

    \I__3232\ : InMux
    port map (
            O => \N__15901\,
            I => \N__15887\
        );

    \I__3231\ : Span4Mux_h
    port map (
            O => \N__15896\,
            I => \N__15884\
        );

    \I__3230\ : LocalMux
    port map (
            O => \N__15893\,
            I => \N__15879\
        );

    \I__3229\ : LocalMux
    port map (
            O => \N__15890\,
            I => \N__15879\
        );

    \I__3228\ : LocalMux
    port map (
            O => \N__15887\,
            I => \b2v_inst.borradoZ0\
        );

    \I__3227\ : Odrv4
    port map (
            O => \N__15884\,
            I => \b2v_inst.borradoZ0\
        );

    \I__3226\ : Odrv12
    port map (
            O => \N__15879\,
            I => \b2v_inst.borradoZ0\
        );

    \I__3225\ : InMux
    port map (
            O => \N__15872\,
            I => \N__15868\
        );

    \I__3224\ : InMux
    port map (
            O => \N__15871\,
            I => \N__15862\
        );

    \I__3223\ : LocalMux
    port map (
            O => \N__15868\,
            I => \N__15859\
        );

    \I__3222\ : InMux
    port map (
            O => \N__15867\,
            I => \N__15854\
        );

    \I__3221\ : InMux
    port map (
            O => \N__15866\,
            I => \N__15854\
        );

    \I__3220\ : InMux
    port map (
            O => \N__15865\,
            I => \N__15851\
        );

    \I__3219\ : LocalMux
    port map (
            O => \N__15862\,
            I => \N__15848\
        );

    \I__3218\ : Span4Mux_h
    port map (
            O => \N__15859\,
            I => \N__15841\
        );

    \I__3217\ : LocalMux
    port map (
            O => \N__15854\,
            I => \N__15838\
        );

    \I__3216\ : LocalMux
    port map (
            O => \N__15851\,
            I => \N__15835\
        );

    \I__3215\ : Span4Mux_h
    port map (
            O => \N__15848\,
            I => \N__15832\
        );

    \I__3214\ : InMux
    port map (
            O => \N__15847\,
            I => \N__15829\
        );

    \I__3213\ : InMux
    port map (
            O => \N__15846\,
            I => \N__15822\
        );

    \I__3212\ : InMux
    port map (
            O => \N__15845\,
            I => \N__15822\
        );

    \I__3211\ : InMux
    port map (
            O => \N__15844\,
            I => \N__15822\
        );

    \I__3210\ : Odrv4
    port map (
            O => \N__15841\,
            I => \b2v_inst.stateZ0Z_5\
        );

    \I__3209\ : Odrv12
    port map (
            O => \N__15838\,
            I => \b2v_inst.stateZ0Z_5\
        );

    \I__3208\ : Odrv4
    port map (
            O => \N__15835\,
            I => \b2v_inst.stateZ0Z_5\
        );

    \I__3207\ : Odrv4
    port map (
            O => \N__15832\,
            I => \b2v_inst.stateZ0Z_5\
        );

    \I__3206\ : LocalMux
    port map (
            O => \N__15829\,
            I => \b2v_inst.stateZ0Z_5\
        );

    \I__3205\ : LocalMux
    port map (
            O => \N__15822\,
            I => \b2v_inst.stateZ0Z_5\
        );

    \I__3204\ : CascadeMux
    port map (
            O => \N__15809\,
            I => \b2v_inst.N_7_1_cascade_\
        );

    \I__3203\ : CascadeMux
    port map (
            O => \N__15806\,
            I => \b2v_inst.g2_2_cascade_\
        );

    \I__3202\ : InMux
    port map (
            O => \N__15803\,
            I => \N__15800\
        );

    \I__3201\ : LocalMux
    port map (
            O => \N__15800\,
            I => \b2v_inst.g1\
        );

    \I__3200\ : InMux
    port map (
            O => \N__15797\,
            I => \N__15794\
        );

    \I__3199\ : LocalMux
    port map (
            O => \N__15794\,
            I => \b2v_inst.un2_indice_21_s0_0_6\
        );

    \I__3198\ : CascadeMux
    port map (
            O => \N__15791\,
            I => \b2v_inst.N_253_cascade_\
        );

    \I__3197\ : InMux
    port map (
            O => \N__15788\,
            I => \N__15782\
        );

    \I__3196\ : InMux
    port map (
            O => \N__15787\,
            I => \N__15782\
        );

    \I__3195\ : LocalMux
    port map (
            O => \N__15782\,
            I => \N__15779\
        );

    \I__3194\ : Odrv4
    port map (
            O => \N__15779\,
            I => \b2v_inst.state_fastZ0Z_17\
        );

    \I__3193\ : InMux
    port map (
            O => \N__15776\,
            I => \N__15770\
        );

    \I__3192\ : InMux
    port map (
            O => \N__15775\,
            I => \N__15770\
        );

    \I__3191\ : LocalMux
    port map (
            O => \N__15770\,
            I => \N__15767\
        );

    \I__3190\ : Odrv4
    port map (
            O => \N__15767\,
            I => \b2v_inst.state_fastZ0Z_15\
        );

    \I__3189\ : CascadeMux
    port map (
            O => \N__15764\,
            I => \b2v_inst.N_253_i_cascade_\
        );

    \I__3188\ : InMux
    port map (
            O => \N__15761\,
            I => \N__15758\
        );

    \I__3187\ : LocalMux
    port map (
            O => \N__15758\,
            I => \N__15755\
        );

    \I__3186\ : Odrv4
    port map (
            O => \N__15755\,
            I => \b2v_inst.dir_mem_3_RNO_0Z0Z_3\
        );

    \I__3185\ : CascadeMux
    port map (
            O => \N__15752\,
            I => \b2v_inst1.r_RX_Bytece_0_0_1_cascade_\
        );

    \I__3184\ : InMux
    port map (
            O => \N__15749\,
            I => \N__15746\
        );

    \I__3183\ : LocalMux
    port map (
            O => \N__15746\,
            I => \N__15743\
        );

    \I__3182\ : Span4Mux_h
    port map (
            O => \N__15743\,
            I => \N__15739\
        );

    \I__3181\ : InMux
    port map (
            O => \N__15742\,
            I => \N__15736\
        );

    \I__3180\ : Odrv4
    port map (
            O => \N__15739\,
            I => \SYNTHESIZED_WIRE_10_1\
        );

    \I__3179\ : LocalMux
    port map (
            O => \N__15736\,
            I => \SYNTHESIZED_WIRE_10_1\
        );

    \I__3178\ : InMux
    port map (
            O => \N__15731\,
            I => \N__15728\
        );

    \I__3177\ : LocalMux
    port map (
            O => \N__15728\,
            I => \b2v_inst.dir_mem_2_RNO_0Z0Z_6\
        );

    \I__3176\ : InMux
    port map (
            O => \N__15725\,
            I => \N__15722\
        );

    \I__3175\ : LocalMux
    port map (
            O => \N__15722\,
            I => \N__15716\
        );

    \I__3174\ : InMux
    port map (
            O => \N__15721\,
            I => \N__15711\
        );

    \I__3173\ : InMux
    port map (
            O => \N__15720\,
            I => \N__15711\
        );

    \I__3172\ : CascadeMux
    port map (
            O => \N__15719\,
            I => \N__15708\
        );

    \I__3171\ : Span4Mux_h
    port map (
            O => \N__15716\,
            I => \N__15705\
        );

    \I__3170\ : LocalMux
    port map (
            O => \N__15711\,
            I => \N__15702\
        );

    \I__3169\ : InMux
    port map (
            O => \N__15708\,
            I => \N__15699\
        );

    \I__3168\ : Span4Mux_v
    port map (
            O => \N__15705\,
            I => \N__15696\
        );

    \I__3167\ : Span12Mux_v
    port map (
            O => \N__15702\,
            I => \N__15693\
        );

    \I__3166\ : LocalMux
    port map (
            O => \N__15699\,
            I => \SYNTHESIZED_WIRE_9\
        );

    \I__3165\ : Odrv4
    port map (
            O => \N__15696\,
            I => \SYNTHESIZED_WIRE_9\
        );

    \I__3164\ : Odrv12
    port map (
            O => \N__15693\,
            I => \SYNTHESIZED_WIRE_9\
        );

    \I__3163\ : CascadeMux
    port map (
            O => \N__15686\,
            I => \N__15674\
        );

    \I__3162\ : CascadeMux
    port map (
            O => \N__15685\,
            I => \N__15671\
        );

    \I__3161\ : InMux
    port map (
            O => \N__15684\,
            I => \N__15668\
        );

    \I__3160\ : InMux
    port map (
            O => \N__15683\,
            I => \N__15665\
        );

    \I__3159\ : InMux
    port map (
            O => \N__15682\,
            I => \N__15660\
        );

    \I__3158\ : InMux
    port map (
            O => \N__15681\,
            I => \N__15660\
        );

    \I__3157\ : InMux
    port map (
            O => \N__15680\,
            I => \N__15655\
        );

    \I__3156\ : InMux
    port map (
            O => \N__15679\,
            I => \N__15655\
        );

    \I__3155\ : InMux
    port map (
            O => \N__15678\,
            I => \N__15652\
        );

    \I__3154\ : InMux
    port map (
            O => \N__15677\,
            I => \N__15645\
        );

    \I__3153\ : InMux
    port map (
            O => \N__15674\,
            I => \N__15645\
        );

    \I__3152\ : InMux
    port map (
            O => \N__15671\,
            I => \N__15645\
        );

    \I__3151\ : LocalMux
    port map (
            O => \N__15668\,
            I => \N__15642\
        );

    \I__3150\ : LocalMux
    port map (
            O => \N__15665\,
            I => \N__15639\
        );

    \I__3149\ : LocalMux
    port map (
            O => \N__15660\,
            I => \N__15634\
        );

    \I__3148\ : LocalMux
    port map (
            O => \N__15655\,
            I => \N__15634\
        );

    \I__3147\ : LocalMux
    port map (
            O => \N__15652\,
            I => \N__15629\
        );

    \I__3146\ : LocalMux
    port map (
            O => \N__15645\,
            I => \N__15626\
        );

    \I__3145\ : Span12Mux_h
    port map (
            O => \N__15642\,
            I => \N__15621\
        );

    \I__3144\ : Span12Mux_s8_h
    port map (
            O => \N__15639\,
            I => \N__15621\
        );

    \I__3143\ : Span4Mux_h
    port map (
            O => \N__15634\,
            I => \N__15618\
        );

    \I__3142\ : InMux
    port map (
            O => \N__15633\,
            I => \N__15613\
        );

    \I__3141\ : InMux
    port map (
            O => \N__15632\,
            I => \N__15613\
        );

    \I__3140\ : Span4Mux_v
    port map (
            O => \N__15629\,
            I => \N__15608\
        );

    \I__3139\ : Span4Mux_v
    port map (
            O => \N__15626\,
            I => \N__15608\
        );

    \I__3138\ : Odrv12
    port map (
            O => \N__15621\,
            I => \b2v_inst.stateZ0Z_16\
        );

    \I__3137\ : Odrv4
    port map (
            O => \N__15618\,
            I => \b2v_inst.stateZ0Z_16\
        );

    \I__3136\ : LocalMux
    port map (
            O => \N__15613\,
            I => \b2v_inst.stateZ0Z_16\
        );

    \I__3135\ : Odrv4
    port map (
            O => \N__15608\,
            I => \b2v_inst.stateZ0Z_16\
        );

    \I__3134\ : InMux
    port map (
            O => \N__15599\,
            I => \N__15581\
        );

    \I__3133\ : InMux
    port map (
            O => \N__15598\,
            I => \N__15581\
        );

    \I__3132\ : InMux
    port map (
            O => \N__15597\,
            I => \N__15581\
        );

    \I__3131\ : InMux
    port map (
            O => \N__15596\,
            I => \N__15581\
        );

    \I__3130\ : InMux
    port map (
            O => \N__15595\,
            I => \N__15581\
        );

    \I__3129\ : InMux
    port map (
            O => \N__15594\,
            I => \N__15581\
        );

    \I__3128\ : LocalMux
    port map (
            O => \N__15581\,
            I => \N__15578\
        );

    \I__3127\ : Span4Mux_v
    port map (
            O => \N__15578\,
            I => \N__15572\
        );

    \I__3126\ : InMux
    port map (
            O => \N__15577\,
            I => \N__15567\
        );

    \I__3125\ : InMux
    port map (
            O => \N__15576\,
            I => \N__15567\
        );

    \I__3124\ : CascadeMux
    port map (
            O => \N__15575\,
            I => \N__15560\
        );

    \I__3123\ : Span4Mux_v
    port map (
            O => \N__15572\,
            I => \N__15554\
        );

    \I__3122\ : LocalMux
    port map (
            O => \N__15567\,
            I => \N__15554\
        );

    \I__3121\ : InMux
    port map (
            O => \N__15566\,
            I => \N__15541\
        );

    \I__3120\ : InMux
    port map (
            O => \N__15565\,
            I => \N__15541\
        );

    \I__3119\ : InMux
    port map (
            O => \N__15564\,
            I => \N__15541\
        );

    \I__3118\ : InMux
    port map (
            O => \N__15563\,
            I => \N__15541\
        );

    \I__3117\ : InMux
    port map (
            O => \N__15560\,
            I => \N__15541\
        );

    \I__3116\ : InMux
    port map (
            O => \N__15559\,
            I => \N__15541\
        );

    \I__3115\ : Span4Mux_h
    port map (
            O => \N__15554\,
            I => \N__15536\
        );

    \I__3114\ : LocalMux
    port map (
            O => \N__15541\,
            I => \N__15536\
        );

    \I__3113\ : Span4Mux_v
    port map (
            O => \N__15536\,
            I => \N__15531\
        );

    \I__3112\ : InMux
    port map (
            O => \N__15535\,
            I => \N__15526\
        );

    \I__3111\ : InMux
    port map (
            O => \N__15534\,
            I => \N__15526\
        );

    \I__3110\ : Odrv4
    port map (
            O => \N__15531\,
            I => \b2v_inst.ignorar_anteriorZ0\
        );

    \I__3109\ : LocalMux
    port map (
            O => \N__15526\,
            I => \b2v_inst.ignorar_anteriorZ0\
        );

    \I__3108\ : CEMux
    port map (
            O => \N__15521\,
            I => \N__15518\
        );

    \I__3107\ : LocalMux
    port map (
            O => \N__15518\,
            I => \N__15515\
        );

    \I__3106\ : Span4Mux_h
    port map (
            O => \N__15515\,
            I => \N__15512\
        );

    \I__3105\ : Span4Mux_h
    port map (
            O => \N__15512\,
            I => \N__15509\
        );

    \I__3104\ : Odrv4
    port map (
            O => \N__15509\,
            I => \b2v_inst.un1_state_19_0\
        );

    \I__3103\ : CascadeMux
    port map (
            O => \N__15506\,
            I => \N__15503\
        );

    \I__3102\ : InMux
    port map (
            O => \N__15503\,
            I => \N__15500\
        );

    \I__3101\ : LocalMux
    port map (
            O => \N__15500\,
            I => \N__15497\
        );

    \I__3100\ : Span4Mux_v
    port map (
            O => \N__15497\,
            I => \N__15494\
        );

    \I__3099\ : Odrv4
    port map (
            O => \N__15494\,
            I => \b2v_inst.N_5\
        );

    \I__3098\ : CEMux
    port map (
            O => \N__15491\,
            I => \N__15487\
        );

    \I__3097\ : CEMux
    port map (
            O => \N__15490\,
            I => \N__15484\
        );

    \I__3096\ : LocalMux
    port map (
            O => \N__15487\,
            I => \N__15481\
        );

    \I__3095\ : LocalMux
    port map (
            O => \N__15484\,
            I => \N__15478\
        );

    \I__3094\ : Span4Mux_h
    port map (
            O => \N__15481\,
            I => \N__15474\
        );

    \I__3093\ : Span4Mux_h
    port map (
            O => \N__15478\,
            I => \N__15471\
        );

    \I__3092\ : InMux
    port map (
            O => \N__15477\,
            I => \N__15466\
        );

    \I__3091\ : Span4Mux_v
    port map (
            O => \N__15474\,
            I => \N__15463\
        );

    \I__3090\ : Span4Mux_h
    port map (
            O => \N__15471\,
            I => \N__15460\
        );

    \I__3089\ : InMux
    port map (
            O => \N__15470\,
            I => \N__15457\
        );

    \I__3088\ : InMux
    port map (
            O => \N__15469\,
            I => \N__15454\
        );

    \I__3087\ : LocalMux
    port map (
            O => \N__15466\,
            I => \N__15451\
        );

    \I__3086\ : Odrv4
    port map (
            O => \N__15463\,
            I => \b2v_inst.stateZ0Z_10\
        );

    \I__3085\ : Odrv4
    port map (
            O => \N__15460\,
            I => \b2v_inst.stateZ0Z_10\
        );

    \I__3084\ : LocalMux
    port map (
            O => \N__15457\,
            I => \b2v_inst.stateZ0Z_10\
        );

    \I__3083\ : LocalMux
    port map (
            O => \N__15454\,
            I => \b2v_inst.stateZ0Z_10\
        );

    \I__3082\ : Odrv4
    port map (
            O => \N__15451\,
            I => \b2v_inst.stateZ0Z_10\
        );

    \I__3081\ : InMux
    port map (
            O => \N__15440\,
            I => \N__15434\
        );

    \I__3080\ : InMux
    port map (
            O => \N__15439\,
            I => \N__15434\
        );

    \I__3079\ : LocalMux
    port map (
            O => \N__15434\,
            I => \b2v_inst.stateZ0Z_1\
        );

    \I__3078\ : CascadeMux
    port map (
            O => \N__15431\,
            I => \N__15428\
        );

    \I__3077\ : InMux
    port map (
            O => \N__15428\,
            I => \N__15425\
        );

    \I__3076\ : LocalMux
    port map (
            O => \N__15425\,
            I => \N__15422\
        );

    \I__3075\ : Odrv4
    port map (
            O => \N__15422\,
            I => \b2v_inst.dir_mem_3Z0Z_4\
        );

    \I__3074\ : CascadeMux
    port map (
            O => \N__15419\,
            I => \b2v_inst.addr_ram_1_0_iv_i_1_4_cascade_\
        );

    \I__3073\ : CascadeMux
    port map (
            O => \N__15416\,
            I => \N__15413\
        );

    \I__3072\ : InMux
    port map (
            O => \N__15413\,
            I => \N__15409\
        );

    \I__3071\ : CascadeMux
    port map (
            O => \N__15412\,
            I => \N__15406\
        );

    \I__3070\ : LocalMux
    port map (
            O => \N__15409\,
            I => \N__15403\
        );

    \I__3069\ : InMux
    port map (
            O => \N__15406\,
            I => \N__15400\
        );

    \I__3068\ : Span4Mux_v
    port map (
            O => \N__15403\,
            I => \N__15395\
        );

    \I__3067\ : LocalMux
    port map (
            O => \N__15400\,
            I => \N__15395\
        );

    \I__3066\ : Span4Mux_h
    port map (
            O => \N__15395\,
            I => \N__15392\
        );

    \I__3065\ : Odrv4
    port map (
            O => \N__15392\,
            I => \N_163\
        );

    \I__3064\ : CascadeMux
    port map (
            O => \N__15389\,
            I => \b2v_inst.g0_11_1_cascade_\
        );

    \I__3063\ : InMux
    port map (
            O => \N__15386\,
            I => \N__15383\
        );

    \I__3062\ : LocalMux
    port map (
            O => \N__15383\,
            I => \b2v_inst.dir_mem_1Z0Z_4\
        );

    \I__3061\ : InMux
    port map (
            O => \N__15380\,
            I => \N__15377\
        );

    \I__3060\ : LocalMux
    port map (
            O => \N__15377\,
            I => \N__15366\
        );

    \I__3059\ : InMux
    port map (
            O => \N__15376\,
            I => \N__15363\
        );

    \I__3058\ : InMux
    port map (
            O => \N__15375\,
            I => \N__15360\
        );

    \I__3057\ : InMux
    port map (
            O => \N__15374\,
            I => \N__15357\
        );

    \I__3056\ : InMux
    port map (
            O => \N__15373\,
            I => \N__15350\
        );

    \I__3055\ : InMux
    port map (
            O => \N__15372\,
            I => \N__15350\
        );

    \I__3054\ : InMux
    port map (
            O => \N__15371\,
            I => \N__15350\
        );

    \I__3053\ : InMux
    port map (
            O => \N__15370\,
            I => \N__15345\
        );

    \I__3052\ : InMux
    port map (
            O => \N__15369\,
            I => \N__15345\
        );

    \I__3051\ : Odrv4
    port map (
            O => \N__15366\,
            I => \b2v_inst.N_235\
        );

    \I__3050\ : LocalMux
    port map (
            O => \N__15363\,
            I => \b2v_inst.N_235\
        );

    \I__3049\ : LocalMux
    port map (
            O => \N__15360\,
            I => \b2v_inst.N_235\
        );

    \I__3048\ : LocalMux
    port map (
            O => \N__15357\,
            I => \b2v_inst.N_235\
        );

    \I__3047\ : LocalMux
    port map (
            O => \N__15350\,
            I => \b2v_inst.N_235\
        );

    \I__3046\ : LocalMux
    port map (
            O => \N__15345\,
            I => \b2v_inst.N_235\
        );

    \I__3045\ : InMux
    port map (
            O => \N__15332\,
            I => \N__15329\
        );

    \I__3044\ : LocalMux
    port map (
            O => \N__15329\,
            I => \b2v_inst.addr_ram_1_0_iv_i_0_4\
        );

    \I__3043\ : CascadeMux
    port map (
            O => \N__15326\,
            I => \N__15321\
        );

    \I__3042\ : CascadeMux
    port map (
            O => \N__15325\,
            I => \N__15318\
        );

    \I__3041\ : InMux
    port map (
            O => \N__15324\,
            I => \N__15312\
        );

    \I__3040\ : InMux
    port map (
            O => \N__15321\,
            I => \N__15301\
        );

    \I__3039\ : InMux
    port map (
            O => \N__15318\,
            I => \N__15301\
        );

    \I__3038\ : InMux
    port map (
            O => \N__15317\,
            I => \N__15301\
        );

    \I__3037\ : InMux
    port map (
            O => \N__15316\,
            I => \N__15301\
        );

    \I__3036\ : InMux
    port map (
            O => \N__15315\,
            I => \N__15301\
        );

    \I__3035\ : LocalMux
    port map (
            O => \N__15312\,
            I => \b2v_inst.dir_mem_315_0\
        );

    \I__3034\ : LocalMux
    port map (
            O => \N__15301\,
            I => \b2v_inst.dir_mem_315_0\
        );

    \I__3033\ : InMux
    port map (
            O => \N__15296\,
            I => \N__15293\
        );

    \I__3032\ : LocalMux
    port map (
            O => \N__15293\,
            I => \N__15290\
        );

    \I__3031\ : Odrv4
    port map (
            O => \N__15290\,
            I => \b2v_inst.dir_mem_3Z0Z_3\
        );

    \I__3030\ : InMux
    port map (
            O => \N__15287\,
            I => \N__15284\
        );

    \I__3029\ : LocalMux
    port map (
            O => \N__15284\,
            I => \N__15281\
        );

    \I__3028\ : Span4Mux_h
    port map (
            O => \N__15281\,
            I => \N__15278\
        );

    \I__3027\ : Odrv4
    port map (
            O => \N__15278\,
            I => \b2v_inst.dir_mem_3Z0Z_7\
        );

    \I__3026\ : CEMux
    port map (
            O => \N__15275\,
            I => \N__15271\
        );

    \I__3025\ : CEMux
    port map (
            O => \N__15274\,
            I => \N__15268\
        );

    \I__3024\ : LocalMux
    port map (
            O => \N__15271\,
            I => \N__15263\
        );

    \I__3023\ : LocalMux
    port map (
            O => \N__15268\,
            I => \N__15263\
        );

    \I__3022\ : Span4Mux_v
    port map (
            O => \N__15263\,
            I => \N__15260\
        );

    \I__3021\ : Span4Mux_v
    port map (
            O => \N__15260\,
            I => \N__15257\
        );

    \I__3020\ : Sp12to4
    port map (
            O => \N__15257\,
            I => \N__15254\
        );

    \I__3019\ : Odrv12
    port map (
            O => \N__15254\,
            I => \b2v_inst.N_138_i\
        );

    \I__3018\ : InMux
    port map (
            O => \N__15251\,
            I => \N__15248\
        );

    \I__3017\ : LocalMux
    port map (
            O => \N__15248\,
            I => \N__15245\
        );

    \I__3016\ : Span4Mux_v
    port map (
            O => \N__15245\,
            I => \N__15242\
        );

    \I__3015\ : Odrv4
    port map (
            O => \N__15242\,
            I => \b2v_inst1.r_RX_Bytece_0_5\
        );

    \I__3014\ : CEMux
    port map (
            O => \N__15239\,
            I => \N__15236\
        );

    \I__3013\ : LocalMux
    port map (
            O => \N__15236\,
            I => \N__15231\
        );

    \I__3012\ : CEMux
    port map (
            O => \N__15235\,
            I => \N__15228\
        );

    \I__3011\ : InMux
    port map (
            O => \N__15234\,
            I => \N__15225\
        );

    \I__3010\ : Span4Mux_h
    port map (
            O => \N__15231\,
            I => \N__15219\
        );

    \I__3009\ : LocalMux
    port map (
            O => \N__15228\,
            I => \N__15219\
        );

    \I__3008\ : LocalMux
    port map (
            O => \N__15225\,
            I => \N__15216\
        );

    \I__3007\ : CascadeMux
    port map (
            O => \N__15224\,
            I => \N__15210\
        );

    \I__3006\ : Span4Mux_v
    port map (
            O => \N__15219\,
            I => \N__15207\
        );

    \I__3005\ : Span4Mux_h
    port map (
            O => \N__15216\,
            I => \N__15204\
        );

    \I__3004\ : InMux
    port map (
            O => \N__15215\,
            I => \N__15197\
        );

    \I__3003\ : InMux
    port map (
            O => \N__15214\,
            I => \N__15197\
        );

    \I__3002\ : InMux
    port map (
            O => \N__15213\,
            I => \N__15197\
        );

    \I__3001\ : InMux
    port map (
            O => \N__15210\,
            I => \N__15194\
        );

    \I__3000\ : Odrv4
    port map (
            O => \N__15207\,
            I => \b2v_inst.stateZ0Z_14\
        );

    \I__2999\ : Odrv4
    port map (
            O => \N__15204\,
            I => \b2v_inst.stateZ0Z_14\
        );

    \I__2998\ : LocalMux
    port map (
            O => \N__15197\,
            I => \b2v_inst.stateZ0Z_14\
        );

    \I__2997\ : LocalMux
    port map (
            O => \N__15194\,
            I => \b2v_inst.stateZ0Z_14\
        );

    \I__2996\ : InMux
    port map (
            O => \N__15185\,
            I => \N__15177\
        );

    \I__2995\ : InMux
    port map (
            O => \N__15184\,
            I => \N__15174\
        );

    \I__2994\ : InMux
    port map (
            O => \N__15183\,
            I => \N__15165\
        );

    \I__2993\ : InMux
    port map (
            O => \N__15182\,
            I => \N__15165\
        );

    \I__2992\ : InMux
    port map (
            O => \N__15181\,
            I => \N__15165\
        );

    \I__2991\ : InMux
    port map (
            O => \N__15180\,
            I => \N__15165\
        );

    \I__2990\ : LocalMux
    port map (
            O => \N__15177\,
            I => \N__15162\
        );

    \I__2989\ : LocalMux
    port map (
            O => \N__15174\,
            I => \N__15157\
        );

    \I__2988\ : LocalMux
    port map (
            O => \N__15165\,
            I => \N__15157\
        );

    \I__2987\ : Span12Mux_h
    port map (
            O => \N__15162\,
            I => \N__15154\
        );

    \I__2986\ : Span4Mux_v
    port map (
            O => \N__15157\,
            I => \N__15151\
        );

    \I__2985\ : Odrv12
    port map (
            O => \N__15154\,
            I => \b2v_inst.stateZ0Z_6\
        );

    \I__2984\ : Odrv4
    port map (
            O => \N__15151\,
            I => \b2v_inst.stateZ0Z_6\
        );

    \I__2983\ : InMux
    port map (
            O => \N__15146\,
            I => \N__15140\
        );

    \I__2982\ : InMux
    port map (
            O => \N__15145\,
            I => \N__15140\
        );

    \I__2981\ : LocalMux
    port map (
            O => \N__15140\,
            I => \N__15135\
        );

    \I__2980\ : InMux
    port map (
            O => \N__15139\,
            I => \N__15132\
        );

    \I__2979\ : InMux
    port map (
            O => \N__15138\,
            I => \N__15129\
        );

    \I__2978\ : Span4Mux_v
    port map (
            O => \N__15135\,
            I => \N__15126\
        );

    \I__2977\ : LocalMux
    port map (
            O => \N__15132\,
            I => \b2v_inst.state_RNITETBZ0Z_0\
        );

    \I__2976\ : LocalMux
    port map (
            O => \N__15129\,
            I => \b2v_inst.state_RNITETBZ0Z_0\
        );

    \I__2975\ : Odrv4
    port map (
            O => \N__15126\,
            I => \b2v_inst.state_RNITETBZ0Z_0\
        );

    \I__2974\ : CascadeMux
    port map (
            O => \N__15119\,
            I => \b2v_inst.N_351_cascade_\
        );

    \I__2973\ : InMux
    port map (
            O => \N__15116\,
            I => \N__15113\
        );

    \I__2972\ : LocalMux
    port map (
            O => \N__15113\,
            I => \b2v_inst.addr_ram_1_iv_i_1_3\
        );

    \I__2971\ : CascadeMux
    port map (
            O => \N__15110\,
            I => \b2v_inst.addr_ram_1_iv_i_2_3_cascade_\
        );

    \I__2970\ : CascadeMux
    port map (
            O => \N__15107\,
            I => \N__15104\
        );

    \I__2969\ : InMux
    port map (
            O => \N__15104\,
            I => \N__15100\
        );

    \I__2968\ : CascadeMux
    port map (
            O => \N__15103\,
            I => \N__15097\
        );

    \I__2967\ : LocalMux
    port map (
            O => \N__15100\,
            I => \N__15094\
        );

    \I__2966\ : InMux
    port map (
            O => \N__15097\,
            I => \N__15091\
        );

    \I__2965\ : Span4Mux_v
    port map (
            O => \N__15094\,
            I => \N__15086\
        );

    \I__2964\ : LocalMux
    port map (
            O => \N__15091\,
            I => \N__15086\
        );

    \I__2963\ : Span4Mux_h
    port map (
            O => \N__15086\,
            I => \N__15083\
        );

    \I__2962\ : Odrv4
    port map (
            O => \N__15083\,
            I => \N_58\
        );

    \I__2961\ : InMux
    port map (
            O => \N__15080\,
            I => \N__15077\
        );

    \I__2960\ : LocalMux
    port map (
            O => \N__15077\,
            I => \N__15074\
        );

    \I__2959\ : Span4Mux_v
    port map (
            O => \N__15074\,
            I => \N__15070\
        );

    \I__2958\ : InMux
    port map (
            O => \N__15073\,
            I => \N__15067\
        );

    \I__2957\ : Odrv4
    port map (
            O => \N__15070\,
            I => \b2v_inst.stateZ0Z_0\
        );

    \I__2956\ : LocalMux
    port map (
            O => \N__15067\,
            I => \b2v_inst.stateZ0Z_0\
        );

    \I__2955\ : CascadeMux
    port map (
            O => \N__15062\,
            I => \N__15055\
        );

    \I__2954\ : InMux
    port map (
            O => \N__15061\,
            I => \N__15046\
        );

    \I__2953\ : InMux
    port map (
            O => \N__15060\,
            I => \N__15046\
        );

    \I__2952\ : InMux
    port map (
            O => \N__15059\,
            I => \N__15046\
        );

    \I__2951\ : InMux
    port map (
            O => \N__15058\,
            I => \N__15043\
        );

    \I__2950\ : InMux
    port map (
            O => \N__15055\,
            I => \N__15036\
        );

    \I__2949\ : InMux
    port map (
            O => \N__15054\,
            I => \N__15036\
        );

    \I__2948\ : InMux
    port map (
            O => \N__15053\,
            I => \N__15036\
        );

    \I__2947\ : LocalMux
    port map (
            O => \N__15046\,
            I => \b2v_inst.cuentaZ0Z_5\
        );

    \I__2946\ : LocalMux
    port map (
            O => \N__15043\,
            I => \b2v_inst.cuentaZ0Z_5\
        );

    \I__2945\ : LocalMux
    port map (
            O => \N__15036\,
            I => \b2v_inst.cuentaZ0Z_5\
        );

    \I__2944\ : CascadeMux
    port map (
            O => \N__15029\,
            I => \N__15023\
        );

    \I__2943\ : InMux
    port map (
            O => \N__15028\,
            I => \N__15017\
        );

    \I__2942\ : InMux
    port map (
            O => \N__15027\,
            I => \N__15008\
        );

    \I__2941\ : InMux
    port map (
            O => \N__15026\,
            I => \N__15008\
        );

    \I__2940\ : InMux
    port map (
            O => \N__15023\,
            I => \N__15008\
        );

    \I__2939\ : InMux
    port map (
            O => \N__15022\,
            I => \N__15008\
        );

    \I__2938\ : InMux
    port map (
            O => \N__15021\,
            I => \N__15003\
        );

    \I__2937\ : InMux
    port map (
            O => \N__15020\,
            I => \N__15003\
        );

    \I__2936\ : LocalMux
    port map (
            O => \N__15017\,
            I => \N__14998\
        );

    \I__2935\ : LocalMux
    port map (
            O => \N__15008\,
            I => \N__14998\
        );

    \I__2934\ : LocalMux
    port map (
            O => \N__15003\,
            I => \b2v_inst.cuentaZ0Z_4\
        );

    \I__2933\ : Odrv4
    port map (
            O => \N__14998\,
            I => \b2v_inst.cuentaZ0Z_4\
        );

    \I__2932\ : CascadeMux
    port map (
            O => \N__14993\,
            I => \b2v_inst.un4_cuenta_ac0_9_0_cascade_\
        );

    \I__2931\ : InMux
    port map (
            O => \N__14990\,
            I => \N__14981\
        );

    \I__2930\ : InMux
    port map (
            O => \N__14989\,
            I => \N__14978\
        );

    \I__2929\ : InMux
    port map (
            O => \N__14988\,
            I => \N__14975\
        );

    \I__2928\ : InMux
    port map (
            O => \N__14987\,
            I => \N__14966\
        );

    \I__2927\ : InMux
    port map (
            O => \N__14986\,
            I => \N__14966\
        );

    \I__2926\ : InMux
    port map (
            O => \N__14985\,
            I => \N__14966\
        );

    \I__2925\ : InMux
    port map (
            O => \N__14984\,
            I => \N__14966\
        );

    \I__2924\ : LocalMux
    port map (
            O => \N__14981\,
            I => \b2v_inst.un4_cuenta_c4\
        );

    \I__2923\ : LocalMux
    port map (
            O => \N__14978\,
            I => \b2v_inst.un4_cuenta_c4\
        );

    \I__2922\ : LocalMux
    port map (
            O => \N__14975\,
            I => \b2v_inst.un4_cuenta_c4\
        );

    \I__2921\ : LocalMux
    port map (
            O => \N__14966\,
            I => \b2v_inst.un4_cuenta_c4\
        );

    \I__2920\ : InMux
    port map (
            O => \N__14957\,
            I => \N__14949\
        );

    \I__2919\ : InMux
    port map (
            O => \N__14956\,
            I => \N__14942\
        );

    \I__2918\ : InMux
    port map (
            O => \N__14955\,
            I => \N__14942\
        );

    \I__2917\ : InMux
    port map (
            O => \N__14954\,
            I => \N__14942\
        );

    \I__2916\ : InMux
    port map (
            O => \N__14953\,
            I => \N__14939\
        );

    \I__2915\ : InMux
    port map (
            O => \N__14952\,
            I => \N__14936\
        );

    \I__2914\ : LocalMux
    port map (
            O => \N__14949\,
            I => \b2v_inst.cuentaZ0Z_6\
        );

    \I__2913\ : LocalMux
    port map (
            O => \N__14942\,
            I => \b2v_inst.cuentaZ0Z_6\
        );

    \I__2912\ : LocalMux
    port map (
            O => \N__14939\,
            I => \b2v_inst.cuentaZ0Z_6\
        );

    \I__2911\ : LocalMux
    port map (
            O => \N__14936\,
            I => \b2v_inst.cuentaZ0Z_6\
        );

    \I__2910\ : InMux
    port map (
            O => \N__14927\,
            I => \N__14919\
        );

    \I__2909\ : InMux
    port map (
            O => \N__14926\,
            I => \N__14919\
        );

    \I__2908\ : InMux
    port map (
            O => \N__14925\,
            I => \N__14916\
        );

    \I__2907\ : InMux
    port map (
            O => \N__14924\,
            I => \N__14913\
        );

    \I__2906\ : LocalMux
    port map (
            O => \N__14919\,
            I => \b2v_inst.cuentaZ0Z_7\
        );

    \I__2905\ : LocalMux
    port map (
            O => \N__14916\,
            I => \b2v_inst.cuentaZ0Z_7\
        );

    \I__2904\ : LocalMux
    port map (
            O => \N__14913\,
            I => \b2v_inst.cuentaZ0Z_7\
        );

    \I__2903\ : CEMux
    port map (
            O => \N__14906\,
            I => \N__14902\
        );

    \I__2902\ : CEMux
    port map (
            O => \N__14905\,
            I => \N__14899\
        );

    \I__2901\ : LocalMux
    port map (
            O => \N__14902\,
            I => \N__14892\
        );

    \I__2900\ : LocalMux
    port map (
            O => \N__14899\,
            I => \N__14892\
        );

    \I__2899\ : CEMux
    port map (
            O => \N__14898\,
            I => \N__14889\
        );

    \I__2898\ : CEMux
    port map (
            O => \N__14897\,
            I => \N__14886\
        );

    \I__2897\ : Span4Mux_v
    port map (
            O => \N__14892\,
            I => \N__14883\
        );

    \I__2896\ : LocalMux
    port map (
            O => \N__14889\,
            I => \N__14880\
        );

    \I__2895\ : LocalMux
    port map (
            O => \N__14886\,
            I => \b2v_inst.N_399_i\
        );

    \I__2894\ : Odrv4
    port map (
            O => \N__14883\,
            I => \b2v_inst.N_399_i\
        );

    \I__2893\ : Odrv4
    port map (
            O => \N__14880\,
            I => \b2v_inst.N_399_i\
        );

    \I__2892\ : InMux
    port map (
            O => \N__14873\,
            I => \N__14869\
        );

    \I__2891\ : InMux
    port map (
            O => \N__14872\,
            I => \N__14866\
        );

    \I__2890\ : LocalMux
    port map (
            O => \N__14869\,
            I => \N__14863\
        );

    \I__2889\ : LocalMux
    port map (
            O => \N__14866\,
            I => \N__14860\
        );

    \I__2888\ : Span4Mux_h
    port map (
            O => \N__14863\,
            I => \N__14853\
        );

    \I__2887\ : Span4Mux_v
    port map (
            O => \N__14860\,
            I => \N__14850\
        );

    \I__2886\ : InMux
    port map (
            O => \N__14859\,
            I => \N__14847\
        );

    \I__2885\ : InMux
    port map (
            O => \N__14858\,
            I => \N__14844\
        );

    \I__2884\ : InMux
    port map (
            O => \N__14857\,
            I => \N__14839\
        );

    \I__2883\ : InMux
    port map (
            O => \N__14856\,
            I => \N__14839\
        );

    \I__2882\ : Span4Mux_h
    port map (
            O => \N__14853\,
            I => \N__14834\
        );

    \I__2881\ : Span4Mux_h
    port map (
            O => \N__14850\,
            I => \N__14834\
        );

    \I__2880\ : LocalMux
    port map (
            O => \N__14847\,
            I => \b2v_inst.N_227\
        );

    \I__2879\ : LocalMux
    port map (
            O => \N__14844\,
            I => \b2v_inst.N_227\
        );

    \I__2878\ : LocalMux
    port map (
            O => \N__14839\,
            I => \b2v_inst.N_227\
        );

    \I__2877\ : Odrv4
    port map (
            O => \N__14834\,
            I => \b2v_inst.N_227\
        );

    \I__2876\ : InMux
    port map (
            O => \N__14825\,
            I => \N__14821\
        );

    \I__2875\ : InMux
    port map (
            O => \N__14824\,
            I => \N__14817\
        );

    \I__2874\ : LocalMux
    port map (
            O => \N__14821\,
            I => \N__14814\
        );

    \I__2873\ : InMux
    port map (
            O => \N__14820\,
            I => \N__14811\
        );

    \I__2872\ : LocalMux
    port map (
            O => \N__14817\,
            I => \N__14808\
        );

    \I__2871\ : Odrv4
    port map (
            O => \N__14814\,
            I => \b2v_inst.N_232\
        );

    \I__2870\ : LocalMux
    port map (
            O => \N__14811\,
            I => \b2v_inst.N_232\
        );

    \I__2869\ : Odrv12
    port map (
            O => \N__14808\,
            I => \b2v_inst.N_232\
        );

    \I__2868\ : CascadeMux
    port map (
            O => \N__14801\,
            I => \b2v_inst.N_232_cascade_\
        );

    \I__2867\ : InMux
    port map (
            O => \N__14798\,
            I => \N__14788\
        );

    \I__2866\ : InMux
    port map (
            O => \N__14797\,
            I => \N__14782\
        );

    \I__2865\ : CascadeMux
    port map (
            O => \N__14796\,
            I => \N__14778\
        );

    \I__2864\ : InMux
    port map (
            O => \N__14795\,
            I => \N__14769\
        );

    \I__2863\ : InMux
    port map (
            O => \N__14794\,
            I => \N__14769\
        );

    \I__2862\ : InMux
    port map (
            O => \N__14793\,
            I => \N__14769\
        );

    \I__2861\ : InMux
    port map (
            O => \N__14792\,
            I => \N__14769\
        );

    \I__2860\ : InMux
    port map (
            O => \N__14791\,
            I => \N__14766\
        );

    \I__2859\ : LocalMux
    port map (
            O => \N__14788\,
            I => \N__14763\
        );

    \I__2858\ : InMux
    port map (
            O => \N__14787\,
            I => \N__14756\
        );

    \I__2857\ : InMux
    port map (
            O => \N__14786\,
            I => \N__14756\
        );

    \I__2856\ : InMux
    port map (
            O => \N__14785\,
            I => \N__14756\
        );

    \I__2855\ : LocalMux
    port map (
            O => \N__14782\,
            I => \N__14753\
        );

    \I__2854\ : InMux
    port map (
            O => \N__14781\,
            I => \N__14750\
        );

    \I__2853\ : InMux
    port map (
            O => \N__14778\,
            I => \N__14747\
        );

    \I__2852\ : LocalMux
    port map (
            O => \N__14769\,
            I => \N__14744\
        );

    \I__2851\ : LocalMux
    port map (
            O => \N__14766\,
            I => \N__14741\
        );

    \I__2850\ : Span4Mux_v
    port map (
            O => \N__14763\,
            I => \N__14736\
        );

    \I__2849\ : LocalMux
    port map (
            O => \N__14756\,
            I => \N__14736\
        );

    \I__2848\ : Span4Mux_v
    port map (
            O => \N__14753\,
            I => \N__14731\
        );

    \I__2847\ : LocalMux
    port map (
            O => \N__14750\,
            I => \N__14731\
        );

    \I__2846\ : LocalMux
    port map (
            O => \N__14747\,
            I => \N__14728\
        );

    \I__2845\ : Span4Mux_v
    port map (
            O => \N__14744\,
            I => \N__14725\
        );

    \I__2844\ : Span4Mux_v
    port map (
            O => \N__14741\,
            I => \N__14718\
        );

    \I__2843\ : Span4Mux_v
    port map (
            O => \N__14736\,
            I => \N__14718\
        );

    \I__2842\ : Span4Mux_v
    port map (
            O => \N__14731\,
            I => \N__14718\
        );

    \I__2841\ : Span4Mux_v
    port map (
            O => \N__14728\,
            I => \N__14713\
        );

    \I__2840\ : Span4Mux_h
    port map (
            O => \N__14725\,
            I => \N__14713\
        );

    \I__2839\ : Span4Mux_h
    port map (
            O => \N__14718\,
            I => \N__14710\
        );

    \I__2838\ : Odrv4
    port map (
            O => \N__14713\,
            I => \b2v_inst.stateZ0Z_7\
        );

    \I__2837\ : Odrv4
    port map (
            O => \N__14710\,
            I => \b2v_inst.stateZ0Z_7\
        );

    \I__2836\ : InMux
    port map (
            O => \N__14705\,
            I => \N__14701\
        );

    \I__2835\ : InMux
    port map (
            O => \N__14704\,
            I => \N__14698\
        );

    \I__2834\ : LocalMux
    port map (
            O => \N__14701\,
            I => \N__14695\
        );

    \I__2833\ : LocalMux
    port map (
            O => \N__14698\,
            I => \N__14690\
        );

    \I__2832\ : Span4Mux_v
    port map (
            O => \N__14695\,
            I => \N__14687\
        );

    \I__2831\ : InMux
    port map (
            O => \N__14694\,
            I => \N__14684\
        );

    \I__2830\ : InMux
    port map (
            O => \N__14693\,
            I => \N__14681\
        );

    \I__2829\ : Span4Mux_h
    port map (
            O => \N__14690\,
            I => \N__14678\
        );

    \I__2828\ : Span4Mux_h
    port map (
            O => \N__14687\,
            I => \N__14675\
        );

    \I__2827\ : LocalMux
    port map (
            O => \N__14684\,
            I => \N__14670\
        );

    \I__2826\ : LocalMux
    port map (
            O => \N__14681\,
            I => \N__14670\
        );

    \I__2825\ : Odrv4
    port map (
            O => \N__14678\,
            I => \SYNTHESIZED_WIRE_1_5\
        );

    \I__2824\ : Odrv4
    port map (
            O => \N__14675\,
            I => \SYNTHESIZED_WIRE_1_5\
        );

    \I__2823\ : Odrv12
    port map (
            O => \N__14670\,
            I => \SYNTHESIZED_WIRE_1_5\
        );

    \I__2822\ : InMux
    port map (
            O => \N__14663\,
            I => \N__14660\
        );

    \I__2821\ : LocalMux
    port map (
            O => \N__14660\,
            I => \N__14655\
        );

    \I__2820\ : InMux
    port map (
            O => \N__14659\,
            I => \N__14652\
        );

    \I__2819\ : InMux
    port map (
            O => \N__14658\,
            I => \N__14649\
        );

    \I__2818\ : Span4Mux_v
    port map (
            O => \N__14655\,
            I => \N__14643\
        );

    \I__2817\ : LocalMux
    port map (
            O => \N__14652\,
            I => \N__14643\
        );

    \I__2816\ : LocalMux
    port map (
            O => \N__14649\,
            I => \N__14640\
        );

    \I__2815\ : InMux
    port map (
            O => \N__14648\,
            I => \N__14637\
        );

    \I__2814\ : Span4Mux_h
    port map (
            O => \N__14643\,
            I => \N__14634\
        );

    \I__2813\ : Span4Mux_h
    port map (
            O => \N__14640\,
            I => \N__14631\
        );

    \I__2812\ : LocalMux
    port map (
            O => \N__14637\,
            I => \b2v_inst.reg_anteriorZ0Z_5\
        );

    \I__2811\ : Odrv4
    port map (
            O => \N__14634\,
            I => \b2v_inst.reg_anteriorZ0Z_5\
        );

    \I__2810\ : Odrv4
    port map (
            O => \N__14631\,
            I => \b2v_inst.reg_anteriorZ0Z_5\
        );

    \I__2809\ : CascadeMux
    port map (
            O => \N__14624\,
            I => \b2v_inst.un4_cuenta_ac0_11_0_cascade_\
        );

    \I__2808\ : InMux
    port map (
            O => \N__14621\,
            I => \N__14618\
        );

    \I__2807\ : LocalMux
    port map (
            O => \N__14618\,
            I => \N__14615\
        );

    \I__2806\ : Odrv4
    port map (
            O => \N__14615\,
            I => \b2v_inst.N_491\
        );

    \I__2805\ : CascadeMux
    port map (
            O => \N__14612\,
            I => \b2v_inst.cuenta_5_i_o2_0_0_1_cascade_\
        );

    \I__2804\ : CascadeMux
    port map (
            O => \N__14609\,
            I => \b2v_inst.state_ns_a2_0_o2_1_0_2_cascade_\
        );

    \I__2803\ : InMux
    port map (
            O => \N__14606\,
            I => \N__14602\
        );

    \I__2802\ : InMux
    port map (
            O => \N__14605\,
            I => \N__14599\
        );

    \I__2801\ : LocalMux
    port map (
            O => \N__14602\,
            I => \b2v_inst.cuenta_5_i_o2_0_0_1\
        );

    \I__2800\ : LocalMux
    port map (
            O => \N__14599\,
            I => \b2v_inst.cuenta_5_i_o2_0_0_1\
        );

    \I__2799\ : CascadeMux
    port map (
            O => \N__14594\,
            I => \b2v_inst.state_17_rep1_RNICDKZ0Z34_cascade_\
        );

    \I__2798\ : InMux
    port map (
            O => \N__14591\,
            I => \N__14588\
        );

    \I__2797\ : LocalMux
    port map (
            O => \N__14588\,
            I => \b2v_inst.cuenta_RNIO2VO3Z0Z_4\
        );

    \I__2796\ : InMux
    port map (
            O => \N__14585\,
            I => \N__14576\
        );

    \I__2795\ : InMux
    port map (
            O => \N__14584\,
            I => \N__14576\
        );

    \I__2794\ : InMux
    port map (
            O => \N__14583\,
            I => \N__14576\
        );

    \I__2793\ : LocalMux
    port map (
            O => \N__14576\,
            I => \b2v_inst.N_374\
        );

    \I__2792\ : InMux
    port map (
            O => \N__14573\,
            I => \N__14570\
        );

    \I__2791\ : LocalMux
    port map (
            O => \N__14570\,
            I => \N__14567\
        );

    \I__2790\ : Span4Mux_h
    port map (
            O => \N__14567\,
            I => \N__14564\
        );

    \I__2789\ : Odrv4
    port map (
            O => \N__14564\,
            I => \b2v_inst1.r_RX_Bytece_0_3\
        );

    \I__2788\ : InMux
    port map (
            O => \N__14561\,
            I => \N__14558\
        );

    \I__2787\ : LocalMux
    port map (
            O => \N__14558\,
            I => \N__14555\
        );

    \I__2786\ : Span4Mux_h
    port map (
            O => \N__14555\,
            I => \N__14552\
        );

    \I__2785\ : Odrv4
    port map (
            O => \N__14552\,
            I => \b2v_inst1.r_RX_Bytece_0_0_4\
        );

    \I__2784\ : InMux
    port map (
            O => \N__14549\,
            I => \N__14546\
        );

    \I__2783\ : LocalMux
    port map (
            O => \N__14546\,
            I => \N__14542\
        );

    \I__2782\ : InMux
    port map (
            O => \N__14545\,
            I => \N__14539\
        );

    \I__2781\ : Span4Mux_v
    port map (
            O => \N__14542\,
            I => \N__14536\
        );

    \I__2780\ : LocalMux
    port map (
            O => \N__14539\,
            I => \N__14533\
        );

    \I__2779\ : Span4Mux_h
    port map (
            O => \N__14536\,
            I => \N__14530\
        );

    \I__2778\ : Odrv12
    port map (
            O => \N__14533\,
            I => b2v_inst_data_a_escribir_3
        );

    \I__2777\ : Odrv4
    port map (
            O => \N__14530\,
            I => b2v_inst_data_a_escribir_3
        );

    \I__2776\ : InMux
    port map (
            O => \N__14525\,
            I => \N__14522\
        );

    \I__2775\ : LocalMux
    port map (
            O => \N__14522\,
            I => \N__14519\
        );

    \I__2774\ : Odrv4
    port map (
            O => \N__14519\,
            I => \b2v_inst3.data_to_sendZ0Z_3\
        );

    \I__2773\ : InMux
    port map (
            O => \N__14516\,
            I => \N__14513\
        );

    \I__2772\ : LocalMux
    port map (
            O => \N__14513\,
            I => \N__14510\
        );

    \I__2771\ : Span12Mux_v
    port map (
            O => \N__14510\,
            I => \N__14506\
        );

    \I__2770\ : InMux
    port map (
            O => \N__14509\,
            I => \N__14503\
        );

    \I__2769\ : Odrv12
    port map (
            O => \N__14506\,
            I => b2v_inst_data_a_escribir_4
        );

    \I__2768\ : LocalMux
    port map (
            O => \N__14503\,
            I => b2v_inst_data_a_escribir_4
        );

    \I__2767\ : CascadeMux
    port map (
            O => \N__14498\,
            I => \N__14495\
        );

    \I__2766\ : InMux
    port map (
            O => \N__14495\,
            I => \N__14492\
        );

    \I__2765\ : LocalMux
    port map (
            O => \N__14492\,
            I => \b2v_inst3.data_to_sendZ0Z_4\
        );

    \I__2764\ : InMux
    port map (
            O => \N__14489\,
            I => \N__14486\
        );

    \I__2763\ : LocalMux
    port map (
            O => \N__14486\,
            I => \N__14482\
        );

    \I__2762\ : InMux
    port map (
            O => \N__14485\,
            I => \N__14479\
        );

    \I__2761\ : Span4Mux_h
    port map (
            O => \N__14482\,
            I => \N__14476\
        );

    \I__2760\ : LocalMux
    port map (
            O => \N__14479\,
            I => \N__14473\
        );

    \I__2759\ : Span4Mux_v
    port map (
            O => \N__14476\,
            I => \N__14470\
        );

    \I__2758\ : Odrv12
    port map (
            O => \N__14473\,
            I => b2v_inst_data_a_escribir_5
        );

    \I__2757\ : Odrv4
    port map (
            O => \N__14470\,
            I => b2v_inst_data_a_escribir_5
        );

    \I__2756\ : CascadeMux
    port map (
            O => \N__14465\,
            I => \N__14462\
        );

    \I__2755\ : InMux
    port map (
            O => \N__14462\,
            I => \N__14459\
        );

    \I__2754\ : LocalMux
    port map (
            O => \N__14459\,
            I => \b2v_inst3.data_to_sendZ0Z_5\
        );

    \I__2753\ : InMux
    port map (
            O => \N__14456\,
            I => \N__14452\
        );

    \I__2752\ : InMux
    port map (
            O => \N__14455\,
            I => \N__14449\
        );

    \I__2751\ : LocalMux
    port map (
            O => \N__14452\,
            I => \N__14446\
        );

    \I__2750\ : LocalMux
    port map (
            O => \N__14449\,
            I => \N__14443\
        );

    \I__2749\ : Span4Mux_h
    port map (
            O => \N__14446\,
            I => \N__14440\
        );

    \I__2748\ : Span4Mux_v
    port map (
            O => \N__14443\,
            I => \N__14437\
        );

    \I__2747\ : Span4Mux_h
    port map (
            O => \N__14440\,
            I => \N__14434\
        );

    \I__2746\ : Odrv4
    port map (
            O => \N__14437\,
            I => b2v_inst_data_a_escribir_6
        );

    \I__2745\ : Odrv4
    port map (
            O => \N__14434\,
            I => b2v_inst_data_a_escribir_6
        );

    \I__2744\ : CascadeMux
    port map (
            O => \N__14429\,
            I => \N__14426\
        );

    \I__2743\ : InMux
    port map (
            O => \N__14426\,
            I => \N__14423\
        );

    \I__2742\ : LocalMux
    port map (
            O => \N__14423\,
            I => \b2v_inst3.data_to_sendZ0Z_6\
        );

    \I__2741\ : InMux
    port map (
            O => \N__14420\,
            I => \N__14410\
        );

    \I__2740\ : InMux
    port map (
            O => \N__14419\,
            I => \N__14405\
        );

    \I__2739\ : InMux
    port map (
            O => \N__14418\,
            I => \N__14405\
        );

    \I__2738\ : InMux
    port map (
            O => \N__14417\,
            I => \N__14394\
        );

    \I__2737\ : InMux
    port map (
            O => \N__14416\,
            I => \N__14394\
        );

    \I__2736\ : InMux
    port map (
            O => \N__14415\,
            I => \N__14394\
        );

    \I__2735\ : InMux
    port map (
            O => \N__14414\,
            I => \N__14394\
        );

    \I__2734\ : InMux
    port map (
            O => \N__14413\,
            I => \N__14394\
        );

    \I__2733\ : LocalMux
    port map (
            O => \N__14410\,
            I => \N__14389\
        );

    \I__2732\ : LocalMux
    port map (
            O => \N__14405\,
            I => \N__14389\
        );

    \I__2731\ : LocalMux
    port map (
            O => \N__14394\,
            I => \N__14386\
        );

    \I__2730\ : Span4Mux_v
    port map (
            O => \N__14389\,
            I => \N__14383\
        );

    \I__2729\ : Span4Mux_v
    port map (
            O => \N__14386\,
            I => \N__14380\
        );

    \I__2728\ : Odrv4
    port map (
            O => \N__14383\,
            I => \N_458\
        );

    \I__2727\ : Odrv4
    port map (
            O => \N__14380\,
            I => \N_458\
        );

    \I__2726\ : CascadeMux
    port map (
            O => \N__14375\,
            I => \N__14372\
        );

    \I__2725\ : InMux
    port map (
            O => \N__14372\,
            I => \N__14368\
        );

    \I__2724\ : InMux
    port map (
            O => \N__14371\,
            I => \N__14365\
        );

    \I__2723\ : LocalMux
    port map (
            O => \N__14368\,
            I => \N__14362\
        );

    \I__2722\ : LocalMux
    port map (
            O => \N__14365\,
            I => \N__14359\
        );

    \I__2721\ : Span4Mux_h
    port map (
            O => \N__14362\,
            I => \N__14356\
        );

    \I__2720\ : Span4Mux_h
    port map (
            O => \N__14359\,
            I => \N__14353\
        );

    \I__2719\ : Odrv4
    port map (
            O => \N__14356\,
            I => b2v_inst_data_a_escribir_7
        );

    \I__2718\ : Odrv4
    port map (
            O => \N__14353\,
            I => b2v_inst_data_a_escribir_7
        );

    \I__2717\ : InMux
    port map (
            O => \N__14348\,
            I => \N__14328\
        );

    \I__2716\ : InMux
    port map (
            O => \N__14347\,
            I => \N__14328\
        );

    \I__2715\ : InMux
    port map (
            O => \N__14346\,
            I => \N__14328\
        );

    \I__2714\ : InMux
    port map (
            O => \N__14345\,
            I => \N__14328\
        );

    \I__2713\ : InMux
    port map (
            O => \N__14344\,
            I => \N__14328\
        );

    \I__2712\ : InMux
    port map (
            O => \N__14343\,
            I => \N__14323\
        );

    \I__2711\ : InMux
    port map (
            O => \N__14342\,
            I => \N__14323\
        );

    \I__2710\ : InMux
    port map (
            O => \N__14341\,
            I => \N__14314\
        );

    \I__2709\ : InMux
    port map (
            O => \N__14340\,
            I => \N__14314\
        );

    \I__2708\ : InMux
    port map (
            O => \N__14339\,
            I => \N__14314\
        );

    \I__2707\ : LocalMux
    port map (
            O => \N__14328\,
            I => \N__14311\
        );

    \I__2706\ : LocalMux
    port map (
            O => \N__14323\,
            I => \N__14308\
        );

    \I__2705\ : InMux
    port map (
            O => \N__14322\,
            I => \N__14303\
        );

    \I__2704\ : InMux
    port map (
            O => \N__14321\,
            I => \N__14303\
        );

    \I__2703\ : LocalMux
    port map (
            O => \N__14314\,
            I => \N__14300\
        );

    \I__2702\ : Span4Mux_v
    port map (
            O => \N__14311\,
            I => \N__14295\
        );

    \I__2701\ : Span4Mux_h
    port map (
            O => \N__14308\,
            I => \N__14292\
        );

    \I__2700\ : LocalMux
    port map (
            O => \N__14303\,
            I => \N__14287\
        );

    \I__2699\ : Span12Mux_h
    port map (
            O => \N__14300\,
            I => \N__14287\
        );

    \I__2698\ : InMux
    port map (
            O => \N__14299\,
            I => \N__14282\
        );

    \I__2697\ : InMux
    port map (
            O => \N__14298\,
            I => \N__14282\
        );

    \I__2696\ : Span4Mux_v
    port map (
            O => \N__14295\,
            I => \N__14279\
        );

    \I__2695\ : Odrv4
    port map (
            O => \N__14292\,
            I => \N_230\
        );

    \I__2694\ : Odrv12
    port map (
            O => \N__14287\,
            I => \N_230\
        );

    \I__2693\ : LocalMux
    port map (
            O => \N__14282\,
            I => \N_230\
        );

    \I__2692\ : Odrv4
    port map (
            O => \N__14279\,
            I => \N_230\
        );

    \I__2691\ : CascadeMux
    port map (
            O => \N__14270\,
            I => \N__14266\
        );

    \I__2690\ : InMux
    port map (
            O => \N__14269\,
            I => \N__14261\
        );

    \I__2689\ : InMux
    port map (
            O => \N__14266\,
            I => \N__14261\
        );

    \I__2688\ : LocalMux
    port map (
            O => \N__14261\,
            I => \b2v_inst3.data_to_sendZ0Z_7\
        );

    \I__2687\ : CEMux
    port map (
            O => \N__14258\,
            I => \N__14255\
        );

    \I__2686\ : LocalMux
    port map (
            O => \N__14255\,
            I => \N__14251\
        );

    \I__2685\ : CEMux
    port map (
            O => \N__14254\,
            I => \N__14248\
        );

    \I__2684\ : Odrv12
    port map (
            O => \N__14251\,
            I => \b2v_inst3.un2_n_fsm_state_0_sqmuxa_2_0_i_0\
        );

    \I__2683\ : LocalMux
    port map (
            O => \N__14248\,
            I => \b2v_inst3.un2_n_fsm_state_0_sqmuxa_2_0_i_0\
        );

    \I__2682\ : InMux
    port map (
            O => \N__14243\,
            I => \N__14238\
        );

    \I__2681\ : InMux
    port map (
            O => \N__14242\,
            I => \N__14235\
        );

    \I__2680\ : InMux
    port map (
            O => \N__14241\,
            I => \N__14232\
        );

    \I__2679\ : LocalMux
    port map (
            O => \N__14238\,
            I => \N__14228\
        );

    \I__2678\ : LocalMux
    port map (
            O => \N__14235\,
            I => \N__14225\
        );

    \I__2677\ : LocalMux
    port map (
            O => \N__14232\,
            I => \N__14222\
        );

    \I__2676\ : InMux
    port map (
            O => \N__14231\,
            I => \N__14219\
        );

    \I__2675\ : Span4Mux_h
    port map (
            O => \N__14228\,
            I => \N__14216\
        );

    \I__2674\ : Span4Mux_v
    port map (
            O => \N__14225\,
            I => \N__14209\
        );

    \I__2673\ : Span4Mux_h
    port map (
            O => \N__14222\,
            I => \N__14209\
        );

    \I__2672\ : LocalMux
    port map (
            O => \N__14219\,
            I => \N__14209\
        );

    \I__2671\ : Odrv4
    port map (
            O => \N__14216\,
            I => \SYNTHESIZED_WIRE_1_6\
        );

    \I__2670\ : Odrv4
    port map (
            O => \N__14209\,
            I => \SYNTHESIZED_WIRE_1_6\
        );

    \I__2669\ : InMux
    port map (
            O => \N__14204\,
            I => \N__14201\
        );

    \I__2668\ : LocalMux
    port map (
            O => \N__14201\,
            I => \N__14195\
        );

    \I__2667\ : InMux
    port map (
            O => \N__14200\,
            I => \N__14192\
        );

    \I__2666\ : InMux
    port map (
            O => \N__14199\,
            I => \N__14189\
        );

    \I__2665\ : InMux
    port map (
            O => \N__14198\,
            I => \N__14186\
        );

    \I__2664\ : Span4Mux_h
    port map (
            O => \N__14195\,
            I => \N__14181\
        );

    \I__2663\ : LocalMux
    port map (
            O => \N__14192\,
            I => \N__14181\
        );

    \I__2662\ : LocalMux
    port map (
            O => \N__14189\,
            I => \N__14178\
        );

    \I__2661\ : LocalMux
    port map (
            O => \N__14186\,
            I => \b2v_inst.reg_anteriorZ0Z_6\
        );

    \I__2660\ : Odrv4
    port map (
            O => \N__14181\,
            I => \b2v_inst.reg_anteriorZ0Z_6\
        );

    \I__2659\ : Odrv12
    port map (
            O => \N__14178\,
            I => \b2v_inst.reg_anteriorZ0Z_6\
        );

    \I__2658\ : CascadeMux
    port map (
            O => \N__14171\,
            I => \b2v_inst.dir_mem_315_0_cascade_\
        );

    \I__2657\ : InMux
    port map (
            O => \N__14168\,
            I => \N__14165\
        );

    \I__2656\ : LocalMux
    port map (
            O => \N__14165\,
            I => \b2v_inst.dir_mem_3Z0Z_1\
        );

    \I__2655\ : InMux
    port map (
            O => \N__14162\,
            I => \N__14159\
        );

    \I__2654\ : LocalMux
    port map (
            O => \N__14159\,
            I => \b2v_inst.addr_ram_1_0_iv_i_1_1\
        );

    \I__2653\ : InMux
    port map (
            O => \N__14156\,
            I => \N__14153\
        );

    \I__2652\ : LocalMux
    port map (
            O => \N__14153\,
            I => \b2v_inst.dir_mem_3Z0Z_0\
        );

    \I__2651\ : CascadeMux
    port map (
            O => \N__14150\,
            I => \N__14147\
        );

    \I__2650\ : InMux
    port map (
            O => \N__14147\,
            I => \N__14144\
        );

    \I__2649\ : LocalMux
    port map (
            O => \N__14144\,
            I => \N__14141\
        );

    \I__2648\ : Span4Mux_v
    port map (
            O => \N__14141\,
            I => \N__14138\
        );

    \I__2647\ : Odrv4
    port map (
            O => \N__14138\,
            I => \b2v_inst.dir_mem_3Z0Z_5\
        );

    \I__2646\ : InMux
    port map (
            O => \N__14135\,
            I => \N__14132\
        );

    \I__2645\ : LocalMux
    port map (
            O => \N__14132\,
            I => \N__14129\
        );

    \I__2644\ : Odrv4
    port map (
            O => \N__14129\,
            I => \b2v_inst.dir_mem_3Z0Z_6\
        );

    \I__2643\ : InMux
    port map (
            O => \N__14126\,
            I => \N__14123\
        );

    \I__2642\ : LocalMux
    port map (
            O => \N__14123\,
            I => \N__14120\
        );

    \I__2641\ : Span4Mux_v
    port map (
            O => \N__14120\,
            I => \N__14117\
        );

    \I__2640\ : Span4Mux_h
    port map (
            O => \N__14117\,
            I => \N__14114\
        );

    \I__2639\ : Odrv4
    port map (
            O => \N__14114\,
            I => \N_205_i\
        );

    \I__2638\ : CascadeMux
    port map (
            O => \N__14111\,
            I => \N__14108\
        );

    \I__2637\ : InMux
    port map (
            O => \N__14108\,
            I => \N__14105\
        );

    \I__2636\ : LocalMux
    port map (
            O => \N__14105\,
            I => \N__14102\
        );

    \I__2635\ : Odrv4
    port map (
            O => \N__14102\,
            I => \b2v_inst.dir_mem_2Z0Z_6\
        );

    \I__2634\ : CascadeMux
    port map (
            O => \N__14099\,
            I => \b2v_inst.N_235_cascade_\
        );

    \I__2633\ : InMux
    port map (
            O => \N__14096\,
            I => \N__14089\
        );

    \I__2632\ : InMux
    port map (
            O => \N__14095\,
            I => \N__14089\
        );

    \I__2631\ : InMux
    port map (
            O => \N__14094\,
            I => \N__14086\
        );

    \I__2630\ : LocalMux
    port map (
            O => \N__14089\,
            I => \N__14083\
        );

    \I__2629\ : LocalMux
    port map (
            O => \N__14086\,
            I => \N__14078\
        );

    \I__2628\ : Span4Mux_h
    port map (
            O => \N__14083\,
            I => \N__14078\
        );

    \I__2627\ : Span4Mux_v
    port map (
            O => \N__14078\,
            I => \N__14075\
        );

    \I__2626\ : Odrv4
    port map (
            O => \N__14075\,
            I => \b2v_inst.stateZ0Z_11\
        );

    \I__2625\ : CascadeMux
    port map (
            O => \N__14072\,
            I => \b2v_inst.N_237_cascade_\
        );

    \I__2624\ : InMux
    port map (
            O => \N__14069\,
            I => \N__14066\
        );

    \I__2623\ : LocalMux
    port map (
            O => \N__14066\,
            I => \b2v_inst.addr_ram_1_iv_i_2_0\
        );

    \I__2622\ : CascadeMux
    port map (
            O => \N__14063\,
            I => \b2v_inst.addr_ram_1_iv_i_1_0_cascade_\
        );

    \I__2621\ : CascadeMux
    port map (
            O => \N__14060\,
            I => \N__14056\
        );

    \I__2620\ : CascadeMux
    port map (
            O => \N__14059\,
            I => \N__14053\
        );

    \I__2619\ : InMux
    port map (
            O => \N__14056\,
            I => \N__14050\
        );

    \I__2618\ : InMux
    port map (
            O => \N__14053\,
            I => \N__14047\
        );

    \I__2617\ : LocalMux
    port map (
            O => \N__14050\,
            I => \N__14044\
        );

    \I__2616\ : LocalMux
    port map (
            O => \N__14047\,
            I => \N__14041\
        );

    \I__2615\ : Span4Mux_v
    port map (
            O => \N__14044\,
            I => \N__14038\
        );

    \I__2614\ : Odrv4
    port map (
            O => \N__14041\,
            I => \N_167\
        );

    \I__2613\ : Odrv4
    port map (
            O => \N__14038\,
            I => \N_167\
        );

    \I__2612\ : InMux
    port map (
            O => \N__14033\,
            I => \N__14030\
        );

    \I__2611\ : LocalMux
    port map (
            O => \N__14030\,
            I => \b2v_inst.addr_ram_1_0_iv_i_0_1\
        );

    \I__2610\ : CascadeMux
    port map (
            O => \N__14027\,
            I => \N__14023\
        );

    \I__2609\ : CascadeMux
    port map (
            O => \N__14026\,
            I => \N__14020\
        );

    \I__2608\ : InMux
    port map (
            O => \N__14023\,
            I => \N__14017\
        );

    \I__2607\ : InMux
    port map (
            O => \N__14020\,
            I => \N__14014\
        );

    \I__2606\ : LocalMux
    port map (
            O => \N__14017\,
            I => \N__14011\
        );

    \I__2605\ : LocalMux
    port map (
            O => \N__14014\,
            I => \N__14006\
        );

    \I__2604\ : Span4Mux_v
    port map (
            O => \N__14011\,
            I => \N__14006\
        );

    \I__2603\ : Odrv4
    port map (
            O => \N__14006\,
            I => \N_60\
        );

    \I__2602\ : CascadeMux
    port map (
            O => \N__14003\,
            I => \b2v_inst.addr_ram_1_0_iv_i_0_2_cascade_\
        );

    \I__2601\ : CascadeMux
    port map (
            O => \N__14000\,
            I => \N__13996\
        );

    \I__2600\ : CascadeMux
    port map (
            O => \N__13999\,
            I => \N__13993\
        );

    \I__2599\ : InMux
    port map (
            O => \N__13996\,
            I => \N__13990\
        );

    \I__2598\ : InMux
    port map (
            O => \N__13993\,
            I => \N__13987\
        );

    \I__2597\ : LocalMux
    port map (
            O => \N__13990\,
            I => \N__13984\
        );

    \I__2596\ : LocalMux
    port map (
            O => \N__13987\,
            I => \N__13981\
        );

    \I__2595\ : Span4Mux_h
    port map (
            O => \N__13984\,
            I => \N__13978\
        );

    \I__2594\ : Odrv4
    port map (
            O => \N__13981\,
            I => \N_56\
        );

    \I__2593\ : Odrv4
    port map (
            O => \N__13978\,
            I => \N_56\
        );

    \I__2592\ : CascadeMux
    port map (
            O => \N__13973\,
            I => \b2v_inst.N_236_cascade_\
        );

    \I__2591\ : InMux
    port map (
            O => \N__13970\,
            I => \N__13967\
        );

    \I__2590\ : LocalMux
    port map (
            O => \N__13967\,
            I => \N__13964\
        );

    \I__2589\ : Span4Mux_h
    port map (
            O => \N__13964\,
            I => \N__13959\
        );

    \I__2588\ : InMux
    port map (
            O => \N__13963\,
            I => \N__13954\
        );

    \I__2587\ : InMux
    port map (
            O => \N__13962\,
            I => \N__13954\
        );

    \I__2586\ : Odrv4
    port map (
            O => \N__13959\,
            I => \b2v_inst.stateZ0Z_9\
        );

    \I__2585\ : LocalMux
    port map (
            O => \N__13954\,
            I => \b2v_inst.stateZ0Z_9\
        );

    \I__2584\ : CascadeMux
    port map (
            O => \N__13949\,
            I => \b2v_inst.N_399_cascade_\
        );

    \I__2583\ : InMux
    port map (
            O => \N__13946\,
            I => \N__13943\
        );

    \I__2582\ : LocalMux
    port map (
            O => \N__13943\,
            I => \b2v_inst.addr_ram_1_iv_i_1_6\
        );

    \I__2581\ : CascadeMux
    port map (
            O => \N__13940\,
            I => \b2v_inst.addr_ram_1_iv_i_2_6_cascade_\
        );

    \I__2580\ : CascadeMux
    port map (
            O => \N__13937\,
            I => \N__13933\
        );

    \I__2579\ : CascadeMux
    port map (
            O => \N__13936\,
            I => \N__13930\
        );

    \I__2578\ : InMux
    port map (
            O => \N__13933\,
            I => \N__13927\
        );

    \I__2577\ : InMux
    port map (
            O => \N__13930\,
            I => \N__13924\
        );

    \I__2576\ : LocalMux
    port map (
            O => \N__13927\,
            I => \N__13919\
        );

    \I__2575\ : LocalMux
    port map (
            O => \N__13924\,
            I => \N__13919\
        );

    \I__2574\ : Span4Mux_v
    port map (
            O => \N__13919\,
            I => \N__13916\
        );

    \I__2573\ : Odrv4
    port map (
            O => \N__13916\,
            I => \N_165\
        );

    \I__2572\ : CEMux
    port map (
            O => \N__13913\,
            I => \N__13909\
        );

    \I__2571\ : CEMux
    port map (
            O => \N__13912\,
            I => \N__13906\
        );

    \I__2570\ : LocalMux
    port map (
            O => \N__13909\,
            I => \N__13903\
        );

    \I__2569\ : LocalMux
    port map (
            O => \N__13906\,
            I => \N__13900\
        );

    \I__2568\ : Span4Mux_h
    port map (
            O => \N__13903\,
            I => \N__13895\
        );

    \I__2567\ : Span4Mux_h
    port map (
            O => \N__13900\,
            I => \N__13895\
        );

    \I__2566\ : Span4Mux_h
    port map (
            O => \N__13895\,
            I => \N__13889\
        );

    \I__2565\ : InMux
    port map (
            O => \N__13894\,
            I => \N__13886\
        );

    \I__2564\ : InMux
    port map (
            O => \N__13893\,
            I => \N__13881\
        );

    \I__2563\ : InMux
    port map (
            O => \N__13892\,
            I => \N__13881\
        );

    \I__2562\ : Odrv4
    port map (
            O => \N__13889\,
            I => \b2v_inst.stateZ0Z_12\
        );

    \I__2561\ : LocalMux
    port map (
            O => \N__13886\,
            I => \b2v_inst.stateZ0Z_12\
        );

    \I__2560\ : LocalMux
    port map (
            O => \N__13881\,
            I => \b2v_inst.stateZ0Z_12\
        );

    \I__2559\ : CascadeMux
    port map (
            O => \N__13874\,
            I => \b2v_inst.un2_cuentalto7_3_cascade_\
        );

    \I__2558\ : CascadeMux
    port map (
            O => \N__13871\,
            I => \b2v_inst.N_351_0_cascade_\
        );

    \I__2557\ : CascadeMux
    port map (
            O => \N__13868\,
            I => \N__13864\
        );

    \I__2556\ : InMux
    port map (
            O => \N__13867\,
            I => \N__13861\
        );

    \I__2555\ : InMux
    port map (
            O => \N__13864\,
            I => \N__13858\
        );

    \I__2554\ : LocalMux
    port map (
            O => \N__13861\,
            I => \b2v_inst.cuenta_fastZ0Z_4\
        );

    \I__2553\ : LocalMux
    port map (
            O => \N__13858\,
            I => \b2v_inst.cuenta_fastZ0Z_4\
        );

    \I__2552\ : InMux
    port map (
            O => \N__13853\,
            I => \N__13848\
        );

    \I__2551\ : InMux
    port map (
            O => \N__13852\,
            I => \N__13845\
        );

    \I__2550\ : InMux
    port map (
            O => \N__13851\,
            I => \N__13842\
        );

    \I__2549\ : LocalMux
    port map (
            O => \N__13848\,
            I => \b2v_inst.cuenta_RNIQ56K_0Z0Z_3\
        );

    \I__2548\ : LocalMux
    port map (
            O => \N__13845\,
            I => \b2v_inst.cuenta_RNIQ56K_0Z0Z_3\
        );

    \I__2547\ : LocalMux
    port map (
            O => \N__13842\,
            I => \b2v_inst.cuenta_RNIQ56K_0Z0Z_3\
        );

    \I__2546\ : InMux
    port map (
            O => \N__13835\,
            I => \N__13832\
        );

    \I__2545\ : LocalMux
    port map (
            O => \N__13832\,
            I => \b2v_inst.N_376_1\
        );

    \I__2544\ : InMux
    port map (
            O => \N__13829\,
            I => \N__13823\
        );

    \I__2543\ : InMux
    port map (
            O => \N__13828\,
            I => \N__13823\
        );

    \I__2542\ : LocalMux
    port map (
            O => \N__13823\,
            I => \b2v_inst.cuenta_RNIQI4FZ0Z_2\
        );

    \I__2541\ : CascadeMux
    port map (
            O => \N__13820\,
            I => \N__13817\
        );

    \I__2540\ : InMux
    port map (
            O => \N__13817\,
            I => \N__13811\
        );

    \I__2539\ : InMux
    port map (
            O => \N__13816\,
            I => \N__13811\
        );

    \I__2538\ : LocalMux
    port map (
            O => \N__13811\,
            I => \b2v_inst.cuenta_RNIR03AZ0Z_1\
        );

    \I__2537\ : CascadeMux
    port map (
            O => \N__13808\,
            I => \b2v_inst.N_376_1_cascade_\
        );

    \I__2536\ : CascadeMux
    port map (
            O => \N__13805\,
            I => \N__13797\
        );

    \I__2535\ : InMux
    port map (
            O => \N__13804\,
            I => \N__13793\
        );

    \I__2534\ : InMux
    port map (
            O => \N__13803\,
            I => \N__13790\
        );

    \I__2533\ : InMux
    port map (
            O => \N__13802\,
            I => \N__13787\
        );

    \I__2532\ : InMux
    port map (
            O => \N__13801\,
            I => \N__13778\
        );

    \I__2531\ : InMux
    port map (
            O => \N__13800\,
            I => \N__13778\
        );

    \I__2530\ : InMux
    port map (
            O => \N__13797\,
            I => \N__13778\
        );

    \I__2529\ : InMux
    port map (
            O => \N__13796\,
            I => \N__13778\
        );

    \I__2528\ : LocalMux
    port map (
            O => \N__13793\,
            I => \b2v_inst.cuentaZ0Z_1\
        );

    \I__2527\ : LocalMux
    port map (
            O => \N__13790\,
            I => \b2v_inst.cuentaZ0Z_1\
        );

    \I__2526\ : LocalMux
    port map (
            O => \N__13787\,
            I => \b2v_inst.cuentaZ0Z_1\
        );

    \I__2525\ : LocalMux
    port map (
            O => \N__13778\,
            I => \b2v_inst.cuentaZ0Z_1\
        );

    \I__2524\ : InMux
    port map (
            O => \N__13769\,
            I => \N__13766\
        );

    \I__2523\ : LocalMux
    port map (
            O => \N__13766\,
            I => \N__13763\
        );

    \I__2522\ : Odrv4
    port map (
            O => \N__13763\,
            I => \b2v_inst.cuenta_5_i_a2_0_3\
        );

    \I__2521\ : InMux
    port map (
            O => \N__13760\,
            I => \N__13754\
        );

    \I__2520\ : InMux
    port map (
            O => \N__13759\,
            I => \N__13751\
        );

    \I__2519\ : InMux
    port map (
            O => \N__13758\,
            I => \N__13746\
        );

    \I__2518\ : InMux
    port map (
            O => \N__13757\,
            I => \N__13746\
        );

    \I__2517\ : LocalMux
    port map (
            O => \N__13754\,
            I => \N__13734\
        );

    \I__2516\ : LocalMux
    port map (
            O => \N__13751\,
            I => \N__13734\
        );

    \I__2515\ : LocalMux
    port map (
            O => \N__13746\,
            I => \N__13734\
        );

    \I__2514\ : InMux
    port map (
            O => \N__13745\,
            I => \N__13723\
        );

    \I__2513\ : InMux
    port map (
            O => \N__13744\,
            I => \N__13723\
        );

    \I__2512\ : InMux
    port map (
            O => \N__13743\,
            I => \N__13723\
        );

    \I__2511\ : InMux
    port map (
            O => \N__13742\,
            I => \N__13723\
        );

    \I__2510\ : InMux
    port map (
            O => \N__13741\,
            I => \N__13723\
        );

    \I__2509\ : Odrv4
    port map (
            O => \N__13734\,
            I => \b2v_inst.cuentaZ0Z_0\
        );

    \I__2508\ : LocalMux
    port map (
            O => \N__13723\,
            I => \b2v_inst.cuentaZ0Z_0\
        );

    \I__2507\ : InMux
    port map (
            O => \N__13718\,
            I => \N__13715\
        );

    \I__2506\ : LocalMux
    port map (
            O => \N__13715\,
            I => \b2v_inst.N_377\
        );

    \I__2505\ : CascadeMux
    port map (
            O => \N__13712\,
            I => \b2v_inst.N_491_cascade_\
        );

    \I__2504\ : InMux
    port map (
            O => \N__13709\,
            I => \N__13706\
        );

    \I__2503\ : LocalMux
    port map (
            O => \N__13706\,
            I => \N__13703\
        );

    \I__2502\ : Span4Mux_h
    port map (
            O => \N__13703\,
            I => \N__13700\
        );

    \I__2501\ : Odrv4
    port map (
            O => \N__13700\,
            I => \b2v_inst.state_RNIFQKOZ0Z_17\
        );

    \I__2500\ : CascadeMux
    port map (
            O => \N__13697\,
            I => \b2v_inst.state_RNIFQKOZ0Z_17_cascade_\
        );

    \I__2499\ : CascadeMux
    port map (
            O => \N__13694\,
            I => \b2v_inst.cuenta_5_i_a2_2_0_1_cascade_\
        );

    \I__2498\ : CascadeMux
    port map (
            O => \N__13691\,
            I => \b2v_inst.un4_cuenta_c4_cascade_\
        );

    \I__2497\ : CascadeMux
    port map (
            O => \N__13688\,
            I => \N__13683\
        );

    \I__2496\ : InMux
    port map (
            O => \N__13687\,
            I => \N__13680\
        );

    \I__2495\ : InMux
    port map (
            O => \N__13686\,
            I => \N__13675\
        );

    \I__2494\ : InMux
    port map (
            O => \N__13683\,
            I => \N__13675\
        );

    \I__2493\ : LocalMux
    port map (
            O => \N__13680\,
            I => \b2v_inst.cuentaZ0Z_3\
        );

    \I__2492\ : LocalMux
    port map (
            O => \N__13675\,
            I => \b2v_inst.cuentaZ0Z_3\
        );

    \I__2491\ : InMux
    port map (
            O => \N__13670\,
            I => \N__13662\
        );

    \I__2490\ : InMux
    port map (
            O => \N__13669\,
            I => \N__13659\
        );

    \I__2489\ : InMux
    port map (
            O => \N__13668\,
            I => \N__13650\
        );

    \I__2488\ : InMux
    port map (
            O => \N__13667\,
            I => \N__13650\
        );

    \I__2487\ : InMux
    port map (
            O => \N__13666\,
            I => \N__13650\
        );

    \I__2486\ : InMux
    port map (
            O => \N__13665\,
            I => \N__13650\
        );

    \I__2485\ : LocalMux
    port map (
            O => \N__13662\,
            I => \b2v_inst.cuentaZ0Z_2\
        );

    \I__2484\ : LocalMux
    port map (
            O => \N__13659\,
            I => \b2v_inst.cuentaZ0Z_2\
        );

    \I__2483\ : LocalMux
    port map (
            O => \N__13650\,
            I => \b2v_inst.cuentaZ0Z_2\
        );

    \I__2482\ : InMux
    port map (
            O => \N__13643\,
            I => \N__13639\
        );

    \I__2481\ : InMux
    port map (
            O => \N__13642\,
            I => \N__13635\
        );

    \I__2480\ : LocalMux
    port map (
            O => \N__13639\,
            I => \N__13632\
        );

    \I__2479\ : InMux
    port map (
            O => \N__13638\,
            I => \N__13629\
        );

    \I__2478\ : LocalMux
    port map (
            O => \N__13635\,
            I => \N__13626\
        );

    \I__2477\ : Span4Mux_v
    port map (
            O => \N__13632\,
            I => \N__13623\
        );

    \I__2476\ : LocalMux
    port map (
            O => \N__13629\,
            I => \N__13620\
        );

    \I__2475\ : Span4Mux_v
    port map (
            O => \N__13626\,
            I => \N__13612\
        );

    \I__2474\ : Span4Mux_h
    port map (
            O => \N__13623\,
            I => \N__13612\
        );

    \I__2473\ : Span4Mux_h
    port map (
            O => \N__13620\,
            I => \N__13612\
        );

    \I__2472\ : InMux
    port map (
            O => \N__13619\,
            I => \N__13609\
        );

    \I__2471\ : Odrv4
    port map (
            O => \N__13612\,
            I => \SYNTHESIZED_WIRE_1_7\
        );

    \I__2470\ : LocalMux
    port map (
            O => \N__13609\,
            I => \SYNTHESIZED_WIRE_1_7\
        );

    \I__2469\ : InMux
    port map (
            O => \N__13604\,
            I => \N__13598\
        );

    \I__2468\ : CascadeMux
    port map (
            O => \N__13603\,
            I => \N__13595\
        );

    \I__2467\ : InMux
    port map (
            O => \N__13602\,
            I => \N__13592\
        );

    \I__2466\ : InMux
    port map (
            O => \N__13601\,
            I => \N__13589\
        );

    \I__2465\ : LocalMux
    port map (
            O => \N__13598\,
            I => \N__13586\
        );

    \I__2464\ : InMux
    port map (
            O => \N__13595\,
            I => \N__13583\
        );

    \I__2463\ : LocalMux
    port map (
            O => \N__13592\,
            I => \N__13578\
        );

    \I__2462\ : LocalMux
    port map (
            O => \N__13589\,
            I => \N__13578\
        );

    \I__2461\ : Span4Mux_h
    port map (
            O => \N__13586\,
            I => \N__13575\
        );

    \I__2460\ : LocalMux
    port map (
            O => \N__13583\,
            I => \b2v_inst.reg_anteriorZ0Z_7\
        );

    \I__2459\ : Odrv4
    port map (
            O => \N__13578\,
            I => \b2v_inst.reg_anteriorZ0Z_7\
        );

    \I__2458\ : Odrv4
    port map (
            O => \N__13575\,
            I => \b2v_inst.reg_anteriorZ0Z_7\
        );

    \I__2457\ : InMux
    port map (
            O => \N__13568\,
            I => \N__13565\
        );

    \I__2456\ : LocalMux
    port map (
            O => \N__13565\,
            I => \N__13562\
        );

    \I__2455\ : Span4Mux_h
    port map (
            O => \N__13562\,
            I => \N__13559\
        );

    \I__2454\ : Span4Mux_v
    port map (
            O => \N__13559\,
            I => \N__13556\
        );

    \I__2453\ : Odrv4
    port map (
            O => \N__13556\,
            I => \b2v_inst.data_a_escribir9_7_and\
        );

    \I__2452\ : InMux
    port map (
            O => \N__13553\,
            I => \N__13549\
        );

    \I__2451\ : InMux
    port map (
            O => \N__13552\,
            I => \N__13546\
        );

    \I__2450\ : LocalMux
    port map (
            O => \N__13549\,
            I => \N__13542\
        );

    \I__2449\ : LocalMux
    port map (
            O => \N__13546\,
            I => \N__13539\
        );

    \I__2448\ : InMux
    port map (
            O => \N__13545\,
            I => \N__13536\
        );

    \I__2447\ : Span4Mux_h
    port map (
            O => \N__13542\,
            I => \N__13532\
        );

    \I__2446\ : Span12Mux_h
    port map (
            O => \N__13539\,
            I => \N__13529\
        );

    \I__2445\ : LocalMux
    port map (
            O => \N__13536\,
            I => \N__13526\
        );

    \I__2444\ : InMux
    port map (
            O => \N__13535\,
            I => \N__13523\
        );

    \I__2443\ : Odrv4
    port map (
            O => \N__13532\,
            I => \SYNTHESIZED_WIRE_1_4\
        );

    \I__2442\ : Odrv12
    port map (
            O => \N__13529\,
            I => \SYNTHESIZED_WIRE_1_4\
        );

    \I__2441\ : Odrv12
    port map (
            O => \N__13526\,
            I => \SYNTHESIZED_WIRE_1_4\
        );

    \I__2440\ : LocalMux
    port map (
            O => \N__13523\,
            I => \SYNTHESIZED_WIRE_1_4\
        );

    \I__2439\ : InMux
    port map (
            O => \N__13514\,
            I => \N__13510\
        );

    \I__2438\ : InMux
    port map (
            O => \N__13513\,
            I => \N__13505\
        );

    \I__2437\ : LocalMux
    port map (
            O => \N__13510\,
            I => \N__13502\
        );

    \I__2436\ : InMux
    port map (
            O => \N__13509\,
            I => \N__13499\
        );

    \I__2435\ : InMux
    port map (
            O => \N__13508\,
            I => \N__13496\
        );

    \I__2434\ : LocalMux
    port map (
            O => \N__13505\,
            I => \N__13493\
        );

    \I__2433\ : Span4Mux_v
    port map (
            O => \N__13502\,
            I => \N__13488\
        );

    \I__2432\ : LocalMux
    port map (
            O => \N__13499\,
            I => \N__13488\
        );

    \I__2431\ : LocalMux
    port map (
            O => \N__13496\,
            I => \b2v_inst.reg_anteriorZ0Z_4\
        );

    \I__2430\ : Odrv4
    port map (
            O => \N__13493\,
            I => \b2v_inst.reg_anteriorZ0Z_4\
        );

    \I__2429\ : Odrv4
    port map (
            O => \N__13488\,
            I => \b2v_inst.reg_anteriorZ0Z_4\
        );

    \I__2428\ : InMux
    port map (
            O => \N__13481\,
            I => \N__13477\
        );

    \I__2427\ : CascadeMux
    port map (
            O => \N__13480\,
            I => \N__13474\
        );

    \I__2426\ : LocalMux
    port map (
            O => \N__13477\,
            I => \N__13471\
        );

    \I__2425\ : InMux
    port map (
            O => \N__13474\,
            I => \N__13468\
        );

    \I__2424\ : Span4Mux_h
    port map (
            O => \N__13471\,
            I => \N__13463\
        );

    \I__2423\ : LocalMux
    port map (
            O => \N__13468\,
            I => \N__13463\
        );

    \I__2422\ : Odrv4
    port map (
            O => \N__13463\,
            I => b2v_inst_data_a_escribir_1
        );

    \I__2421\ : InMux
    port map (
            O => \N__13460\,
            I => \N__13456\
        );

    \I__2420\ : CascadeMux
    port map (
            O => \N__13459\,
            I => \N__13453\
        );

    \I__2419\ : LocalMux
    port map (
            O => \N__13456\,
            I => \N__13450\
        );

    \I__2418\ : InMux
    port map (
            O => \N__13453\,
            I => \N__13447\
        );

    \I__2417\ : Span4Mux_v
    port map (
            O => \N__13450\,
            I => \N__13444\
        );

    \I__2416\ : LocalMux
    port map (
            O => \N__13447\,
            I => \N__13441\
        );

    \I__2415\ : Odrv4
    port map (
            O => \N__13444\,
            I => b2v_inst_data_a_escribir_0
        );

    \I__2414\ : Odrv4
    port map (
            O => \N__13441\,
            I => b2v_inst_data_a_escribir_0
        );

    \I__2413\ : CascadeMux
    port map (
            O => \N__13436\,
            I => \N__13433\
        );

    \I__2412\ : InMux
    port map (
            O => \N__13433\,
            I => \N__13430\
        );

    \I__2411\ : LocalMux
    port map (
            O => \N__13430\,
            I => \b2v_inst3.data_to_sendZ0Z_1\
        );

    \I__2410\ : InMux
    port map (
            O => \N__13427\,
            I => \N__13424\
        );

    \I__2409\ : LocalMux
    port map (
            O => \N__13424\,
            I => \N__13421\
        );

    \I__2408\ : Span12Mux_v
    port map (
            O => \N__13421\,
            I => \N__13418\
        );

    \I__2407\ : Odrv12
    port map (
            O => \N__13418\,
            I => \b2v_inst3.data_to_sendZ0Z_0\
        );

    \I__2406\ : CascadeMux
    port map (
            O => \N__13415\,
            I => \N__13412\
        );

    \I__2405\ : InMux
    port map (
            O => \N__13412\,
            I => \N__13408\
        );

    \I__2404\ : InMux
    port map (
            O => \N__13411\,
            I => \N__13405\
        );

    \I__2403\ : LocalMux
    port map (
            O => \N__13408\,
            I => \N__13402\
        );

    \I__2402\ : LocalMux
    port map (
            O => \N__13405\,
            I => \N__13399\
        );

    \I__2401\ : Span4Mux_h
    port map (
            O => \N__13402\,
            I => \N__13394\
        );

    \I__2400\ : Span4Mux_h
    port map (
            O => \N__13399\,
            I => \N__13394\
        );

    \I__2399\ : Odrv4
    port map (
            O => \N__13394\,
            I => b2v_inst_data_a_escribir_2
        );

    \I__2398\ : CascadeMux
    port map (
            O => \N__13391\,
            I => \N__13388\
        );

    \I__2397\ : InMux
    port map (
            O => \N__13388\,
            I => \N__13385\
        );

    \I__2396\ : LocalMux
    port map (
            O => \N__13385\,
            I => \b2v_inst3.data_to_sendZ0Z_2\
        );

    \I__2395\ : CascadeMux
    port map (
            O => \N__13382\,
            I => \N__13376\
        );

    \I__2394\ : InMux
    port map (
            O => \N__13381\,
            I => \N__13373\
        );

    \I__2393\ : InMux
    port map (
            O => \N__13380\,
            I => \N__13370\
        );

    \I__2392\ : InMux
    port map (
            O => \N__13379\,
            I => \N__13365\
        );

    \I__2391\ : InMux
    port map (
            O => \N__13376\,
            I => \N__13365\
        );

    \I__2390\ : LocalMux
    port map (
            O => \N__13373\,
            I => \b2v_inst3.fsm_state_RNIEPSN1Z0Z_0\
        );

    \I__2389\ : LocalMux
    port map (
            O => \N__13370\,
            I => \b2v_inst3.fsm_state_RNIEPSN1Z0Z_0\
        );

    \I__2388\ : LocalMux
    port map (
            O => \N__13365\,
            I => \b2v_inst3.fsm_state_RNIEPSN1Z0Z_0\
        );

    \I__2387\ : InMux
    port map (
            O => \N__13358\,
            I => \N__13352\
        );

    \I__2386\ : InMux
    port map (
            O => \N__13357\,
            I => \N__13344\
        );

    \I__2385\ : InMux
    port map (
            O => \N__13356\,
            I => \N__13339\
        );

    \I__2384\ : InMux
    port map (
            O => \N__13355\,
            I => \N__13339\
        );

    \I__2383\ : LocalMux
    port map (
            O => \N__13352\,
            I => \N__13336\
        );

    \I__2382\ : InMux
    port map (
            O => \N__13351\,
            I => \N__13333\
        );

    \I__2381\ : InMux
    port map (
            O => \N__13350\,
            I => \N__13330\
        );

    \I__2380\ : InMux
    port map (
            O => \N__13349\,
            I => \N__13325\
        );

    \I__2379\ : InMux
    port map (
            O => \N__13348\,
            I => \N__13325\
        );

    \I__2378\ : InMux
    port map (
            O => \N__13347\,
            I => \N__13322\
        );

    \I__2377\ : LocalMux
    port map (
            O => \N__13344\,
            I => \N__13317\
        );

    \I__2376\ : LocalMux
    port map (
            O => \N__13339\,
            I => \N__13317\
        );

    \I__2375\ : Odrv4
    port map (
            O => \N__13336\,
            I => \b2v_inst3.N_105_7\
        );

    \I__2374\ : LocalMux
    port map (
            O => \N__13333\,
            I => \b2v_inst3.N_105_7\
        );

    \I__2373\ : LocalMux
    port map (
            O => \N__13330\,
            I => \b2v_inst3.N_105_7\
        );

    \I__2372\ : LocalMux
    port map (
            O => \N__13325\,
            I => \b2v_inst3.N_105_7\
        );

    \I__2371\ : LocalMux
    port map (
            O => \N__13322\,
            I => \b2v_inst3.N_105_7\
        );

    \I__2370\ : Odrv4
    port map (
            O => \N__13317\,
            I => \b2v_inst3.N_105_7\
        );

    \I__2369\ : InMux
    port map (
            O => \N__13304\,
            I => \N__13297\
        );

    \I__2368\ : InMux
    port map (
            O => \N__13303\,
            I => \N__13294\
        );

    \I__2367\ : InMux
    port map (
            O => \N__13302\,
            I => \N__13287\
        );

    \I__2366\ : InMux
    port map (
            O => \N__13301\,
            I => \N__13287\
        );

    \I__2365\ : InMux
    port map (
            O => \N__13300\,
            I => \N__13287\
        );

    \I__2364\ : LocalMux
    port map (
            O => \N__13297\,
            I => \b2v_inst3.bit_counterZ0Z_0\
        );

    \I__2363\ : LocalMux
    port map (
            O => \N__13294\,
            I => \b2v_inst3.bit_counterZ0Z_0\
        );

    \I__2362\ : LocalMux
    port map (
            O => \N__13287\,
            I => \b2v_inst3.bit_counterZ0Z_0\
        );

    \I__2361\ : CascadeMux
    port map (
            O => \N__13280\,
            I => \N__13277\
        );

    \I__2360\ : InMux
    port map (
            O => \N__13277\,
            I => \N__13274\
        );

    \I__2359\ : LocalMux
    port map (
            O => \N__13274\,
            I => \b2v_inst.state_ns_a2_0_a2_0_1_2\
        );

    \I__2358\ : CascadeMux
    port map (
            O => \N__13271\,
            I => \N__13268\
        );

    \I__2357\ : InMux
    port map (
            O => \N__13268\,
            I => \N__13263\
        );

    \I__2356\ : CascadeMux
    port map (
            O => \N__13267\,
            I => \N__13260\
        );

    \I__2355\ : CascadeMux
    port map (
            O => \N__13266\,
            I => \N__13257\
        );

    \I__2354\ : LocalMux
    port map (
            O => \N__13263\,
            I => \N__13254\
        );

    \I__2353\ : InMux
    port map (
            O => \N__13260\,
            I => \N__13251\
        );

    \I__2352\ : InMux
    port map (
            O => \N__13257\,
            I => \N__13248\
        );

    \I__2351\ : Odrv4
    port map (
            O => \N__13254\,
            I => \b2v_inst.reg_ancho_3_i_7\
        );

    \I__2350\ : LocalMux
    port map (
            O => \N__13251\,
            I => \b2v_inst.reg_ancho_3_i_7\
        );

    \I__2349\ : LocalMux
    port map (
            O => \N__13248\,
            I => \b2v_inst.reg_ancho_3_i_7\
        );

    \I__2348\ : InMux
    port map (
            O => \N__13241\,
            I => \bfn_6_18_0_\
        );

    \I__2347\ : CascadeMux
    port map (
            O => \N__13238\,
            I => \N__13234\
        );

    \I__2346\ : InMux
    port map (
            O => \N__13237\,
            I => \N__13224\
        );

    \I__2345\ : InMux
    port map (
            O => \N__13234\,
            I => \N__13220\
        );

    \I__2344\ : InMux
    port map (
            O => \N__13233\,
            I => \N__13215\
        );

    \I__2343\ : InMux
    port map (
            O => \N__13232\,
            I => \N__13210\
        );

    \I__2342\ : InMux
    port map (
            O => \N__13231\,
            I => \N__13210\
        );

    \I__2341\ : InMux
    port map (
            O => \N__13230\,
            I => \N__13207\
        );

    \I__2340\ : InMux
    port map (
            O => \N__13229\,
            I => \N__13204\
        );

    \I__2339\ : InMux
    port map (
            O => \N__13228\,
            I => \N__13199\
        );

    \I__2338\ : InMux
    port map (
            O => \N__13227\,
            I => \N__13199\
        );

    \I__2337\ : LocalMux
    port map (
            O => \N__13224\,
            I => \N__13196\
        );

    \I__2336\ : InMux
    port map (
            O => \N__13223\,
            I => \N__13193\
        );

    \I__2335\ : LocalMux
    port map (
            O => \N__13220\,
            I => \N__13190\
        );

    \I__2334\ : InMux
    port map (
            O => \N__13219\,
            I => \N__13185\
        );

    \I__2333\ : InMux
    port map (
            O => \N__13218\,
            I => \N__13185\
        );

    \I__2332\ : LocalMux
    port map (
            O => \N__13215\,
            I => \N__13180\
        );

    \I__2331\ : LocalMux
    port map (
            O => \N__13210\,
            I => \N__13180\
        );

    \I__2330\ : LocalMux
    port map (
            O => \N__13207\,
            I => \N__13173\
        );

    \I__2329\ : LocalMux
    port map (
            O => \N__13204\,
            I => \N__13173\
        );

    \I__2328\ : LocalMux
    port map (
            O => \N__13199\,
            I => \N__13173\
        );

    \I__2327\ : Span4Mux_v
    port map (
            O => \N__13196\,
            I => \N__13170\
        );

    \I__2326\ : LocalMux
    port map (
            O => \N__13193\,
            I => \N__13163\
        );

    \I__2325\ : Span12Mux_s8_v
    port map (
            O => \N__13190\,
            I => \N__13163\
        );

    \I__2324\ : LocalMux
    port map (
            O => \N__13185\,
            I => \N__13163\
        );

    \I__2323\ : Span4Mux_h
    port map (
            O => \N__13180\,
            I => \N__13158\
        );

    \I__2322\ : Span4Mux_h
    port map (
            O => \N__13173\,
            I => \N__13158\
        );

    \I__2321\ : Odrv4
    port map (
            O => \N__13170\,
            I => \b2v_inst.un3_valor_max2_THRU_CO\
        );

    \I__2320\ : Odrv12
    port map (
            O => \N__13163\,
            I => \b2v_inst.un3_valor_max2_THRU_CO\
        );

    \I__2319\ : Odrv4
    port map (
            O => \N__13158\,
            I => \b2v_inst.un3_valor_max2_THRU_CO\
        );

    \I__2318\ : IoInMux
    port map (
            O => \N__13151\,
            I => \N__13148\
        );

    \I__2317\ : LocalMux
    port map (
            O => \N__13148\,
            I => \N__13145\
        );

    \I__2316\ : Span4Mux_s2_h
    port map (
            O => \N__13145\,
            I => \N__13142\
        );

    \I__2315\ : Sp12to4
    port map (
            O => \N__13142\,
            I => \N__13138\
        );

    \I__2314\ : InMux
    port map (
            O => \N__13141\,
            I => \N__13135\
        );

    \I__2313\ : Span12Mux_v
    port map (
            O => \N__13138\,
            I => \N__13130\
        );

    \I__2312\ : LocalMux
    port map (
            O => \N__13135\,
            I => \N__13130\
        );

    \I__2311\ : Odrv12
    port map (
            O => \N__13130\,
            I => reset_i
        );

    \I__2310\ : InMux
    port map (
            O => \N__13127\,
            I => \N__13124\
        );

    \I__2309\ : LocalMux
    port map (
            O => \N__13124\,
            I => \N__13121\
        );

    \I__2308\ : Span4Mux_v
    port map (
            O => \N__13121\,
            I => \N__13118\
        );

    \I__2307\ : Odrv4
    port map (
            O => \N__13118\,
            I => \b2v_inst3.un2_n_fsm_state_0_sqmuxa_2_0_i\
        );

    \I__2306\ : InMux
    port map (
            O => \N__13115\,
            I => \N__13112\
        );

    \I__2305\ : LocalMux
    port map (
            O => \N__13112\,
            I => \N__13109\
        );

    \I__2304\ : Span4Mux_h
    port map (
            O => \N__13109\,
            I => \N__13106\
        );

    \I__2303\ : Odrv4
    port map (
            O => \N__13106\,
            I => \b2v_inst1.r_RX_Bytece_0_6\
        );

    \I__2302\ : InMux
    port map (
            O => \N__13103\,
            I => \N__13099\
        );

    \I__2301\ : InMux
    port map (
            O => \N__13102\,
            I => \N__13096\
        );

    \I__2300\ : LocalMux
    port map (
            O => \N__13099\,
            I => \N__13092\
        );

    \I__2299\ : LocalMux
    port map (
            O => \N__13096\,
            I => \N__13089\
        );

    \I__2298\ : InMux
    port map (
            O => \N__13095\,
            I => \N__13086\
        );

    \I__2297\ : Span4Mux_h
    port map (
            O => \N__13092\,
            I => \N__13080\
        );

    \I__2296\ : Span4Mux_h
    port map (
            O => \N__13089\,
            I => \N__13080\
        );

    \I__2295\ : LocalMux
    port map (
            O => \N__13086\,
            I => \N__13077\
        );

    \I__2294\ : InMux
    port map (
            O => \N__13085\,
            I => \N__13074\
        );

    \I__2293\ : Odrv4
    port map (
            O => \N__13080\,
            I => \SYNTHESIZED_WIRE_1_0\
        );

    \I__2292\ : Odrv4
    port map (
            O => \N__13077\,
            I => \SYNTHESIZED_WIRE_1_0\
        );

    \I__2291\ : LocalMux
    port map (
            O => \N__13074\,
            I => \SYNTHESIZED_WIRE_1_0\
        );

    \I__2290\ : InMux
    port map (
            O => \N__13067\,
            I => \N__13064\
        );

    \I__2289\ : LocalMux
    port map (
            O => \N__13064\,
            I => \N__13061\
        );

    \I__2288\ : Span4Mux_v
    port map (
            O => \N__13061\,
            I => \N__13055\
        );

    \I__2287\ : InMux
    port map (
            O => \N__13060\,
            I => \N__13052\
        );

    \I__2286\ : InMux
    port map (
            O => \N__13059\,
            I => \N__13049\
        );

    \I__2285\ : InMux
    port map (
            O => \N__13058\,
            I => \N__13046\
        );

    \I__2284\ : Span4Mux_h
    port map (
            O => \N__13055\,
            I => \N__13041\
        );

    \I__2283\ : LocalMux
    port map (
            O => \N__13052\,
            I => \N__13041\
        );

    \I__2282\ : LocalMux
    port map (
            O => \N__13049\,
            I => \N__13038\
        );

    \I__2281\ : LocalMux
    port map (
            O => \N__13046\,
            I => \b2v_inst.reg_anteriorZ0Z_0\
        );

    \I__2280\ : Odrv4
    port map (
            O => \N__13041\,
            I => \b2v_inst.reg_anteriorZ0Z_0\
        );

    \I__2279\ : Odrv12
    port map (
            O => \N__13038\,
            I => \b2v_inst.reg_anteriorZ0Z_0\
        );

    \I__2278\ : InMux
    port map (
            O => \N__13031\,
            I => \N__13028\
        );

    \I__2277\ : LocalMux
    port map (
            O => \N__13028\,
            I => \N__13024\
        );

    \I__2276\ : InMux
    port map (
            O => \N__13027\,
            I => \N__13021\
        );

    \I__2275\ : Span4Mux_h
    port map (
            O => \N__13024\,
            I => \N__13017\
        );

    \I__2274\ : LocalMux
    port map (
            O => \N__13021\,
            I => \N__13014\
        );

    \I__2273\ : InMux
    port map (
            O => \N__13020\,
            I => \N__13011\
        );

    \I__2272\ : Span4Mux_v
    port map (
            O => \N__13017\,
            I => \N__13005\
        );

    \I__2271\ : Span4Mux_h
    port map (
            O => \N__13014\,
            I => \N__13005\
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__13011\,
            I => \N__13002\
        );

    \I__2269\ : InMux
    port map (
            O => \N__13010\,
            I => \N__12999\
        );

    \I__2268\ : Odrv4
    port map (
            O => \N__13005\,
            I => \SYNTHESIZED_WIRE_1_1\
        );

    \I__2267\ : Odrv4
    port map (
            O => \N__13002\,
            I => \SYNTHESIZED_WIRE_1_1\
        );

    \I__2266\ : LocalMux
    port map (
            O => \N__12999\,
            I => \SYNTHESIZED_WIRE_1_1\
        );

    \I__2265\ : InMux
    port map (
            O => \N__12992\,
            I => \N__12988\
        );

    \I__2264\ : InMux
    port map (
            O => \N__12991\,
            I => \N__12983\
        );

    \I__2263\ : LocalMux
    port map (
            O => \N__12988\,
            I => \N__12980\
        );

    \I__2262\ : InMux
    port map (
            O => \N__12987\,
            I => \N__12977\
        );

    \I__2261\ : InMux
    port map (
            O => \N__12986\,
            I => \N__12974\
        );

    \I__2260\ : LocalMux
    port map (
            O => \N__12983\,
            I => \N__12971\
        );

    \I__2259\ : Span4Mux_v
    port map (
            O => \N__12980\,
            I => \N__12966\
        );

    \I__2258\ : LocalMux
    port map (
            O => \N__12977\,
            I => \N__12966\
        );

    \I__2257\ : LocalMux
    port map (
            O => \N__12974\,
            I => \b2v_inst.reg_anteriorZ0Z_1\
        );

    \I__2256\ : Odrv4
    port map (
            O => \N__12971\,
            I => \b2v_inst.reg_anteriorZ0Z_1\
        );

    \I__2255\ : Odrv4
    port map (
            O => \N__12966\,
            I => \b2v_inst.reg_anteriorZ0Z_1\
        );

    \I__2254\ : InMux
    port map (
            O => \N__12959\,
            I => \N__12955\
        );

    \I__2253\ : InMux
    port map (
            O => \N__12958\,
            I => \N__12952\
        );

    \I__2252\ : LocalMux
    port map (
            O => \N__12955\,
            I => \N__12948\
        );

    \I__2251\ : LocalMux
    port map (
            O => \N__12952\,
            I => \N__12945\
        );

    \I__2250\ : InMux
    port map (
            O => \N__12951\,
            I => \N__12942\
        );

    \I__2249\ : Span4Mux_h
    port map (
            O => \N__12948\,
            I => \N__12936\
        );

    \I__2248\ : Span4Mux_h
    port map (
            O => \N__12945\,
            I => \N__12936\
        );

    \I__2247\ : LocalMux
    port map (
            O => \N__12942\,
            I => \N__12933\
        );

    \I__2246\ : InMux
    port map (
            O => \N__12941\,
            I => \N__12930\
        );

    \I__2245\ : Odrv4
    port map (
            O => \N__12936\,
            I => \SYNTHESIZED_WIRE_1_2\
        );

    \I__2244\ : Odrv12
    port map (
            O => \N__12933\,
            I => \SYNTHESIZED_WIRE_1_2\
        );

    \I__2243\ : LocalMux
    port map (
            O => \N__12930\,
            I => \SYNTHESIZED_WIRE_1_2\
        );

    \I__2242\ : CascadeMux
    port map (
            O => \N__12923\,
            I => \N__12920\
        );

    \I__2241\ : InMux
    port map (
            O => \N__12920\,
            I => \N__12916\
        );

    \I__2240\ : InMux
    port map (
            O => \N__12919\,
            I => \N__12911\
        );

    \I__2239\ : LocalMux
    port map (
            O => \N__12916\,
            I => \N__12908\
        );

    \I__2238\ : InMux
    port map (
            O => \N__12915\,
            I => \N__12905\
        );

    \I__2237\ : InMux
    port map (
            O => \N__12914\,
            I => \N__12902\
        );

    \I__2236\ : LocalMux
    port map (
            O => \N__12911\,
            I => \N__12899\
        );

    \I__2235\ : Span4Mux_v
    port map (
            O => \N__12908\,
            I => \N__12894\
        );

    \I__2234\ : LocalMux
    port map (
            O => \N__12905\,
            I => \N__12894\
        );

    \I__2233\ : LocalMux
    port map (
            O => \N__12902\,
            I => \b2v_inst.reg_anteriorZ0Z_2\
        );

    \I__2232\ : Odrv4
    port map (
            O => \N__12899\,
            I => \b2v_inst.reg_anteriorZ0Z_2\
        );

    \I__2231\ : Odrv4
    port map (
            O => \N__12894\,
            I => \b2v_inst.reg_anteriorZ0Z_2\
        );

    \I__2230\ : InMux
    port map (
            O => \N__12887\,
            I => \N__12883\
        );

    \I__2229\ : InMux
    port map (
            O => \N__12886\,
            I => \N__12880\
        );

    \I__2228\ : LocalMux
    port map (
            O => \N__12883\,
            I => \N__12876\
        );

    \I__2227\ : LocalMux
    port map (
            O => \N__12880\,
            I => \N__12873\
        );

    \I__2226\ : InMux
    port map (
            O => \N__12879\,
            I => \N__12870\
        );

    \I__2225\ : Span4Mux_h
    port map (
            O => \N__12876\,
            I => \N__12864\
        );

    \I__2224\ : Span4Mux_h
    port map (
            O => \N__12873\,
            I => \N__12864\
        );

    \I__2223\ : LocalMux
    port map (
            O => \N__12870\,
            I => \N__12861\
        );

    \I__2222\ : InMux
    port map (
            O => \N__12869\,
            I => \N__12858\
        );

    \I__2221\ : Odrv4
    port map (
            O => \N__12864\,
            I => \SYNTHESIZED_WIRE_1_3\
        );

    \I__2220\ : Odrv4
    port map (
            O => \N__12861\,
            I => \SYNTHESIZED_WIRE_1_3\
        );

    \I__2219\ : LocalMux
    port map (
            O => \N__12858\,
            I => \SYNTHESIZED_WIRE_1_3\
        );

    \I__2218\ : InMux
    port map (
            O => \N__12851\,
            I => \N__12848\
        );

    \I__2217\ : LocalMux
    port map (
            O => \N__12848\,
            I => \N__12842\
        );

    \I__2216\ : CascadeMux
    port map (
            O => \N__12847\,
            I => \N__12839\
        );

    \I__2215\ : InMux
    port map (
            O => \N__12846\,
            I => \N__12836\
        );

    \I__2214\ : InMux
    port map (
            O => \N__12845\,
            I => \N__12833\
        );

    \I__2213\ : Span4Mux_h
    port map (
            O => \N__12842\,
            I => \N__12830\
        );

    \I__2212\ : InMux
    port map (
            O => \N__12839\,
            I => \N__12827\
        );

    \I__2211\ : LocalMux
    port map (
            O => \N__12836\,
            I => \N__12824\
        );

    \I__2210\ : LocalMux
    port map (
            O => \N__12833\,
            I => \N__12821\
        );

    \I__2209\ : Odrv4
    port map (
            O => \N__12830\,
            I => \b2v_inst.reg_anteriorZ0Z_3\
        );

    \I__2208\ : LocalMux
    port map (
            O => \N__12827\,
            I => \b2v_inst.reg_anteriorZ0Z_3\
        );

    \I__2207\ : Odrv4
    port map (
            O => \N__12824\,
            I => \b2v_inst.reg_anteriorZ0Z_3\
        );

    \I__2206\ : Odrv4
    port map (
            O => \N__12821\,
            I => \b2v_inst.reg_anteriorZ0Z_3\
        );

    \I__2205\ : InMux
    port map (
            O => \N__12812\,
            I => \N__12809\
        );

    \I__2204\ : LocalMux
    port map (
            O => \N__12809\,
            I => \N__12804\
        );

    \I__2203\ : InMux
    port map (
            O => \N__12808\,
            I => \N__12801\
        );

    \I__2202\ : InMux
    port map (
            O => \N__12807\,
            I => \N__12798\
        );

    \I__2201\ : Odrv12
    port map (
            O => \N__12804\,
            I => \b2v_inst.reg_ancho_3Z0Z_6\
        );

    \I__2200\ : LocalMux
    port map (
            O => \N__12801\,
            I => \b2v_inst.reg_ancho_3Z0Z_6\
        );

    \I__2199\ : LocalMux
    port map (
            O => \N__12798\,
            I => \b2v_inst.reg_ancho_3Z0Z_6\
        );

    \I__2198\ : InMux
    port map (
            O => \N__12791\,
            I => \N__12788\
        );

    \I__2197\ : LocalMux
    port map (
            O => \N__12788\,
            I => \N__12785\
        );

    \I__2196\ : Span4Mux_h
    port map (
            O => \N__12785\,
            I => \N__12780\
        );

    \I__2195\ : InMux
    port map (
            O => \N__12784\,
            I => \N__12777\
        );

    \I__2194\ : InMux
    port map (
            O => \N__12783\,
            I => \N__12774\
        );

    \I__2193\ : Odrv4
    port map (
            O => \N__12780\,
            I => \b2v_inst.reg_ancho_3Z0Z_5\
        );

    \I__2192\ : LocalMux
    port map (
            O => \N__12777\,
            I => \b2v_inst.reg_ancho_3Z0Z_5\
        );

    \I__2191\ : LocalMux
    port map (
            O => \N__12774\,
            I => \b2v_inst.reg_ancho_3Z0Z_5\
        );

    \I__2190\ : CascadeMux
    port map (
            O => \N__12767\,
            I => \N__12764\
        );

    \I__2189\ : InMux
    port map (
            O => \N__12764\,
            I => \N__12759\
        );

    \I__2188\ : CascadeMux
    port map (
            O => \N__12763\,
            I => \N__12756\
        );

    \I__2187\ : CascadeMux
    port map (
            O => \N__12762\,
            I => \N__12753\
        );

    \I__2186\ : LocalMux
    port map (
            O => \N__12759\,
            I => \N__12750\
        );

    \I__2185\ : InMux
    port map (
            O => \N__12756\,
            I => \N__12747\
        );

    \I__2184\ : InMux
    port map (
            O => \N__12753\,
            I => \N__12744\
        );

    \I__2183\ : Odrv4
    port map (
            O => \N__12750\,
            I => \b2v_inst.reg_ancho_3_i_0\
        );

    \I__2182\ : LocalMux
    port map (
            O => \N__12747\,
            I => \b2v_inst.reg_ancho_3_i_0\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__12744\,
            I => \b2v_inst.reg_ancho_3_i_0\
        );

    \I__2180\ : CascadeMux
    port map (
            O => \N__12737\,
            I => \N__12732\
        );

    \I__2179\ : CascadeMux
    port map (
            O => \N__12736\,
            I => \N__12729\
        );

    \I__2178\ : CascadeMux
    port map (
            O => \N__12735\,
            I => \N__12726\
        );

    \I__2177\ : InMux
    port map (
            O => \N__12732\,
            I => \N__12723\
        );

    \I__2176\ : InMux
    port map (
            O => \N__12729\,
            I => \N__12720\
        );

    \I__2175\ : InMux
    port map (
            O => \N__12726\,
            I => \N__12717\
        );

    \I__2174\ : LocalMux
    port map (
            O => \N__12723\,
            I => \N__12714\
        );

    \I__2173\ : LocalMux
    port map (
            O => \N__12720\,
            I => \b2v_inst.reg_ancho_3_i_1\
        );

    \I__2172\ : LocalMux
    port map (
            O => \N__12717\,
            I => \b2v_inst.reg_ancho_3_i_1\
        );

    \I__2171\ : Odrv12
    port map (
            O => \N__12714\,
            I => \b2v_inst.reg_ancho_3_i_1\
        );

    \I__2170\ : CascadeMux
    port map (
            O => \N__12707\,
            I => \N__12704\
        );

    \I__2169\ : InMux
    port map (
            O => \N__12704\,
            I => \N__12699\
        );

    \I__2168\ : CascadeMux
    port map (
            O => \N__12703\,
            I => \N__12696\
        );

    \I__2167\ : CascadeMux
    port map (
            O => \N__12702\,
            I => \N__12693\
        );

    \I__2166\ : LocalMux
    port map (
            O => \N__12699\,
            I => \N__12690\
        );

    \I__2165\ : InMux
    port map (
            O => \N__12696\,
            I => \N__12687\
        );

    \I__2164\ : InMux
    port map (
            O => \N__12693\,
            I => \N__12684\
        );

    \I__2163\ : Odrv4
    port map (
            O => \N__12690\,
            I => \b2v_inst.reg_ancho_3_i_2\
        );

    \I__2162\ : LocalMux
    port map (
            O => \N__12687\,
            I => \b2v_inst.reg_ancho_3_i_2\
        );

    \I__2161\ : LocalMux
    port map (
            O => \N__12684\,
            I => \b2v_inst.reg_ancho_3_i_2\
        );

    \I__2160\ : CascadeMux
    port map (
            O => \N__12677\,
            I => \N__12672\
        );

    \I__2159\ : CascadeMux
    port map (
            O => \N__12676\,
            I => \N__12669\
        );

    \I__2158\ : CascadeMux
    port map (
            O => \N__12675\,
            I => \N__12666\
        );

    \I__2157\ : InMux
    port map (
            O => \N__12672\,
            I => \N__12663\
        );

    \I__2156\ : InMux
    port map (
            O => \N__12669\,
            I => \N__12660\
        );

    \I__2155\ : InMux
    port map (
            O => \N__12666\,
            I => \N__12657\
        );

    \I__2154\ : LocalMux
    port map (
            O => \N__12663\,
            I => \N__12654\
        );

    \I__2153\ : LocalMux
    port map (
            O => \N__12660\,
            I => \b2v_inst.reg_ancho_3_i_3\
        );

    \I__2152\ : LocalMux
    port map (
            O => \N__12657\,
            I => \b2v_inst.reg_ancho_3_i_3\
        );

    \I__2151\ : Odrv12
    port map (
            O => \N__12654\,
            I => \b2v_inst.reg_ancho_3_i_3\
        );

    \I__2150\ : CascadeMux
    port map (
            O => \N__12647\,
            I => \N__12644\
        );

    \I__2149\ : InMux
    port map (
            O => \N__12644\,
            I => \N__12639\
        );

    \I__2148\ : CascadeMux
    port map (
            O => \N__12643\,
            I => \N__12636\
        );

    \I__2147\ : CascadeMux
    port map (
            O => \N__12642\,
            I => \N__12633\
        );

    \I__2146\ : LocalMux
    port map (
            O => \N__12639\,
            I => \N__12630\
        );

    \I__2145\ : InMux
    port map (
            O => \N__12636\,
            I => \N__12627\
        );

    \I__2144\ : InMux
    port map (
            O => \N__12633\,
            I => \N__12624\
        );

    \I__2143\ : Odrv4
    port map (
            O => \N__12630\,
            I => \b2v_inst.reg_ancho_3_i_4\
        );

    \I__2142\ : LocalMux
    port map (
            O => \N__12627\,
            I => \b2v_inst.reg_ancho_3_i_4\
        );

    \I__2141\ : LocalMux
    port map (
            O => \N__12624\,
            I => \b2v_inst.reg_ancho_3_i_4\
        );

    \I__2140\ : CascadeMux
    port map (
            O => \N__12617\,
            I => \N__12614\
        );

    \I__2139\ : InMux
    port map (
            O => \N__12614\,
            I => \N__12609\
        );

    \I__2138\ : CascadeMux
    port map (
            O => \N__12613\,
            I => \N__12606\
        );

    \I__2137\ : CascadeMux
    port map (
            O => \N__12612\,
            I => \N__12603\
        );

    \I__2136\ : LocalMux
    port map (
            O => \N__12609\,
            I => \N__12600\
        );

    \I__2135\ : InMux
    port map (
            O => \N__12606\,
            I => \N__12597\
        );

    \I__2134\ : InMux
    port map (
            O => \N__12603\,
            I => \N__12594\
        );

    \I__2133\ : Odrv4
    port map (
            O => \N__12600\,
            I => \b2v_inst.reg_ancho_3_i_5\
        );

    \I__2132\ : LocalMux
    port map (
            O => \N__12597\,
            I => \b2v_inst.reg_ancho_3_i_5\
        );

    \I__2131\ : LocalMux
    port map (
            O => \N__12594\,
            I => \b2v_inst.reg_ancho_3_i_5\
        );

    \I__2130\ : CascadeMux
    port map (
            O => \N__12587\,
            I => \N__12584\
        );

    \I__2129\ : InMux
    port map (
            O => \N__12584\,
            I => \N__12579\
        );

    \I__2128\ : CascadeMux
    port map (
            O => \N__12583\,
            I => \N__12576\
        );

    \I__2127\ : CascadeMux
    port map (
            O => \N__12582\,
            I => \N__12573\
        );

    \I__2126\ : LocalMux
    port map (
            O => \N__12579\,
            I => \N__12570\
        );

    \I__2125\ : InMux
    port map (
            O => \N__12576\,
            I => \N__12567\
        );

    \I__2124\ : InMux
    port map (
            O => \N__12573\,
            I => \N__12564\
        );

    \I__2123\ : Odrv4
    port map (
            O => \N__12570\,
            I => \b2v_inst.reg_ancho_3_i_6\
        );

    \I__2122\ : LocalMux
    port map (
            O => \N__12567\,
            I => \b2v_inst.reg_ancho_3_i_6\
        );

    \I__2121\ : LocalMux
    port map (
            O => \N__12564\,
            I => \b2v_inst.reg_ancho_3_i_6\
        );

    \I__2120\ : InMux
    port map (
            O => \N__12557\,
            I => \N__12553\
        );

    \I__2119\ : InMux
    port map (
            O => \N__12556\,
            I => \N__12550\
        );

    \I__2118\ : LocalMux
    port map (
            O => \N__12553\,
            I => \SYNTHESIZED_WIRE_10_7\
        );

    \I__2117\ : LocalMux
    port map (
            O => \N__12550\,
            I => \SYNTHESIZED_WIRE_10_7\
        );

    \I__2116\ : CascadeMux
    port map (
            O => \N__12545\,
            I => \b2v_inst.addr_ram_1_iv_i_2_5_cascade_\
        );

    \I__2115\ : CascadeMux
    port map (
            O => \N__12542\,
            I => \N__12538\
        );

    \I__2114\ : CascadeMux
    port map (
            O => \N__12541\,
            I => \N__12535\
        );

    \I__2113\ : InMux
    port map (
            O => \N__12538\,
            I => \N__12532\
        );

    \I__2112\ : InMux
    port map (
            O => \N__12535\,
            I => \N__12529\
        );

    \I__2111\ : LocalMux
    port map (
            O => \N__12532\,
            I => \N__12526\
        );

    \I__2110\ : LocalMux
    port map (
            O => \N__12529\,
            I => \N__12523\
        );

    \I__2109\ : Span4Mux_h
    port map (
            O => \N__12526\,
            I => \N__12520\
        );

    \I__2108\ : Odrv4
    port map (
            O => \N__12523\,
            I => \N_54\
        );

    \I__2107\ : Odrv4
    port map (
            O => \N__12520\,
            I => \N_54\
        );

    \I__2106\ : InMux
    port map (
            O => \N__12515\,
            I => \N__12512\
        );

    \I__2105\ : LocalMux
    port map (
            O => \N__12512\,
            I => \b2v_inst.addr_ram_1_iv_i_1_5\
        );

    \I__2104\ : InMux
    port map (
            O => \N__12509\,
            I => \N__12506\
        );

    \I__2103\ : LocalMux
    port map (
            O => \N__12506\,
            I => \b2v_inst.N_341\
        );

    \I__2102\ : CascadeMux
    port map (
            O => \N__12503\,
            I => \b2v_inst.N_404_cascade_\
        );

    \I__2101\ : InMux
    port map (
            O => \N__12500\,
            I => \N__12487\
        );

    \I__2100\ : InMux
    port map (
            O => \N__12499\,
            I => \N__12487\
        );

    \I__2099\ : InMux
    port map (
            O => \N__12498\,
            I => \N__12474\
        );

    \I__2098\ : InMux
    port map (
            O => \N__12497\,
            I => \N__12474\
        );

    \I__2097\ : InMux
    port map (
            O => \N__12496\,
            I => \N__12474\
        );

    \I__2096\ : InMux
    port map (
            O => \N__12495\,
            I => \N__12474\
        );

    \I__2095\ : InMux
    port map (
            O => \N__12494\,
            I => \N__12474\
        );

    \I__2094\ : InMux
    port map (
            O => \N__12493\,
            I => \N__12474\
        );

    \I__2093\ : InMux
    port map (
            O => \N__12492\,
            I => \N__12470\
        );

    \I__2092\ : LocalMux
    port map (
            O => \N__12487\,
            I => \N__12467\
        );

    \I__2091\ : LocalMux
    port map (
            O => \N__12474\,
            I => \N__12464\
        );

    \I__2090\ : InMux
    port map (
            O => \N__12473\,
            I => \N__12461\
        );

    \I__2089\ : LocalMux
    port map (
            O => \N__12470\,
            I => \b2v_inst.cuenta_pixelZ0Z_0\
        );

    \I__2088\ : Odrv12
    port map (
            O => \N__12467\,
            I => \b2v_inst.cuenta_pixelZ0Z_0\
        );

    \I__2087\ : Odrv4
    port map (
            O => \N__12464\,
            I => \b2v_inst.cuenta_pixelZ0Z_0\
        );

    \I__2086\ : LocalMux
    port map (
            O => \N__12461\,
            I => \b2v_inst.cuenta_pixelZ0Z_0\
        );

    \I__2085\ : CascadeMux
    port map (
            O => \N__12452\,
            I => \N__12449\
        );

    \I__2084\ : InMux
    port map (
            O => \N__12449\,
            I => \N__12443\
        );

    \I__2083\ : InMux
    port map (
            O => \N__12448\,
            I => \N__12443\
        );

    \I__2082\ : LocalMux
    port map (
            O => \N__12443\,
            I => \N__12440\
        );

    \I__2081\ : Span4Mux_h
    port map (
            O => \N__12440\,
            I => \N__12434\
        );

    \I__2080\ : CascadeMux
    port map (
            O => \N__12439\,
            I => \N__12431\
        );

    \I__2079\ : CascadeMux
    port map (
            O => \N__12438\,
            I => \N__12428\
        );

    \I__2078\ : CascadeMux
    port map (
            O => \N__12437\,
            I => \N__12423\
        );

    \I__2077\ : Span4Mux_h
    port map (
            O => \N__12434\,
            I => \N__12418\
        );

    \I__2076\ : InMux
    port map (
            O => \N__12431\,
            I => \N__12405\
        );

    \I__2075\ : InMux
    port map (
            O => \N__12428\,
            I => \N__12405\
        );

    \I__2074\ : InMux
    port map (
            O => \N__12427\,
            I => \N__12405\
        );

    \I__2073\ : InMux
    port map (
            O => \N__12426\,
            I => \N__12405\
        );

    \I__2072\ : InMux
    port map (
            O => \N__12423\,
            I => \N__12405\
        );

    \I__2071\ : InMux
    port map (
            O => \N__12422\,
            I => \N__12405\
        );

    \I__2070\ : InMux
    port map (
            O => \N__12421\,
            I => \N__12402\
        );

    \I__2069\ : Odrv4
    port map (
            O => \N__12418\,
            I => \b2v_inst.cuenta_pixelZ0Z_1\
        );

    \I__2068\ : LocalMux
    port map (
            O => \N__12405\,
            I => \b2v_inst.cuenta_pixelZ0Z_1\
        );

    \I__2067\ : LocalMux
    port map (
            O => \N__12402\,
            I => \b2v_inst.cuenta_pixelZ0Z_1\
        );

    \I__2066\ : InMux
    port map (
            O => \N__12395\,
            I => \N__12392\
        );

    \I__2065\ : LocalMux
    port map (
            O => \N__12392\,
            I => \N__12389\
        );

    \I__2064\ : Odrv12
    port map (
            O => \N__12389\,
            I => \b2v_inst.cuenta_pixel_4_i_a2_0_6\
        );

    \I__2063\ : InMux
    port map (
            O => \N__12386\,
            I => \N__12383\
        );

    \I__2062\ : LocalMux
    port map (
            O => \N__12383\,
            I => \N__12380\
        );

    \I__2061\ : Span4Mux_h
    port map (
            O => \N__12380\,
            I => \N__12377\
        );

    \I__2060\ : Odrv4
    port map (
            O => \N__12377\,
            I => \N_213_i\
        );

    \I__2059\ : InMux
    port map (
            O => \N__12374\,
            I => \N__12371\
        );

    \I__2058\ : LocalMux
    port map (
            O => \N__12371\,
            I => \N__12368\
        );

    \I__2057\ : Span4Mux_h
    port map (
            O => \N__12368\,
            I => \N__12365\
        );

    \I__2056\ : Odrv4
    port map (
            O => \N__12365\,
            I => \N_209_i\
        );

    \I__2055\ : InMux
    port map (
            O => \N__12362\,
            I => \N__12359\
        );

    \I__2054\ : LocalMux
    port map (
            O => \N__12359\,
            I => \N__12356\
        );

    \I__2053\ : Span4Mux_h
    port map (
            O => \N__12356\,
            I => \N__12353\
        );

    \I__2052\ : Odrv4
    port map (
            O => \N__12353\,
            I => \N_207_i\
        );

    \I__2051\ : InMux
    port map (
            O => \N__12350\,
            I => \N__12346\
        );

    \I__2050\ : InMux
    port map (
            O => \N__12349\,
            I => \N__12343\
        );

    \I__2049\ : LocalMux
    port map (
            O => \N__12346\,
            I => \SYNTHESIZED_WIRE_10_2\
        );

    \I__2048\ : LocalMux
    port map (
            O => \N__12343\,
            I => \SYNTHESIZED_WIRE_10_2\
        );

    \I__2047\ : InMux
    port map (
            O => \N__12338\,
            I => \N__12334\
        );

    \I__2046\ : InMux
    port map (
            O => \N__12337\,
            I => \N__12331\
        );

    \I__2045\ : LocalMux
    port map (
            O => \N__12334\,
            I => \SYNTHESIZED_WIRE_10_3\
        );

    \I__2044\ : LocalMux
    port map (
            O => \N__12331\,
            I => \SYNTHESIZED_WIRE_10_3\
        );

    \I__2043\ : InMux
    port map (
            O => \N__12326\,
            I => \N__12322\
        );

    \I__2042\ : InMux
    port map (
            O => \N__12325\,
            I => \N__12319\
        );

    \I__2041\ : LocalMux
    port map (
            O => \N__12322\,
            I => \SYNTHESIZED_WIRE_10_4\
        );

    \I__2040\ : LocalMux
    port map (
            O => \N__12319\,
            I => \SYNTHESIZED_WIRE_10_4\
        );

    \I__2039\ : InMux
    port map (
            O => \N__12314\,
            I => \N__12310\
        );

    \I__2038\ : InMux
    port map (
            O => \N__12313\,
            I => \N__12307\
        );

    \I__2037\ : LocalMux
    port map (
            O => \N__12310\,
            I => \SYNTHESIZED_WIRE_10_5\
        );

    \I__2036\ : LocalMux
    port map (
            O => \N__12307\,
            I => \SYNTHESIZED_WIRE_10_5\
        );

    \I__2035\ : CascadeMux
    port map (
            O => \N__12302\,
            I => \N__12298\
        );

    \I__2034\ : InMux
    port map (
            O => \N__12301\,
            I => \N__12295\
        );

    \I__2033\ : InMux
    port map (
            O => \N__12298\,
            I => \N__12292\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__12295\,
            I => \SYNTHESIZED_WIRE_10_6\
        );

    \I__2031\ : LocalMux
    port map (
            O => \N__12292\,
            I => \SYNTHESIZED_WIRE_10_6\
        );

    \I__2030\ : CascadeMux
    port map (
            O => \N__12287\,
            I => \b2v_inst3.next_bit_0_a3_4_cascade_\
        );

    \I__2029\ : InMux
    port map (
            O => \N__12284\,
            I => \N__12281\
        );

    \I__2028\ : LocalMux
    port map (
            O => \N__12281\,
            I => \b2v_inst3.next_bit_0_a3_3\
        );

    \I__2027\ : CascadeMux
    port map (
            O => \N__12278\,
            I => \N__12273\
        );

    \I__2026\ : InMux
    port map (
            O => \N__12277\,
            I => \N__12266\
        );

    \I__2025\ : InMux
    port map (
            O => \N__12276\,
            I => \N__12266\
        );

    \I__2024\ : InMux
    port map (
            O => \N__12273\,
            I => \N__12266\
        );

    \I__2023\ : LocalMux
    port map (
            O => \N__12266\,
            I => \N__12261\
        );

    \I__2022\ : InMux
    port map (
            O => \N__12265\,
            I => \N__12258\
        );

    \I__2021\ : InMux
    port map (
            O => \N__12264\,
            I => \N__12255\
        );

    \I__2020\ : Span4Mux_v
    port map (
            O => \N__12261\,
            I => \N__12252\
        );

    \I__2019\ : LocalMux
    port map (
            O => \N__12258\,
            I => \SYNTHESIZED_WIRE_7\
        );

    \I__2018\ : LocalMux
    port map (
            O => \N__12255\,
            I => \SYNTHESIZED_WIRE_7\
        );

    \I__2017\ : Odrv4
    port map (
            O => \N__12252\,
            I => \SYNTHESIZED_WIRE_7\
        );

    \I__2016\ : CascadeMux
    port map (
            O => \N__12245\,
            I => \b2v_inst3.N_105_7_cascade_\
        );

    \I__2015\ : InMux
    port map (
            O => \N__12242\,
            I => \N__12238\
        );

    \I__2014\ : InMux
    port map (
            O => \N__12241\,
            I => \N__12229\
        );

    \I__2013\ : LocalMux
    port map (
            O => \N__12238\,
            I => \N__12226\
        );

    \I__2012\ : InMux
    port map (
            O => \N__12237\,
            I => \N__12221\
        );

    \I__2011\ : InMux
    port map (
            O => \N__12236\,
            I => \N__12221\
        );

    \I__2010\ : InMux
    port map (
            O => \N__12235\,
            I => \N__12216\
        );

    \I__2009\ : InMux
    port map (
            O => \N__12234\,
            I => \N__12216\
        );

    \I__2008\ : InMux
    port map (
            O => \N__12233\,
            I => \N__12211\
        );

    \I__2007\ : InMux
    port map (
            O => \N__12232\,
            I => \N__12211\
        );

    \I__2006\ : LocalMux
    port map (
            O => \N__12229\,
            I => \b2v_inst3.fsm_stateZ0Z_0\
        );

    \I__2005\ : Odrv4
    port map (
            O => \N__12226\,
            I => \b2v_inst3.fsm_stateZ0Z_0\
        );

    \I__2004\ : LocalMux
    port map (
            O => \N__12221\,
            I => \b2v_inst3.fsm_stateZ0Z_0\
        );

    \I__2003\ : LocalMux
    port map (
            O => \N__12216\,
            I => \b2v_inst3.fsm_stateZ0Z_0\
        );

    \I__2002\ : LocalMux
    port map (
            O => \N__12211\,
            I => \b2v_inst3.fsm_stateZ0Z_0\
        );

    \I__2001\ : CascadeMux
    port map (
            O => \N__12200\,
            I => \N__12195\
        );

    \I__2000\ : InMux
    port map (
            O => \N__12199\,
            I => \N__12188\
        );

    \I__1999\ : InMux
    port map (
            O => \N__12198\,
            I => \N__12188\
        );

    \I__1998\ : InMux
    port map (
            O => \N__12195\,
            I => \N__12181\
        );

    \I__1997\ : InMux
    port map (
            O => \N__12194\,
            I => \N__12181\
        );

    \I__1996\ : InMux
    port map (
            O => \N__12193\,
            I => \N__12181\
        );

    \I__1995\ : LocalMux
    port map (
            O => \N__12188\,
            I => \b2v_inst3.cycle_counterZ0Z_1\
        );

    \I__1994\ : LocalMux
    port map (
            O => \N__12181\,
            I => \b2v_inst3.cycle_counterZ0Z_1\
        );

    \I__1993\ : CascadeMux
    port map (
            O => \N__12176\,
            I => \N__12173\
        );

    \I__1992\ : InMux
    port map (
            O => \N__12173\,
            I => \N__12167\
        );

    \I__1991\ : InMux
    port map (
            O => \N__12172\,
            I => \N__12167\
        );

    \I__1990\ : LocalMux
    port map (
            O => \N__12167\,
            I => \N__12162\
        );

    \I__1989\ : CascadeMux
    port map (
            O => \N__12166\,
            I => \N__12154\
        );

    \I__1988\ : InMux
    port map (
            O => \N__12165\,
            I => \N__12150\
        );

    \I__1987\ : Span4Mux_h
    port map (
            O => \N__12162\,
            I => \N__12147\
        );

    \I__1986\ : InMux
    port map (
            O => \N__12161\,
            I => \N__12142\
        );

    \I__1985\ : InMux
    port map (
            O => \N__12160\,
            I => \N__12142\
        );

    \I__1984\ : InMux
    port map (
            O => \N__12159\,
            I => \N__12135\
        );

    \I__1983\ : InMux
    port map (
            O => \N__12158\,
            I => \N__12135\
        );

    \I__1982\ : InMux
    port map (
            O => \N__12157\,
            I => \N__12135\
        );

    \I__1981\ : InMux
    port map (
            O => \N__12154\,
            I => \N__12130\
        );

    \I__1980\ : InMux
    port map (
            O => \N__12153\,
            I => \N__12130\
        );

    \I__1979\ : LocalMux
    port map (
            O => \N__12150\,
            I => \b2v_inst3.fsm_stateZ0Z_1\
        );

    \I__1978\ : Odrv4
    port map (
            O => \N__12147\,
            I => \b2v_inst3.fsm_stateZ0Z_1\
        );

    \I__1977\ : LocalMux
    port map (
            O => \N__12142\,
            I => \b2v_inst3.fsm_stateZ0Z_1\
        );

    \I__1976\ : LocalMux
    port map (
            O => \N__12135\,
            I => \b2v_inst3.fsm_stateZ0Z_1\
        );

    \I__1975\ : LocalMux
    port map (
            O => \N__12130\,
            I => \b2v_inst3.fsm_stateZ0Z_1\
        );

    \I__1974\ : InMux
    port map (
            O => \N__12119\,
            I => \N__12109\
        );

    \I__1973\ : InMux
    port map (
            O => \N__12118\,
            I => \N__12109\
        );

    \I__1972\ : InMux
    port map (
            O => \N__12117\,
            I => \N__12100\
        );

    \I__1971\ : InMux
    port map (
            O => \N__12116\,
            I => \N__12100\
        );

    \I__1970\ : InMux
    port map (
            O => \N__12115\,
            I => \N__12100\
        );

    \I__1969\ : InMux
    port map (
            O => \N__12114\,
            I => \N__12100\
        );

    \I__1968\ : LocalMux
    port map (
            O => \N__12109\,
            I => \b2v_inst3.cycle_counterZ0Z_0\
        );

    \I__1967\ : LocalMux
    port map (
            O => \N__12100\,
            I => \b2v_inst3.cycle_counterZ0Z_0\
        );

    \I__1966\ : InMux
    port map (
            O => \N__12095\,
            I => \N__12092\
        );

    \I__1965\ : LocalMux
    port map (
            O => \N__12092\,
            I => \b2v_inst3.un1_cycle_counter_5_c2\
        );

    \I__1964\ : CascadeMux
    port map (
            O => \N__12089\,
            I => \N__12085\
        );

    \I__1963\ : CascadeMux
    port map (
            O => \N__12088\,
            I => \N__12082\
        );

    \I__1962\ : InMux
    port map (
            O => \N__12085\,
            I => \N__12076\
        );

    \I__1961\ : InMux
    port map (
            O => \N__12082\,
            I => \N__12071\
        );

    \I__1960\ : InMux
    port map (
            O => \N__12081\,
            I => \N__12071\
        );

    \I__1959\ : InMux
    port map (
            O => \N__12080\,
            I => \N__12066\
        );

    \I__1958\ : InMux
    port map (
            O => \N__12079\,
            I => \N__12066\
        );

    \I__1957\ : LocalMux
    port map (
            O => \N__12076\,
            I => \b2v_inst3.cycle_counterZ0Z_2\
        );

    \I__1956\ : LocalMux
    port map (
            O => \N__12071\,
            I => \b2v_inst3.cycle_counterZ0Z_2\
        );

    \I__1955\ : LocalMux
    port map (
            O => \N__12066\,
            I => \b2v_inst3.cycle_counterZ0Z_2\
        );

    \I__1954\ : InMux
    port map (
            O => \N__12059\,
            I => \N__12053\
        );

    \I__1953\ : InMux
    port map (
            O => \N__12058\,
            I => \N__12050\
        );

    \I__1952\ : InMux
    port map (
            O => \N__12057\,
            I => \N__12045\
        );

    \I__1951\ : InMux
    port map (
            O => \N__12056\,
            I => \N__12045\
        );

    \I__1950\ : LocalMux
    port map (
            O => \N__12053\,
            I => \b2v_inst3.cycle_counterZ0Z_3\
        );

    \I__1949\ : LocalMux
    port map (
            O => \N__12050\,
            I => \b2v_inst3.cycle_counterZ0Z_3\
        );

    \I__1948\ : LocalMux
    port map (
            O => \N__12045\,
            I => \b2v_inst3.cycle_counterZ0Z_3\
        );

    \I__1947\ : CascadeMux
    port map (
            O => \N__12038\,
            I => \b2v_inst3.un1_cycle_counter_5_c2_cascade_\
        );

    \I__1946\ : InMux
    port map (
            O => \N__12035\,
            I => \N__12030\
        );

    \I__1945\ : InMux
    port map (
            O => \N__12034\,
            I => \N__12025\
        );

    \I__1944\ : InMux
    port map (
            O => \N__12033\,
            I => \N__12025\
        );

    \I__1943\ : LocalMux
    port map (
            O => \N__12030\,
            I => \b2v_inst3.cycle_counterZ0Z_4\
        );

    \I__1942\ : LocalMux
    port map (
            O => \N__12025\,
            I => \b2v_inst3.cycle_counterZ0Z_4\
        );

    \I__1941\ : InMux
    port map (
            O => \N__12020\,
            I => \N__12017\
        );

    \I__1940\ : LocalMux
    port map (
            O => \N__12017\,
            I => \N__12014\
        );

    \I__1939\ : Span4Mux_h
    port map (
            O => \N__12014\,
            I => \N__12004\
        );

    \I__1938\ : InMux
    port map (
            O => \N__12013\,
            I => \N__11989\
        );

    \I__1937\ : InMux
    port map (
            O => \N__12012\,
            I => \N__11989\
        );

    \I__1936\ : InMux
    port map (
            O => \N__12011\,
            I => \N__11989\
        );

    \I__1935\ : InMux
    port map (
            O => \N__12010\,
            I => \N__11989\
        );

    \I__1934\ : InMux
    port map (
            O => \N__12009\,
            I => \N__11989\
        );

    \I__1933\ : InMux
    port map (
            O => \N__12008\,
            I => \N__11989\
        );

    \I__1932\ : InMux
    port map (
            O => \N__12007\,
            I => \N__11989\
        );

    \I__1931\ : Odrv4
    port map (
            O => \N__12004\,
            I => \b2v_inst4.un1_pix_count_int_0_sqmuxa_9\
        );

    \I__1930\ : LocalMux
    port map (
            O => \N__11989\,
            I => \b2v_inst4.un1_pix_count_int_0_sqmuxa_9\
        );

    \I__1929\ : InMux
    port map (
            O => \N__11984\,
            I => \N__11981\
        );

    \I__1928\ : LocalMux
    port map (
            O => \N__11981\,
            I => \N__11978\
        );

    \I__1927\ : Span4Mux_v
    port map (
            O => \N__11978\,
            I => \N__11968\
        );

    \I__1926\ : InMux
    port map (
            O => \N__11977\,
            I => \N__11953\
        );

    \I__1925\ : InMux
    port map (
            O => \N__11976\,
            I => \N__11953\
        );

    \I__1924\ : InMux
    port map (
            O => \N__11975\,
            I => \N__11953\
        );

    \I__1923\ : InMux
    port map (
            O => \N__11974\,
            I => \N__11953\
        );

    \I__1922\ : InMux
    port map (
            O => \N__11973\,
            I => \N__11953\
        );

    \I__1921\ : InMux
    port map (
            O => \N__11972\,
            I => \N__11953\
        );

    \I__1920\ : InMux
    port map (
            O => \N__11971\,
            I => \N__11953\
        );

    \I__1919\ : Odrv4
    port map (
            O => \N__11968\,
            I => \b2v_inst4.un1_pix_count_int_0_sqmuxa_11\
        );

    \I__1918\ : LocalMux
    port map (
            O => \N__11953\,
            I => \b2v_inst4.un1_pix_count_int_0_sqmuxa_11\
        );

    \I__1917\ : CascadeMux
    port map (
            O => \N__11948\,
            I => \N__11941\
        );

    \I__1916\ : CascadeMux
    port map (
            O => \N__11947\,
            I => \N__11938\
        );

    \I__1915\ : CascadeMux
    port map (
            O => \N__11946\,
            I => \N__11935\
        );

    \I__1914\ : CascadeMux
    port map (
            O => \N__11945\,
            I => \N__11932\
        );

    \I__1913\ : CascadeMux
    port map (
            O => \N__11944\,
            I => \N__11929\
        );

    \I__1912\ : InMux
    port map (
            O => \N__11941\,
            I => \N__11926\
        );

    \I__1911\ : InMux
    port map (
            O => \N__11938\,
            I => \N__11914\
        );

    \I__1910\ : InMux
    port map (
            O => \N__11935\,
            I => \N__11914\
        );

    \I__1909\ : InMux
    port map (
            O => \N__11932\,
            I => \N__11914\
        );

    \I__1908\ : InMux
    port map (
            O => \N__11929\,
            I => \N__11914\
        );

    \I__1907\ : LocalMux
    port map (
            O => \N__11926\,
            I => \N__11911\
        );

    \I__1906\ : CascadeMux
    port map (
            O => \N__11925\,
            I => \N__11908\
        );

    \I__1905\ : CascadeMux
    port map (
            O => \N__11924\,
            I => \N__11905\
        );

    \I__1904\ : CascadeMux
    port map (
            O => \N__11923\,
            I => \N__11902\
        );

    \I__1903\ : LocalMux
    port map (
            O => \N__11914\,
            I => \N__11897\
        );

    \I__1902\ : Span4Mux_h
    port map (
            O => \N__11911\,
            I => \N__11897\
        );

    \I__1901\ : InMux
    port map (
            O => \N__11908\,
            I => \N__11890\
        );

    \I__1900\ : InMux
    port map (
            O => \N__11905\,
            I => \N__11890\
        );

    \I__1899\ : InMux
    port map (
            O => \N__11902\,
            I => \N__11890\
        );

    \I__1898\ : Span4Mux_h
    port map (
            O => \N__11897\,
            I => \N__11887\
        );

    \I__1897\ : LocalMux
    port map (
            O => \N__11890\,
            I => \b2v_inst4.un1_pix_count_int_0_sqmuxa_10\
        );

    \I__1896\ : Odrv4
    port map (
            O => \N__11887\,
            I => \b2v_inst4.un1_pix_count_int_0_sqmuxa_10\
        );

    \I__1895\ : InMux
    port map (
            O => \N__11882\,
            I => \N__11879\
        );

    \I__1894\ : LocalMux
    port map (
            O => \N__11879\,
            I => \N__11876\
        );

    \I__1893\ : Span4Mux_v
    port map (
            O => \N__11876\,
            I => \N__11873\
        );

    \I__1892\ : Odrv4
    port map (
            O => \N__11873\,
            I => \b2v_inst4.pix_count_int_RNO_0Z0Z_9\
        );

    \I__1891\ : InMux
    port map (
            O => \N__11870\,
            I => \N__11864\
        );

    \I__1890\ : InMux
    port map (
            O => \N__11869\,
            I => \N__11857\
        );

    \I__1889\ : InMux
    port map (
            O => \N__11868\,
            I => \N__11857\
        );

    \I__1888\ : InMux
    port map (
            O => \N__11867\,
            I => \N__11857\
        );

    \I__1887\ : LocalMux
    port map (
            O => \N__11864\,
            I => \N__11852\
        );

    \I__1886\ : LocalMux
    port map (
            O => \N__11857\,
            I => \N__11852\
        );

    \I__1885\ : Span4Mux_h
    port map (
            O => \N__11852\,
            I => \N__11849\
        );

    \I__1884\ : Odrv4
    port map (
            O => \N__11849\,
            I => \SYNTHESIZED_WIRE_2_9\
        );

    \I__1883\ : CascadeMux
    port map (
            O => \N__11846\,
            I => \N__11841\
        );

    \I__1882\ : CascadeMux
    port map (
            O => \N__11845\,
            I => \N__11838\
        );

    \I__1881\ : InMux
    port map (
            O => \N__11844\,
            I => \N__11835\
        );

    \I__1880\ : InMux
    port map (
            O => \N__11841\,
            I => \N__11829\
        );

    \I__1879\ : InMux
    port map (
            O => \N__11838\,
            I => \N__11826\
        );

    \I__1878\ : LocalMux
    port map (
            O => \N__11835\,
            I => \N__11823\
        );

    \I__1877\ : InMux
    port map (
            O => \N__11834\,
            I => \N__11816\
        );

    \I__1876\ : InMux
    port map (
            O => \N__11833\,
            I => \N__11816\
        );

    \I__1875\ : InMux
    port map (
            O => \N__11832\,
            I => \N__11816\
        );

    \I__1874\ : LocalMux
    port map (
            O => \N__11829\,
            I => \N__11813\
        );

    \I__1873\ : LocalMux
    port map (
            O => \N__11826\,
            I => \N__11810\
        );

    \I__1872\ : Odrv12
    port map (
            O => \N__11823\,
            I => \b2v_inst.cuenta_pixelZ0Z_6\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__11816\,
            I => \b2v_inst.cuenta_pixelZ0Z_6\
        );

    \I__1870\ : Odrv4
    port map (
            O => \N__11813\,
            I => \b2v_inst.cuenta_pixelZ0Z_6\
        );

    \I__1869\ : Odrv4
    port map (
            O => \N__11810\,
            I => \b2v_inst.cuenta_pixelZ0Z_6\
        );

    \I__1868\ : CascadeMux
    port map (
            O => \N__11801\,
            I => \N__11798\
        );

    \I__1867\ : InMux
    port map (
            O => \N__11798\,
            I => \N__11795\
        );

    \I__1866\ : LocalMux
    port map (
            O => \N__11795\,
            I => \N__11791\
        );

    \I__1865\ : CascadeMux
    port map (
            O => \N__11794\,
            I => \N__11788\
        );

    \I__1864\ : Span4Mux_v
    port map (
            O => \N__11791\,
            I => \N__11784\
        );

    \I__1863\ : InMux
    port map (
            O => \N__11788\,
            I => \N__11779\
        );

    \I__1862\ : InMux
    port map (
            O => \N__11787\,
            I => \N__11779\
        );

    \I__1861\ : Span4Mux_h
    port map (
            O => \N__11784\,
            I => \N__11776\
        );

    \I__1860\ : LocalMux
    port map (
            O => \N__11779\,
            I => \N__11773\
        );

    \I__1859\ : Odrv4
    port map (
            O => \N__11776\,
            I => \b2v_inst.un11_cuenta_pixel_i_0_o2_0\
        );

    \I__1858\ : Odrv12
    port map (
            O => \N__11773\,
            I => \b2v_inst.un11_cuenta_pixel_i_0_o2_0\
        );

    \I__1857\ : InMux
    port map (
            O => \N__11768\,
            I => \N__11765\
        );

    \I__1856\ : LocalMux
    port map (
            O => \N__11765\,
            I => \N__11761\
        );

    \I__1855\ : CascadeMux
    port map (
            O => \N__11764\,
            I => \N__11756\
        );

    \I__1854\ : Span4Mux_h
    port map (
            O => \N__11761\,
            I => \N__11752\
        );

    \I__1853\ : InMux
    port map (
            O => \N__11760\,
            I => \N__11747\
        );

    \I__1852\ : InMux
    port map (
            O => \N__11759\,
            I => \N__11747\
        );

    \I__1851\ : InMux
    port map (
            O => \N__11756\,
            I => \N__11742\
        );

    \I__1850\ : InMux
    port map (
            O => \N__11755\,
            I => \N__11742\
        );

    \I__1849\ : Odrv4
    port map (
            O => \N__11752\,
            I => \b2v_inst.cuenta_pixelZ0Z_5\
        );

    \I__1848\ : LocalMux
    port map (
            O => \N__11747\,
            I => \b2v_inst.cuenta_pixelZ0Z_5\
        );

    \I__1847\ : LocalMux
    port map (
            O => \N__11742\,
            I => \b2v_inst.cuenta_pixelZ0Z_5\
        );

    \I__1846\ : IoInMux
    port map (
            O => \N__11735\,
            I => \N__11732\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__11732\,
            I => \N__11729\
        );

    \I__1844\ : Span4Mux_s3_v
    port map (
            O => \N__11729\,
            I => \N__11726\
        );

    \I__1843\ : Sp12to4
    port map (
            O => \N__11726\,
            I => \N__11723\
        );

    \I__1842\ : Span12Mux_h
    port map (
            O => \N__11723\,
            I => \N__11720\
        );

    \I__1841\ : Span12Mux_v
    port map (
            O => \N__11720\,
            I => \N__11717\
        );

    \I__1840\ : Odrv12
    port map (
            O => \N__11717\,
            I => uart_tx_o
        );

    \I__1839\ : InMux
    port map (
            O => \N__11714\,
            I => \N__11710\
        );

    \I__1838\ : InMux
    port map (
            O => \N__11713\,
            I => \N__11707\
        );

    \I__1837\ : LocalMux
    port map (
            O => \N__11710\,
            I => \N__11701\
        );

    \I__1836\ : LocalMux
    port map (
            O => \N__11707\,
            I => \N__11701\
        );

    \I__1835\ : InMux
    port map (
            O => \N__11706\,
            I => \N__11698\
        );

    \I__1834\ : Span4Mux_v
    port map (
            O => \N__11701\,
            I => \N__11695\
        );

    \I__1833\ : LocalMux
    port map (
            O => \N__11698\,
            I => \b2v_inst4.stateZ0Z_0\
        );

    \I__1832\ : Odrv4
    port map (
            O => \N__11695\,
            I => \b2v_inst4.stateZ0Z_0\
        );

    \I__1831\ : InMux
    port map (
            O => \N__11690\,
            I => \N__11683\
        );

    \I__1830\ : InMux
    port map (
            O => \N__11689\,
            I => \N__11683\
        );

    \I__1829\ : InMux
    port map (
            O => \N__11688\,
            I => \N__11680\
        );

    \I__1828\ : LocalMux
    port map (
            O => \N__11683\,
            I => \N__11675\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__11680\,
            I => \N__11675\
        );

    \I__1826\ : Odrv4
    port map (
            O => \N__11675\,
            I => \b2v_inst3.cycle_counterZ0Z_6\
        );

    \I__1825\ : InMux
    port map (
            O => \N__11672\,
            I => \N__11662\
        );

    \I__1824\ : InMux
    port map (
            O => \N__11671\,
            I => \N__11662\
        );

    \I__1823\ : InMux
    port map (
            O => \N__11670\,
            I => \N__11662\
        );

    \I__1822\ : InMux
    port map (
            O => \N__11669\,
            I => \N__11659\
        );

    \I__1821\ : LocalMux
    port map (
            O => \N__11662\,
            I => \b2v_inst3.cycle_counterZ0Z_5\
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__11659\,
            I => \b2v_inst3.cycle_counterZ0Z_5\
        );

    \I__1819\ : CascadeMux
    port map (
            O => \N__11654\,
            I => \N__11650\
        );

    \I__1818\ : InMux
    port map (
            O => \N__11653\,
            I => \N__11647\
        );

    \I__1817\ : InMux
    port map (
            O => \N__11650\,
            I => \N__11644\
        );

    \I__1816\ : LocalMux
    port map (
            O => \N__11647\,
            I => \b2v_inst3.cycle_counterZ0Z_7\
        );

    \I__1815\ : LocalMux
    port map (
            O => \N__11644\,
            I => \b2v_inst3.cycle_counterZ0Z_7\
        );

    \I__1814\ : InMux
    port map (
            O => \N__11639\,
            I => \bfn_5_20_0_\
        );

    \I__1813\ : CascadeMux
    port map (
            O => \N__11636\,
            I => \N__11632\
        );

    \I__1812\ : InMux
    port map (
            O => \N__11635\,
            I => \N__11629\
        );

    \I__1811\ : InMux
    port map (
            O => \N__11632\,
            I => \N__11626\
        );

    \I__1810\ : LocalMux
    port map (
            O => \N__11629\,
            I => \N__11623\
        );

    \I__1809\ : LocalMux
    port map (
            O => \N__11626\,
            I => \N__11620\
        );

    \I__1808\ : Span4Mux_v
    port map (
            O => \N__11623\,
            I => \N__11617\
        );

    \I__1807\ : Span4Mux_h
    port map (
            O => \N__11620\,
            I => \N__11614\
        );

    \I__1806\ : Odrv4
    port map (
            O => \N__11617\,
            I => \b2v_inst.valor_max_final52_THRU_CO\
        );

    \I__1805\ : Odrv4
    port map (
            O => \N__11614\,
            I => \b2v_inst.valor_max_final52_THRU_CO\
        );

    \I__1804\ : InMux
    port map (
            O => \N__11609\,
            I => \N__11606\
        );

    \I__1803\ : LocalMux
    port map (
            O => \N__11606\,
            I => \b2v_inst3.un1_bit_counter_3_c2\
        );

    \I__1802\ : CascadeMux
    port map (
            O => \N__11603\,
            I => \b2v_inst3.un1_bit_counter_3_c2_cascade_\
        );

    \I__1801\ : InMux
    port map (
            O => \N__11600\,
            I => \N__11597\
        );

    \I__1800\ : LocalMux
    port map (
            O => \N__11597\,
            I => \b2v_inst3.N_258\
        );

    \I__1799\ : CascadeMux
    port map (
            O => \N__11594\,
            I => \b2v_inst3.N_258_cascade_\
        );

    \I__1798\ : InMux
    port map (
            O => \N__11591\,
            I => \N__11583\
        );

    \I__1797\ : InMux
    port map (
            O => \N__11590\,
            I => \N__11583\
        );

    \I__1796\ : InMux
    port map (
            O => \N__11589\,
            I => \N__11578\
        );

    \I__1795\ : InMux
    port map (
            O => \N__11588\,
            I => \N__11578\
        );

    \I__1794\ : LocalMux
    port map (
            O => \N__11583\,
            I => \b2v_inst3.bit_counterZ0Z_2\
        );

    \I__1793\ : LocalMux
    port map (
            O => \N__11578\,
            I => \b2v_inst3.bit_counterZ0Z_2\
        );

    \I__1792\ : InMux
    port map (
            O => \N__11573\,
            I => \N__11565\
        );

    \I__1791\ : InMux
    port map (
            O => \N__11572\,
            I => \N__11565\
        );

    \I__1790\ : InMux
    port map (
            O => \N__11571\,
            I => \N__11560\
        );

    \I__1789\ : InMux
    port map (
            O => \N__11570\,
            I => \N__11560\
        );

    \I__1788\ : LocalMux
    port map (
            O => \N__11565\,
            I => \b2v_inst3.bit_counterZ1Z_1\
        );

    \I__1787\ : LocalMux
    port map (
            O => \N__11560\,
            I => \b2v_inst3.bit_counterZ1Z_1\
        );

    \I__1786\ : CascadeMux
    port map (
            O => \N__11555\,
            I => \b2v_inst3.N_102_2_cascade_\
        );

    \I__1785\ : CascadeMux
    port map (
            O => \N__11552\,
            I => \N__11547\
        );

    \I__1784\ : InMux
    port map (
            O => \N__11551\,
            I => \N__11540\
        );

    \I__1783\ : InMux
    port map (
            O => \N__11550\,
            I => \N__11540\
        );

    \I__1782\ : InMux
    port map (
            O => \N__11547\,
            I => \N__11540\
        );

    \I__1781\ : LocalMux
    port map (
            O => \N__11540\,
            I => \b2v_inst3.bit_counterZ0Z_3\
        );

    \I__1780\ : InMux
    port map (
            O => \N__11537\,
            I => \N__11533\
        );

    \I__1779\ : InMux
    port map (
            O => \N__11536\,
            I => \N__11530\
        );

    \I__1778\ : LocalMux
    port map (
            O => \N__11533\,
            I => \b2v_inst3.N_436\
        );

    \I__1777\ : LocalMux
    port map (
            O => \N__11530\,
            I => \b2v_inst3.N_436\
        );

    \I__1776\ : InMux
    port map (
            O => \N__11525\,
            I => \N__11522\
        );

    \I__1775\ : LocalMux
    port map (
            O => \N__11522\,
            I => \N__11519\
        );

    \I__1774\ : Span4Mux_h
    port map (
            O => \N__11519\,
            I => \N__11516\
        );

    \I__1773\ : Odrv4
    port map (
            O => \N__11516\,
            I => \b2v_inst.data_a_escribir9_6_and\
        );

    \I__1772\ : CascadeMux
    port map (
            O => \N__11513\,
            I => \N__11507\
        );

    \I__1771\ : InMux
    port map (
            O => \N__11512\,
            I => \N__11503\
        );

    \I__1770\ : InMux
    port map (
            O => \N__11511\,
            I => \N__11500\
        );

    \I__1769\ : InMux
    port map (
            O => \N__11510\,
            I => \N__11497\
        );

    \I__1768\ : InMux
    port map (
            O => \N__11507\,
            I => \N__11494\
        );

    \I__1767\ : InMux
    port map (
            O => \N__11506\,
            I => \N__11491\
        );

    \I__1766\ : LocalMux
    port map (
            O => \N__11503\,
            I => \N__11488\
        );

    \I__1765\ : LocalMux
    port map (
            O => \N__11500\,
            I => \N__11485\
        );

    \I__1764\ : LocalMux
    port map (
            O => \N__11497\,
            I => \b2v_inst.reg_ancho_2Z0Z_0\
        );

    \I__1763\ : LocalMux
    port map (
            O => \N__11494\,
            I => \b2v_inst.reg_ancho_2Z0Z_0\
        );

    \I__1762\ : LocalMux
    port map (
            O => \N__11491\,
            I => \b2v_inst.reg_ancho_2Z0Z_0\
        );

    \I__1761\ : Odrv4
    port map (
            O => \N__11488\,
            I => \b2v_inst.reg_ancho_2Z0Z_0\
        );

    \I__1760\ : Odrv4
    port map (
            O => \N__11485\,
            I => \b2v_inst.reg_ancho_2Z0Z_0\
        );

    \I__1759\ : InMux
    port map (
            O => \N__11474\,
            I => \N__11468\
        );

    \I__1758\ : InMux
    port map (
            O => \N__11473\,
            I => \N__11465\
        );

    \I__1757\ : InMux
    port map (
            O => \N__11472\,
            I => \N__11462\
        );

    \I__1756\ : CascadeMux
    port map (
            O => \N__11471\,
            I => \N__11459\
        );

    \I__1755\ : LocalMux
    port map (
            O => \N__11468\,
            I => \N__11455\
        );

    \I__1754\ : LocalMux
    port map (
            O => \N__11465\,
            I => \N__11452\
        );

    \I__1753\ : LocalMux
    port map (
            O => \N__11462\,
            I => \N__11449\
        );

    \I__1752\ : InMux
    port map (
            O => \N__11459\,
            I => \N__11446\
        );

    \I__1751\ : InMux
    port map (
            O => \N__11458\,
            I => \N__11443\
        );

    \I__1750\ : Span4Mux_h
    port map (
            O => \N__11455\,
            I => \N__11438\
        );

    \I__1749\ : Span4Mux_v
    port map (
            O => \N__11452\,
            I => \N__11438\
        );

    \I__1748\ : Odrv4
    port map (
            O => \N__11449\,
            I => \b2v_inst.reg_ancho_2Z0Z_1\
        );

    \I__1747\ : LocalMux
    port map (
            O => \N__11446\,
            I => \b2v_inst.reg_ancho_2Z0Z_1\
        );

    \I__1746\ : LocalMux
    port map (
            O => \N__11443\,
            I => \b2v_inst.reg_ancho_2Z0Z_1\
        );

    \I__1745\ : Odrv4
    port map (
            O => \N__11438\,
            I => \b2v_inst.reg_ancho_2Z0Z_1\
        );

    \I__1744\ : CascadeMux
    port map (
            O => \N__11429\,
            I => \N__11423\
        );

    \I__1743\ : InMux
    port map (
            O => \N__11428\,
            I => \N__11420\
        );

    \I__1742\ : InMux
    port map (
            O => \N__11427\,
            I => \N__11416\
        );

    \I__1741\ : InMux
    port map (
            O => \N__11426\,
            I => \N__11413\
        );

    \I__1740\ : InMux
    port map (
            O => \N__11423\,
            I => \N__11410\
        );

    \I__1739\ : LocalMux
    port map (
            O => \N__11420\,
            I => \N__11407\
        );

    \I__1738\ : InMux
    port map (
            O => \N__11419\,
            I => \N__11404\
        );

    \I__1737\ : LocalMux
    port map (
            O => \N__11416\,
            I => \N__11401\
        );

    \I__1736\ : LocalMux
    port map (
            O => \N__11413\,
            I => \b2v_inst.reg_ancho_2Z0Z_2\
        );

    \I__1735\ : LocalMux
    port map (
            O => \N__11410\,
            I => \b2v_inst.reg_ancho_2Z0Z_2\
        );

    \I__1734\ : Odrv4
    port map (
            O => \N__11407\,
            I => \b2v_inst.reg_ancho_2Z0Z_2\
        );

    \I__1733\ : LocalMux
    port map (
            O => \N__11404\,
            I => \b2v_inst.reg_ancho_2Z0Z_2\
        );

    \I__1732\ : Odrv4
    port map (
            O => \N__11401\,
            I => \b2v_inst.reg_ancho_2Z0Z_2\
        );

    \I__1731\ : CascadeMux
    port map (
            O => \N__11390\,
            I => \N__11383\
        );

    \I__1730\ : CascadeMux
    port map (
            O => \N__11389\,
            I => \N__11380\
        );

    \I__1729\ : InMux
    port map (
            O => \N__11388\,
            I => \N__11377\
        );

    \I__1728\ : CascadeMux
    port map (
            O => \N__11387\,
            I => \N__11374\
        );

    \I__1727\ : InMux
    port map (
            O => \N__11386\,
            I => \N__11371\
        );

    \I__1726\ : InMux
    port map (
            O => \N__11383\,
            I => \N__11368\
        );

    \I__1725\ : InMux
    port map (
            O => \N__11380\,
            I => \N__11365\
        );

    \I__1724\ : LocalMux
    port map (
            O => \N__11377\,
            I => \N__11362\
        );

    \I__1723\ : InMux
    port map (
            O => \N__11374\,
            I => \N__11359\
        );

    \I__1722\ : LocalMux
    port map (
            O => \N__11371\,
            I => \N__11356\
        );

    \I__1721\ : LocalMux
    port map (
            O => \N__11368\,
            I => \b2v_inst.reg_ancho_2Z0Z_3\
        );

    \I__1720\ : LocalMux
    port map (
            O => \N__11365\,
            I => \b2v_inst.reg_ancho_2Z0Z_3\
        );

    \I__1719\ : Odrv4
    port map (
            O => \N__11362\,
            I => \b2v_inst.reg_ancho_2Z0Z_3\
        );

    \I__1718\ : LocalMux
    port map (
            O => \N__11359\,
            I => \b2v_inst.reg_ancho_2Z0Z_3\
        );

    \I__1717\ : Odrv4
    port map (
            O => \N__11356\,
            I => \b2v_inst.reg_ancho_2Z0Z_3\
        );

    \I__1716\ : InMux
    port map (
            O => \N__11345\,
            I => \N__11341\
        );

    \I__1715\ : InMux
    port map (
            O => \N__11344\,
            I => \N__11338\
        );

    \I__1714\ : LocalMux
    port map (
            O => \N__11341\,
            I => \N__11334\
        );

    \I__1713\ : LocalMux
    port map (
            O => \N__11338\,
            I => \N__11331\
        );

    \I__1712\ : InMux
    port map (
            O => \N__11337\,
            I => \N__11328\
        );

    \I__1711\ : Span4Mux_v
    port map (
            O => \N__11334\,
            I => \N__11319\
        );

    \I__1710\ : Span4Mux_v
    port map (
            O => \N__11331\,
            I => \N__11319\
        );

    \I__1709\ : LocalMux
    port map (
            O => \N__11328\,
            I => \N__11319\
        );

    \I__1708\ : InMux
    port map (
            O => \N__11327\,
            I => \N__11314\
        );

    \I__1707\ : InMux
    port map (
            O => \N__11326\,
            I => \N__11314\
        );

    \I__1706\ : Odrv4
    port map (
            O => \N__11319\,
            I => \b2v_inst.reg_ancho_2Z0Z_4\
        );

    \I__1705\ : LocalMux
    port map (
            O => \N__11314\,
            I => \b2v_inst.reg_ancho_2Z0Z_4\
        );

    \I__1704\ : InMux
    port map (
            O => \N__11309\,
            I => \N__11305\
        );

    \I__1703\ : InMux
    port map (
            O => \N__11308\,
            I => \N__11300\
        );

    \I__1702\ : LocalMux
    port map (
            O => \N__11305\,
            I => \N__11297\
        );

    \I__1701\ : InMux
    port map (
            O => \N__11304\,
            I => \N__11294\
        );

    \I__1700\ : InMux
    port map (
            O => \N__11303\,
            I => \N__11290\
        );

    \I__1699\ : LocalMux
    port map (
            O => \N__11300\,
            I => \N__11287\
        );

    \I__1698\ : Span4Mux_v
    port map (
            O => \N__11297\,
            I => \N__11284\
        );

    \I__1697\ : LocalMux
    port map (
            O => \N__11294\,
            I => \N__11281\
        );

    \I__1696\ : InMux
    port map (
            O => \N__11293\,
            I => \N__11278\
        );

    \I__1695\ : LocalMux
    port map (
            O => \N__11290\,
            I => \b2v_inst.reg_ancho_2Z0Z_5\
        );

    \I__1694\ : Odrv4
    port map (
            O => \N__11287\,
            I => \b2v_inst.reg_ancho_2Z0Z_5\
        );

    \I__1693\ : Odrv4
    port map (
            O => \N__11284\,
            I => \b2v_inst.reg_ancho_2Z0Z_5\
        );

    \I__1692\ : Odrv12
    port map (
            O => \N__11281\,
            I => \b2v_inst.reg_ancho_2Z0Z_5\
        );

    \I__1691\ : LocalMux
    port map (
            O => \N__11278\,
            I => \b2v_inst.reg_ancho_2Z0Z_5\
        );

    \I__1690\ : CascadeMux
    port map (
            O => \N__11267\,
            I => \N__11264\
        );

    \I__1689\ : InMux
    port map (
            O => \N__11264\,
            I => \N__11259\
        );

    \I__1688\ : InMux
    port map (
            O => \N__11263\,
            I => \N__11256\
        );

    \I__1687\ : InMux
    port map (
            O => \N__11262\,
            I => \N__11253\
        );

    \I__1686\ : LocalMux
    port map (
            O => \N__11259\,
            I => \N__11250\
        );

    \I__1685\ : LocalMux
    port map (
            O => \N__11256\,
            I => \N__11247\
        );

    \I__1684\ : LocalMux
    port map (
            O => \N__11253\,
            I => \N__11244\
        );

    \I__1683\ : Span4Mux_v
    port map (
            O => \N__11250\,
            I => \N__11235\
        );

    \I__1682\ : Span4Mux_v
    port map (
            O => \N__11247\,
            I => \N__11235\
        );

    \I__1681\ : Span4Mux_v
    port map (
            O => \N__11244\,
            I => \N__11235\
        );

    \I__1680\ : InMux
    port map (
            O => \N__11243\,
            I => \N__11232\
        );

    \I__1679\ : InMux
    port map (
            O => \N__11242\,
            I => \N__11229\
        );

    \I__1678\ : Odrv4
    port map (
            O => \N__11235\,
            I => \b2v_inst.reg_ancho_2Z0Z_6\
        );

    \I__1677\ : LocalMux
    port map (
            O => \N__11232\,
            I => \b2v_inst.reg_ancho_2Z0Z_6\
        );

    \I__1676\ : LocalMux
    port map (
            O => \N__11229\,
            I => \b2v_inst.reg_ancho_2Z0Z_6\
        );

    \I__1675\ : CascadeMux
    port map (
            O => \N__11222\,
            I => \N__11218\
        );

    \I__1674\ : InMux
    port map (
            O => \N__11221\,
            I => \N__11214\
        );

    \I__1673\ : InMux
    port map (
            O => \N__11218\,
            I => \N__11210\
        );

    \I__1672\ : CascadeMux
    port map (
            O => \N__11217\,
            I => \N__11207\
        );

    \I__1671\ : LocalMux
    port map (
            O => \N__11214\,
            I => \N__11204\
        );

    \I__1670\ : InMux
    port map (
            O => \N__11213\,
            I => \N__11200\
        );

    \I__1669\ : LocalMux
    port map (
            O => \N__11210\,
            I => \N__11197\
        );

    \I__1668\ : InMux
    port map (
            O => \N__11207\,
            I => \N__11194\
        );

    \I__1667\ : Span4Mux_v
    port map (
            O => \N__11204\,
            I => \N__11191\
        );

    \I__1666\ : CascadeMux
    port map (
            O => \N__11203\,
            I => \N__11188\
        );

    \I__1665\ : LocalMux
    port map (
            O => \N__11200\,
            I => \N__11185\
        );

    \I__1664\ : Span4Mux_h
    port map (
            O => \N__11197\,
            I => \N__11178\
        );

    \I__1663\ : LocalMux
    port map (
            O => \N__11194\,
            I => \N__11178\
        );

    \I__1662\ : Span4Mux_h
    port map (
            O => \N__11191\,
            I => \N__11178\
        );

    \I__1661\ : InMux
    port map (
            O => \N__11188\,
            I => \N__11175\
        );

    \I__1660\ : Odrv4
    port map (
            O => \N__11185\,
            I => \b2v_inst.reg_ancho_2Z0Z_7\
        );

    \I__1659\ : Odrv4
    port map (
            O => \N__11178\,
            I => \b2v_inst.reg_ancho_2Z0Z_7\
        );

    \I__1658\ : LocalMux
    port map (
            O => \N__11175\,
            I => \b2v_inst.reg_ancho_2Z0Z_7\
        );

    \I__1657\ : InMux
    port map (
            O => \N__11168\,
            I => \N__11164\
        );

    \I__1656\ : InMux
    port map (
            O => \N__11167\,
            I => \N__11160\
        );

    \I__1655\ : LocalMux
    port map (
            O => \N__11164\,
            I => \N__11157\
        );

    \I__1654\ : InMux
    port map (
            O => \N__11163\,
            I => \N__11152\
        );

    \I__1653\ : LocalMux
    port map (
            O => \N__11160\,
            I => \N__11149\
        );

    \I__1652\ : Span4Mux_h
    port map (
            O => \N__11157\,
            I => \N__11146\
        );

    \I__1651\ : InMux
    port map (
            O => \N__11156\,
            I => \N__11143\
        );

    \I__1650\ : InMux
    port map (
            O => \N__11155\,
            I => \N__11140\
        );

    \I__1649\ : LocalMux
    port map (
            O => \N__11152\,
            I => \b2v_inst.reg_ancho_1Z0Z_1\
        );

    \I__1648\ : Odrv4
    port map (
            O => \N__11149\,
            I => \b2v_inst.reg_ancho_1Z0Z_1\
        );

    \I__1647\ : Odrv4
    port map (
            O => \N__11146\,
            I => \b2v_inst.reg_ancho_1Z0Z_1\
        );

    \I__1646\ : LocalMux
    port map (
            O => \N__11143\,
            I => \b2v_inst.reg_ancho_1Z0Z_1\
        );

    \I__1645\ : LocalMux
    port map (
            O => \N__11140\,
            I => \b2v_inst.reg_ancho_1Z0Z_1\
        );

    \I__1644\ : InMux
    port map (
            O => \N__11129\,
            I => \N__11126\
        );

    \I__1643\ : LocalMux
    port map (
            O => \N__11126\,
            I => \N__11122\
        );

    \I__1642\ : InMux
    port map (
            O => \N__11125\,
            I => \N__11118\
        );

    \I__1641\ : Span4Mux_v
    port map (
            O => \N__11122\,
            I => \N__11115\
        );

    \I__1640\ : InMux
    port map (
            O => \N__11121\,
            I => \N__11112\
        );

    \I__1639\ : LocalMux
    port map (
            O => \N__11118\,
            I => \N__11109\
        );

    \I__1638\ : Odrv4
    port map (
            O => \N__11115\,
            I => \b2v_inst.reg_ancho_3Z0Z_1\
        );

    \I__1637\ : LocalMux
    port map (
            O => \N__11112\,
            I => \b2v_inst.reg_ancho_3Z0Z_1\
        );

    \I__1636\ : Odrv4
    port map (
            O => \N__11109\,
            I => \b2v_inst.reg_ancho_3Z0Z_1\
        );

    \I__1635\ : InMux
    port map (
            O => \N__11102\,
            I => \N__11099\
        );

    \I__1634\ : LocalMux
    port map (
            O => \N__11099\,
            I => \N__11095\
        );

    \I__1633\ : InMux
    port map (
            O => \N__11098\,
            I => \N__11091\
        );

    \I__1632\ : Span4Mux_h
    port map (
            O => \N__11095\,
            I => \N__11088\
        );

    \I__1631\ : InMux
    port map (
            O => \N__11094\,
            I => \N__11085\
        );

    \I__1630\ : LocalMux
    port map (
            O => \N__11091\,
            I => \N__11082\
        );

    \I__1629\ : Odrv4
    port map (
            O => \N__11088\,
            I => \b2v_inst.reg_ancho_3Z0Z_2\
        );

    \I__1628\ : LocalMux
    port map (
            O => \N__11085\,
            I => \b2v_inst.reg_ancho_3Z0Z_2\
        );

    \I__1627\ : Odrv12
    port map (
            O => \N__11082\,
            I => \b2v_inst.reg_ancho_3Z0Z_2\
        );

    \I__1626\ : CascadeMux
    port map (
            O => \N__11075\,
            I => \N__11071\
        );

    \I__1625\ : InMux
    port map (
            O => \N__11074\,
            I => \N__11067\
        );

    \I__1624\ : InMux
    port map (
            O => \N__11071\,
            I => \N__11064\
        );

    \I__1623\ : InMux
    port map (
            O => \N__11070\,
            I => \N__11061\
        );

    \I__1622\ : LocalMux
    port map (
            O => \N__11067\,
            I => \N__11057\
        );

    \I__1621\ : LocalMux
    port map (
            O => \N__11064\,
            I => \N__11051\
        );

    \I__1620\ : LocalMux
    port map (
            O => \N__11061\,
            I => \N__11051\
        );

    \I__1619\ : InMux
    port map (
            O => \N__11060\,
            I => \N__11048\
        );

    \I__1618\ : Span4Mux_h
    port map (
            O => \N__11057\,
            I => \N__11045\
        );

    \I__1617\ : InMux
    port map (
            O => \N__11056\,
            I => \N__11042\
        );

    \I__1616\ : Odrv4
    port map (
            O => \N__11051\,
            I => \b2v_inst.reg_ancho_1Z0Z_2\
        );

    \I__1615\ : LocalMux
    port map (
            O => \N__11048\,
            I => \b2v_inst.reg_ancho_1Z0Z_2\
        );

    \I__1614\ : Odrv4
    port map (
            O => \N__11045\,
            I => \b2v_inst.reg_ancho_1Z0Z_2\
        );

    \I__1613\ : LocalMux
    port map (
            O => \N__11042\,
            I => \b2v_inst.reg_ancho_1Z0Z_2\
        );

    \I__1612\ : InMux
    port map (
            O => \N__11033\,
            I => \N__11029\
        );

    \I__1611\ : InMux
    port map (
            O => \N__11032\,
            I => \N__11026\
        );

    \I__1610\ : LocalMux
    port map (
            O => \N__11029\,
            I => \N__11023\
        );

    \I__1609\ : LocalMux
    port map (
            O => \N__11026\,
            I => \N__11018\
        );

    \I__1608\ : Span4Mux_v
    port map (
            O => \N__11023\,
            I => \N__11015\
        );

    \I__1607\ : CascadeMux
    port map (
            O => \N__11022\,
            I => \N__11012\
        );

    \I__1606\ : InMux
    port map (
            O => \N__11021\,
            I => \N__11008\
        );

    \I__1605\ : Span4Mux_h
    port map (
            O => \N__11018\,
            I => \N__11003\
        );

    \I__1604\ : Span4Mux_h
    port map (
            O => \N__11015\,
            I => \N__11003\
        );

    \I__1603\ : InMux
    port map (
            O => \N__11012\,
            I => \N__11000\
        );

    \I__1602\ : InMux
    port map (
            O => \N__11011\,
            I => \N__10997\
        );

    \I__1601\ : LocalMux
    port map (
            O => \N__11008\,
            I => \b2v_inst.reg_ancho_1Z0Z_3\
        );

    \I__1600\ : Odrv4
    port map (
            O => \N__11003\,
            I => \b2v_inst.reg_ancho_1Z0Z_3\
        );

    \I__1599\ : LocalMux
    port map (
            O => \N__11000\,
            I => \b2v_inst.reg_ancho_1Z0Z_3\
        );

    \I__1598\ : LocalMux
    port map (
            O => \N__10997\,
            I => \b2v_inst.reg_ancho_1Z0Z_3\
        );

    \I__1597\ : InMux
    port map (
            O => \N__10988\,
            I => \N__10985\
        );

    \I__1596\ : LocalMux
    port map (
            O => \N__10985\,
            I => \N__10981\
        );

    \I__1595\ : CascadeMux
    port map (
            O => \N__10984\,
            I => \N__10977\
        );

    \I__1594\ : Span4Mux_v
    port map (
            O => \N__10981\,
            I => \N__10974\
        );

    \I__1593\ : InMux
    port map (
            O => \N__10980\,
            I => \N__10971\
        );

    \I__1592\ : InMux
    port map (
            O => \N__10977\,
            I => \N__10968\
        );

    \I__1591\ : Span4Mux_h
    port map (
            O => \N__10974\,
            I => \N__10963\
        );

    \I__1590\ : LocalMux
    port map (
            O => \N__10971\,
            I => \N__10963\
        );

    \I__1589\ : LocalMux
    port map (
            O => \N__10968\,
            I => \b2v_inst.reg_ancho_3Z0Z_3\
        );

    \I__1588\ : Odrv4
    port map (
            O => \N__10963\,
            I => \b2v_inst.reg_ancho_3Z0Z_3\
        );

    \I__1587\ : InMux
    port map (
            O => \N__10958\,
            I => \N__10955\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__10955\,
            I => \N__10951\
        );

    \I__1585\ : InMux
    port map (
            O => \N__10954\,
            I => \N__10947\
        );

    \I__1584\ : Span4Mux_v
    port map (
            O => \N__10951\,
            I => \N__10943\
        );

    \I__1583\ : InMux
    port map (
            O => \N__10950\,
            I => \N__10939\
        );

    \I__1582\ : LocalMux
    port map (
            O => \N__10947\,
            I => \N__10936\
        );

    \I__1581\ : InMux
    port map (
            O => \N__10946\,
            I => \N__10933\
        );

    \I__1580\ : Span4Mux_h
    port map (
            O => \N__10943\,
            I => \N__10930\
        );

    \I__1579\ : InMux
    port map (
            O => \N__10942\,
            I => \N__10927\
        );

    \I__1578\ : LocalMux
    port map (
            O => \N__10939\,
            I => \b2v_inst.reg_ancho_1Z0Z_4\
        );

    \I__1577\ : Odrv4
    port map (
            O => \N__10936\,
            I => \b2v_inst.reg_ancho_1Z0Z_4\
        );

    \I__1576\ : LocalMux
    port map (
            O => \N__10933\,
            I => \b2v_inst.reg_ancho_1Z0Z_4\
        );

    \I__1575\ : Odrv4
    port map (
            O => \N__10930\,
            I => \b2v_inst.reg_ancho_1Z0Z_4\
        );

    \I__1574\ : LocalMux
    port map (
            O => \N__10927\,
            I => \b2v_inst.reg_ancho_1Z0Z_4\
        );

    \I__1573\ : InMux
    port map (
            O => \N__10916\,
            I => \N__10913\
        );

    \I__1572\ : LocalMux
    port map (
            O => \N__10913\,
            I => \N__10910\
        );

    \I__1571\ : Span4Mux_h
    port map (
            O => \N__10910\,
            I => \N__10906\
        );

    \I__1570\ : InMux
    port map (
            O => \N__10909\,
            I => \N__10902\
        );

    \I__1569\ : Span4Mux_v
    port map (
            O => \N__10906\,
            I => \N__10899\
        );

    \I__1568\ : InMux
    port map (
            O => \N__10905\,
            I => \N__10896\
        );

    \I__1567\ : LocalMux
    port map (
            O => \N__10902\,
            I => \N__10893\
        );

    \I__1566\ : Odrv4
    port map (
            O => \N__10899\,
            I => \b2v_inst.reg_ancho_3Z0Z_4\
        );

    \I__1565\ : LocalMux
    port map (
            O => \N__10896\,
            I => \b2v_inst.reg_ancho_3Z0Z_4\
        );

    \I__1564\ : Odrv4
    port map (
            O => \N__10893\,
            I => \b2v_inst.reg_ancho_3Z0Z_4\
        );

    \I__1563\ : InMux
    port map (
            O => \N__10886\,
            I => \N__10881\
        );

    \I__1562\ : InMux
    port map (
            O => \N__10885\,
            I => \N__10878\
        );

    \I__1561\ : InMux
    port map (
            O => \N__10884\,
            I => \N__10875\
        );

    \I__1560\ : LocalMux
    port map (
            O => \N__10881\,
            I => \N__10872\
        );

    \I__1559\ : LocalMux
    port map (
            O => \N__10878\,
            I => \N__10865\
        );

    \I__1558\ : LocalMux
    port map (
            O => \N__10875\,
            I => \N__10865\
        );

    \I__1557\ : Span4Mux_h
    port map (
            O => \N__10872\,
            I => \N__10862\
        );

    \I__1556\ : InMux
    port map (
            O => \N__10871\,
            I => \N__10859\
        );

    \I__1555\ : InMux
    port map (
            O => \N__10870\,
            I => \N__10856\
        );

    \I__1554\ : Odrv4
    port map (
            O => \N__10865\,
            I => \b2v_inst.reg_ancho_1Z0Z_5\
        );

    \I__1553\ : Odrv4
    port map (
            O => \N__10862\,
            I => \b2v_inst.reg_ancho_1Z0Z_5\
        );

    \I__1552\ : LocalMux
    port map (
            O => \N__10859\,
            I => \b2v_inst.reg_ancho_1Z0Z_5\
        );

    \I__1551\ : LocalMux
    port map (
            O => \N__10856\,
            I => \b2v_inst.reg_ancho_1Z0Z_5\
        );

    \I__1550\ : InMux
    port map (
            O => \N__10847\,
            I => \N__10842\
        );

    \I__1549\ : InMux
    port map (
            O => \N__10846\,
            I => \N__10839\
        );

    \I__1548\ : InMux
    port map (
            O => \N__10845\,
            I => \N__10836\
        );

    \I__1547\ : LocalMux
    port map (
            O => \N__10842\,
            I => \N__10833\
        );

    \I__1546\ : LocalMux
    port map (
            O => \N__10839\,
            I => \N__10830\
        );

    \I__1545\ : LocalMux
    port map (
            O => \N__10836\,
            I => \N__10825\
        );

    \I__1544\ : Span4Mux_h
    port map (
            O => \N__10833\,
            I => \N__10822\
        );

    \I__1543\ : Span4Mux_h
    port map (
            O => \N__10830\,
            I => \N__10819\
        );

    \I__1542\ : InMux
    port map (
            O => \N__10829\,
            I => \N__10816\
        );

    \I__1541\ : InMux
    port map (
            O => \N__10828\,
            I => \N__10813\
        );

    \I__1540\ : Odrv12
    port map (
            O => \N__10825\,
            I => \b2v_inst.reg_ancho_1Z0Z_6\
        );

    \I__1539\ : Odrv4
    port map (
            O => \N__10822\,
            I => \b2v_inst.reg_ancho_1Z0Z_6\
        );

    \I__1538\ : Odrv4
    port map (
            O => \N__10819\,
            I => \b2v_inst.reg_ancho_1Z0Z_6\
        );

    \I__1537\ : LocalMux
    port map (
            O => \N__10816\,
            I => \b2v_inst.reg_ancho_1Z0Z_6\
        );

    \I__1536\ : LocalMux
    port map (
            O => \N__10813\,
            I => \b2v_inst.reg_ancho_1Z0Z_6\
        );

    \I__1535\ : InMux
    port map (
            O => \N__10802\,
            I => \N__10798\
        );

    \I__1534\ : InMux
    port map (
            O => \N__10801\,
            I => \N__10795\
        );

    \I__1533\ : LocalMux
    port map (
            O => \N__10798\,
            I => \N__10790\
        );

    \I__1532\ : LocalMux
    port map (
            O => \N__10795\,
            I => \N__10787\
        );

    \I__1531\ : CascadeMux
    port map (
            O => \N__10794\,
            I => \N__10784\
        );

    \I__1530\ : InMux
    port map (
            O => \N__10793\,
            I => \N__10780\
        );

    \I__1529\ : Span4Mux_v
    port map (
            O => \N__10790\,
            I => \N__10777\
        );

    \I__1528\ : Span4Mux_h
    port map (
            O => \N__10787\,
            I => \N__10774\
        );

    \I__1527\ : InMux
    port map (
            O => \N__10784\,
            I => \N__10771\
        );

    \I__1526\ : InMux
    port map (
            O => \N__10783\,
            I => \N__10768\
        );

    \I__1525\ : LocalMux
    port map (
            O => \N__10780\,
            I => \b2v_inst.reg_ancho_1Z0Z_7\
        );

    \I__1524\ : Odrv4
    port map (
            O => \N__10777\,
            I => \b2v_inst.reg_ancho_1Z0Z_7\
        );

    \I__1523\ : Odrv4
    port map (
            O => \N__10774\,
            I => \b2v_inst.reg_ancho_1Z0Z_7\
        );

    \I__1522\ : LocalMux
    port map (
            O => \N__10771\,
            I => \b2v_inst.reg_ancho_1Z0Z_7\
        );

    \I__1521\ : LocalMux
    port map (
            O => \N__10768\,
            I => \b2v_inst.reg_ancho_1Z0Z_7\
        );

    \I__1520\ : CascadeMux
    port map (
            O => \N__10757\,
            I => \N__10753\
        );

    \I__1519\ : CascadeMux
    port map (
            O => \N__10756\,
            I => \N__10749\
        );

    \I__1518\ : InMux
    port map (
            O => \N__10753\,
            I => \N__10746\
        );

    \I__1517\ : InMux
    port map (
            O => \N__10752\,
            I => \N__10743\
        );

    \I__1516\ : InMux
    port map (
            O => \N__10749\,
            I => \N__10740\
        );

    \I__1515\ : LocalMux
    port map (
            O => \N__10746\,
            I => \N__10735\
        );

    \I__1514\ : LocalMux
    port map (
            O => \N__10743\,
            I => \N__10735\
        );

    \I__1513\ : LocalMux
    port map (
            O => \N__10740\,
            I => \b2v_inst.reg_ancho_3Z0Z_7\
        );

    \I__1512\ : Odrv4
    port map (
            O => \N__10735\,
            I => \b2v_inst.reg_ancho_3Z0Z_7\
        );

    \I__1511\ : InMux
    port map (
            O => \N__10730\,
            I => \bfn_5_18_0_\
        );

    \I__1510\ : InMux
    port map (
            O => \N__10727\,
            I => \N__10724\
        );

    \I__1509\ : LocalMux
    port map (
            O => \N__10724\,
            I => \N__10721\
        );

    \I__1508\ : Span4Mux_h
    port map (
            O => \N__10721\,
            I => \N__10718\
        );

    \I__1507\ : Odrv4
    port map (
            O => \N__10718\,
            I => \b2v_inst.valor_max_final50_THRU_CO\
        );

    \I__1506\ : InMux
    port map (
            O => \N__10715\,
            I => \N__10712\
        );

    \I__1505\ : LocalMux
    port map (
            O => \N__10712\,
            I => \N__10709\
        );

    \I__1504\ : Odrv4
    port map (
            O => \N__10709\,
            I => \b2v_inst.data_a_escribir9_5_and\
        );

    \I__1503\ : InMux
    port map (
            O => \N__10706\,
            I => \N__10702\
        );

    \I__1502\ : InMux
    port map (
            O => \N__10705\,
            I => \N__10697\
        );

    \I__1501\ : LocalMux
    port map (
            O => \N__10702\,
            I => \N__10692\
        );

    \I__1500\ : InMux
    port map (
            O => \N__10701\,
            I => \N__10689\
        );

    \I__1499\ : InMux
    port map (
            O => \N__10700\,
            I => \N__10685\
        );

    \I__1498\ : LocalMux
    port map (
            O => \N__10697\,
            I => \N__10682\
        );

    \I__1497\ : InMux
    port map (
            O => \N__10696\,
            I => \N__10673\
        );

    \I__1496\ : InMux
    port map (
            O => \N__10695\,
            I => \N__10673\
        );

    \I__1495\ : Span4Mux_v
    port map (
            O => \N__10692\,
            I => \N__10668\
        );

    \I__1494\ : LocalMux
    port map (
            O => \N__10689\,
            I => \N__10668\
        );

    \I__1493\ : InMux
    port map (
            O => \N__10688\,
            I => \N__10665\
        );

    \I__1492\ : LocalMux
    port map (
            O => \N__10685\,
            I => \N__10662\
        );

    \I__1491\ : Span4Mux_v
    port map (
            O => \N__10682\,
            I => \N__10659\
        );

    \I__1490\ : InMux
    port map (
            O => \N__10681\,
            I => \N__10654\
        );

    \I__1489\ : InMux
    port map (
            O => \N__10680\,
            I => \N__10654\
        );

    \I__1488\ : InMux
    port map (
            O => \N__10679\,
            I => \N__10649\
        );

    \I__1487\ : InMux
    port map (
            O => \N__10678\,
            I => \N__10649\
        );

    \I__1486\ : LocalMux
    port map (
            O => \N__10673\,
            I => \N__10646\
        );

    \I__1485\ : Span4Mux_h
    port map (
            O => \N__10668\,
            I => \N__10641\
        );

    \I__1484\ : LocalMux
    port map (
            O => \N__10665\,
            I => \N__10641\
        );

    \I__1483\ : Odrv4
    port map (
            O => \N__10662\,
            I => \b2v_inst.un3_valor_max1_THRU_CO\
        );

    \I__1482\ : Odrv4
    port map (
            O => \N__10659\,
            I => \b2v_inst.un3_valor_max1_THRU_CO\
        );

    \I__1481\ : LocalMux
    port map (
            O => \N__10654\,
            I => \b2v_inst.un3_valor_max1_THRU_CO\
        );

    \I__1480\ : LocalMux
    port map (
            O => \N__10649\,
            I => \b2v_inst.un3_valor_max1_THRU_CO\
        );

    \I__1479\ : Odrv4
    port map (
            O => \N__10646\,
            I => \b2v_inst.un3_valor_max1_THRU_CO\
        );

    \I__1478\ : Odrv4
    port map (
            O => \N__10641\,
            I => \b2v_inst.un3_valor_max1_THRU_CO\
        );

    \I__1477\ : InMux
    port map (
            O => \N__10628\,
            I => \N__10625\
        );

    \I__1476\ : LocalMux
    port map (
            O => \N__10625\,
            I => \N__10622\
        );

    \I__1475\ : Odrv4
    port map (
            O => \N__10622\,
            I => \b2v_inst.data_a_escribir_RNO_3Z0Z_6\
        );

    \I__1474\ : InMux
    port map (
            O => \N__10619\,
            I => \N__10616\
        );

    \I__1473\ : LocalMux
    port map (
            O => \N__10616\,
            I => \N__10613\
        );

    \I__1472\ : Span4Mux_h
    port map (
            O => \N__10613\,
            I => \N__10607\
        );

    \I__1471\ : InMux
    port map (
            O => \N__10612\,
            I => \N__10604\
        );

    \I__1470\ : InMux
    port map (
            O => \N__10611\,
            I => \N__10601\
        );

    \I__1469\ : InMux
    port map (
            O => \N__10610\,
            I => \N__10598\
        );

    \I__1468\ : Odrv4
    port map (
            O => \N__10607\,
            I => \b2v_inst.un1_reg_anterior_iv_0_0_a2_6_0_1\
        );

    \I__1467\ : LocalMux
    port map (
            O => \N__10604\,
            I => \b2v_inst.un1_reg_anterior_iv_0_0_a2_6_0_1\
        );

    \I__1466\ : LocalMux
    port map (
            O => \N__10601\,
            I => \b2v_inst.un1_reg_anterior_iv_0_0_a2_6_0_1\
        );

    \I__1465\ : LocalMux
    port map (
            O => \N__10598\,
            I => \b2v_inst.un1_reg_anterior_iv_0_0_a2_6_0_1\
        );

    \I__1464\ : InMux
    port map (
            O => \N__10589\,
            I => \N__10586\
        );

    \I__1463\ : LocalMux
    port map (
            O => \N__10586\,
            I => \b2v_inst.un1_m3_0_0\
        );

    \I__1462\ : InMux
    port map (
            O => \N__10583\,
            I => \N__10580\
        );

    \I__1461\ : LocalMux
    port map (
            O => \N__10580\,
            I => \N__10577\
        );

    \I__1460\ : Odrv4
    port map (
            O => \N__10577\,
            I => \b2v_inst.un1_reg_anterior_iv_0_0_0_6\
        );

    \I__1459\ : CascadeMux
    port map (
            O => \N__10574\,
            I => \b2v_inst.data_a_escribir_RNO_1Z0Z_6_cascade_\
        );

    \I__1458\ : CascadeMux
    port map (
            O => \N__10571\,
            I => \N__10564\
        );

    \I__1457\ : CascadeMux
    port map (
            O => \N__10570\,
            I => \N__10559\
        );

    \I__1456\ : CascadeMux
    port map (
            O => \N__10569\,
            I => \N__10554\
        );

    \I__1455\ : InMux
    port map (
            O => \N__10568\,
            I => \N__10548\
        );

    \I__1454\ : InMux
    port map (
            O => \N__10567\,
            I => \N__10548\
        );

    \I__1453\ : InMux
    port map (
            O => \N__10564\,
            I => \N__10537\
        );

    \I__1452\ : InMux
    port map (
            O => \N__10563\,
            I => \N__10534\
        );

    \I__1451\ : InMux
    port map (
            O => \N__10562\,
            I => \N__10531\
        );

    \I__1450\ : InMux
    port map (
            O => \N__10559\,
            I => \N__10528\
        );

    \I__1449\ : InMux
    port map (
            O => \N__10558\,
            I => \N__10519\
        );

    \I__1448\ : InMux
    port map (
            O => \N__10557\,
            I => \N__10519\
        );

    \I__1447\ : InMux
    port map (
            O => \N__10554\,
            I => \N__10519\
        );

    \I__1446\ : InMux
    port map (
            O => \N__10553\,
            I => \N__10519\
        );

    \I__1445\ : LocalMux
    port map (
            O => \N__10548\,
            I => \N__10507\
        );

    \I__1444\ : InMux
    port map (
            O => \N__10547\,
            I => \N__10494\
        );

    \I__1443\ : InMux
    port map (
            O => \N__10546\,
            I => \N__10494\
        );

    \I__1442\ : InMux
    port map (
            O => \N__10545\,
            I => \N__10494\
        );

    \I__1441\ : InMux
    port map (
            O => \N__10544\,
            I => \N__10494\
        );

    \I__1440\ : InMux
    port map (
            O => \N__10543\,
            I => \N__10494\
        );

    \I__1439\ : InMux
    port map (
            O => \N__10542\,
            I => \N__10494\
        );

    \I__1438\ : InMux
    port map (
            O => \N__10541\,
            I => \N__10489\
        );

    \I__1437\ : InMux
    port map (
            O => \N__10540\,
            I => \N__10489\
        );

    \I__1436\ : LocalMux
    port map (
            O => \N__10537\,
            I => \N__10482\
        );

    \I__1435\ : LocalMux
    port map (
            O => \N__10534\,
            I => \N__10482\
        );

    \I__1434\ : LocalMux
    port map (
            O => \N__10531\,
            I => \N__10482\
        );

    \I__1433\ : LocalMux
    port map (
            O => \N__10528\,
            I => \N__10477\
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__10519\,
            I => \N__10477\
        );

    \I__1431\ : InMux
    port map (
            O => \N__10518\,
            I => \N__10472\
        );

    \I__1430\ : InMux
    port map (
            O => \N__10517\,
            I => \N__10472\
        );

    \I__1429\ : InMux
    port map (
            O => \N__10516\,
            I => \N__10467\
        );

    \I__1428\ : InMux
    port map (
            O => \N__10515\,
            I => \N__10467\
        );

    \I__1427\ : InMux
    port map (
            O => \N__10514\,
            I => \N__10456\
        );

    \I__1426\ : InMux
    port map (
            O => \N__10513\,
            I => \N__10456\
        );

    \I__1425\ : InMux
    port map (
            O => \N__10512\,
            I => \N__10456\
        );

    \I__1424\ : InMux
    port map (
            O => \N__10511\,
            I => \N__10456\
        );

    \I__1423\ : InMux
    port map (
            O => \N__10510\,
            I => \N__10456\
        );

    \I__1422\ : Span4Mux_h
    port map (
            O => \N__10507\,
            I => \N__10451\
        );

    \I__1421\ : LocalMux
    port map (
            O => \N__10494\,
            I => \N__10451\
        );

    \I__1420\ : LocalMux
    port map (
            O => \N__10489\,
            I => \N__10444\
        );

    \I__1419\ : Span4Mux_v
    port map (
            O => \N__10482\,
            I => \N__10444\
        );

    \I__1418\ : Span4Mux_h
    port map (
            O => \N__10477\,
            I => \N__10444\
        );

    \I__1417\ : LocalMux
    port map (
            O => \N__10472\,
            I => \b2v_inst.data_a_escribir10_THRU_CO\
        );

    \I__1416\ : LocalMux
    port map (
            O => \N__10467\,
            I => \b2v_inst.data_a_escribir10_THRU_CO\
        );

    \I__1415\ : LocalMux
    port map (
            O => \N__10456\,
            I => \b2v_inst.data_a_escribir10_THRU_CO\
        );

    \I__1414\ : Odrv4
    port map (
            O => \N__10451\,
            I => \b2v_inst.data_a_escribir10_THRU_CO\
        );

    \I__1413\ : Odrv4
    port map (
            O => \N__10444\,
            I => \b2v_inst.data_a_escribir10_THRU_CO\
        );

    \I__1412\ : InMux
    port map (
            O => \N__10433\,
            I => \N__10420\
        );

    \I__1411\ : InMux
    port map (
            O => \N__10432\,
            I => \N__10420\
        );

    \I__1410\ : InMux
    port map (
            O => \N__10431\,
            I => \N__10414\
        );

    \I__1409\ : InMux
    port map (
            O => \N__10430\,
            I => \N__10414\
        );

    \I__1408\ : InMux
    port map (
            O => \N__10429\,
            I => \N__10411\
        );

    \I__1407\ : InMux
    port map (
            O => \N__10428\,
            I => \N__10406\
        );

    \I__1406\ : InMux
    port map (
            O => \N__10427\,
            I => \N__10406\
        );

    \I__1405\ : InMux
    port map (
            O => \N__10426\,
            I => \N__10401\
        );

    \I__1404\ : InMux
    port map (
            O => \N__10425\,
            I => \N__10401\
        );

    \I__1403\ : LocalMux
    port map (
            O => \N__10420\,
            I => \N__10398\
        );

    \I__1402\ : InMux
    port map (
            O => \N__10419\,
            I => \N__10395\
        );

    \I__1401\ : LocalMux
    port map (
            O => \N__10414\,
            I => \N__10392\
        );

    \I__1400\ : LocalMux
    port map (
            O => \N__10411\,
            I => \N__10383\
        );

    \I__1399\ : LocalMux
    port map (
            O => \N__10406\,
            I => \N__10383\
        );

    \I__1398\ : LocalMux
    port map (
            O => \N__10401\,
            I => \N__10383\
        );

    \I__1397\ : Span4Mux_h
    port map (
            O => \N__10398\,
            I => \N__10383\
        );

    \I__1396\ : LocalMux
    port map (
            O => \N__10395\,
            I => \b2v_inst.N_264\
        );

    \I__1395\ : Odrv4
    port map (
            O => \N__10392\,
            I => \b2v_inst.N_264\
        );

    \I__1394\ : Odrv4
    port map (
            O => \N__10383\,
            I => \b2v_inst.N_264\
        );

    \I__1393\ : InMux
    port map (
            O => \N__10376\,
            I => \N__10373\
        );

    \I__1392\ : LocalMux
    port map (
            O => \N__10373\,
            I => \N__10370\
        );

    \I__1391\ : Odrv4
    port map (
            O => \N__10370\,
            I => \b2v_inst.un1_reg_anterior_iv_0_0_0_7\
        );

    \I__1390\ : CascadeMux
    port map (
            O => \N__10367\,
            I => \b2v_inst.un1_reg_anterior_iv_0_0_3_0_7_cascade_\
        );

    \I__1389\ : InMux
    port map (
            O => \N__10364\,
            I => \N__10361\
        );

    \I__1388\ : LocalMux
    port map (
            O => \N__10361\,
            I => \N__10358\
        );

    \I__1387\ : Span4Mux_h
    port map (
            O => \N__10358\,
            I => \N__10355\
        );

    \I__1386\ : Odrv4
    port map (
            O => \N__10355\,
            I => \b2v_inst.un1_reg_anterior_iv_0_0_2_0_tz_7\
        );

    \I__1385\ : CEMux
    port map (
            O => \N__10352\,
            I => \N__10346\
        );

    \I__1384\ : CEMux
    port map (
            O => \N__10351\,
            I => \N__10343\
        );

    \I__1383\ : CEMux
    port map (
            O => \N__10350\,
            I => \N__10340\
        );

    \I__1382\ : CEMux
    port map (
            O => \N__10349\,
            I => \N__10337\
        );

    \I__1381\ : LocalMux
    port map (
            O => \N__10346\,
            I => \N__10334\
        );

    \I__1380\ : LocalMux
    port map (
            O => \N__10343\,
            I => \N__10330\
        );

    \I__1379\ : LocalMux
    port map (
            O => \N__10340\,
            I => \N__10327\
        );

    \I__1378\ : LocalMux
    port map (
            O => \N__10337\,
            I => \N__10324\
        );

    \I__1377\ : Span4Mux_v
    port map (
            O => \N__10334\,
            I => \N__10321\
        );

    \I__1376\ : CEMux
    port map (
            O => \N__10333\,
            I => \N__10318\
        );

    \I__1375\ : Span4Mux_h
    port map (
            O => \N__10330\,
            I => \N__10315\
        );

    \I__1374\ : Span4Mux_h
    port map (
            O => \N__10327\,
            I => \N__10312\
        );

    \I__1373\ : Span4Mux_h
    port map (
            O => \N__10324\,
            I => \N__10307\
        );

    \I__1372\ : Span4Mux_v
    port map (
            O => \N__10321\,
            I => \N__10307\
        );

    \I__1371\ : LocalMux
    port map (
            O => \N__10318\,
            I => \N__10302\
        );

    \I__1370\ : Span4Mux_h
    port map (
            O => \N__10315\,
            I => \N__10302\
        );

    \I__1369\ : Odrv4
    port map (
            O => \N__10312\,
            I => \b2v_inst.un1_reset_inv_2_0\
        );

    \I__1368\ : Odrv4
    port map (
            O => \N__10307\,
            I => \b2v_inst.un1_reset_inv_2_0\
        );

    \I__1367\ : Odrv4
    port map (
            O => \N__10302\,
            I => \b2v_inst.un1_reset_inv_2_0\
        );

    \I__1366\ : InMux
    port map (
            O => \N__10295\,
            I => \N__10291\
        );

    \I__1365\ : InMux
    port map (
            O => \N__10294\,
            I => \N__10288\
        );

    \I__1364\ : LocalMux
    port map (
            O => \N__10291\,
            I => \N__10283\
        );

    \I__1363\ : LocalMux
    port map (
            O => \N__10288\,
            I => \N__10279\
        );

    \I__1362\ : InMux
    port map (
            O => \N__10287\,
            I => \N__10276\
        );

    \I__1361\ : InMux
    port map (
            O => \N__10286\,
            I => \N__10273\
        );

    \I__1360\ : Span4Mux_v
    port map (
            O => \N__10283\,
            I => \N__10270\
        );

    \I__1359\ : InMux
    port map (
            O => \N__10282\,
            I => \N__10267\
        );

    \I__1358\ : Span4Mux_h
    port map (
            O => \N__10279\,
            I => \N__10264\
        );

    \I__1357\ : LocalMux
    port map (
            O => \N__10276\,
            I => \N__10259\
        );

    \I__1356\ : LocalMux
    port map (
            O => \N__10273\,
            I => \N__10259\
        );

    \I__1355\ : Odrv4
    port map (
            O => \N__10270\,
            I => \b2v_inst.reg_ancho_1Z0Z_0\
        );

    \I__1354\ : LocalMux
    port map (
            O => \N__10267\,
            I => \b2v_inst.reg_ancho_1Z0Z_0\
        );

    \I__1353\ : Odrv4
    port map (
            O => \N__10264\,
            I => \b2v_inst.reg_ancho_1Z0Z_0\
        );

    \I__1352\ : Odrv4
    port map (
            O => \N__10259\,
            I => \b2v_inst.reg_ancho_1Z0Z_0\
        );

    \I__1351\ : InMux
    port map (
            O => \N__10250\,
            I => \N__10247\
        );

    \I__1350\ : LocalMux
    port map (
            O => \N__10247\,
            I => \N__10243\
        );

    \I__1349\ : InMux
    port map (
            O => \N__10246\,
            I => \N__10239\
        );

    \I__1348\ : Span4Mux_v
    port map (
            O => \N__10243\,
            I => \N__10236\
        );

    \I__1347\ : InMux
    port map (
            O => \N__10242\,
            I => \N__10233\
        );

    \I__1346\ : LocalMux
    port map (
            O => \N__10239\,
            I => \N__10230\
        );

    \I__1345\ : Odrv4
    port map (
            O => \N__10236\,
            I => \b2v_inst.reg_ancho_3Z0Z_0\
        );

    \I__1344\ : LocalMux
    port map (
            O => \N__10233\,
            I => \b2v_inst.reg_ancho_3Z0Z_0\
        );

    \I__1343\ : Odrv4
    port map (
            O => \N__10230\,
            I => \b2v_inst.reg_ancho_3Z0Z_0\
        );

    \I__1342\ : CascadeMux
    port map (
            O => \N__10223\,
            I => \N_458_cascade_\
        );

    \I__1341\ : CascadeMux
    port map (
            O => \N__10220\,
            I => \b2v_inst.N_429_cascade_\
        );

    \I__1340\ : InMux
    port map (
            O => \N__10217\,
            I => \N__10214\
        );

    \I__1339\ : LocalMux
    port map (
            O => \N__10214\,
            I => \N__10211\
        );

    \I__1338\ : Span4Mux_h
    port map (
            O => \N__10211\,
            I => \N__10203\
        );

    \I__1337\ : InMux
    port map (
            O => \N__10210\,
            I => \N__10198\
        );

    \I__1336\ : InMux
    port map (
            O => \N__10209\,
            I => \N__10198\
        );

    \I__1335\ : InMux
    port map (
            O => \N__10208\,
            I => \N__10191\
        );

    \I__1334\ : InMux
    port map (
            O => \N__10207\,
            I => \N__10191\
        );

    \I__1333\ : InMux
    port map (
            O => \N__10206\,
            I => \N__10191\
        );

    \I__1332\ : Odrv4
    port map (
            O => \N__10203\,
            I => \b2v_inst.un1_pix_count_anterior_0_N_2_THRU_CO\
        );

    \I__1331\ : LocalMux
    port map (
            O => \N__10198\,
            I => \b2v_inst.un1_pix_count_anterior_0_N_2_THRU_CO\
        );

    \I__1330\ : LocalMux
    port map (
            O => \N__10191\,
            I => \b2v_inst.un1_pix_count_anterior_0_N_2_THRU_CO\
        );

    \I__1329\ : InMux
    port map (
            O => \N__10184\,
            I => \N__10175\
        );

    \I__1328\ : InMux
    port map (
            O => \N__10183\,
            I => \N__10175\
        );

    \I__1327\ : InMux
    port map (
            O => \N__10182\,
            I => \N__10175\
        );

    \I__1326\ : LocalMux
    port map (
            O => \N__10175\,
            I => \b2v_inst.stateZ0Z_3\
        );

    \I__1325\ : CascadeMux
    port map (
            O => \N__10172\,
            I => \N__10168\
        );

    \I__1324\ : IoInMux
    port map (
            O => \N__10171\,
            I => \N__10165\
        );

    \I__1323\ : InMux
    port map (
            O => \N__10168\,
            I => \N__10161\
        );

    \I__1322\ : LocalMux
    port map (
            O => \N__10165\,
            I => \N__10158\
        );

    \I__1321\ : InMux
    port map (
            O => \N__10164\,
            I => \N__10154\
        );

    \I__1320\ : LocalMux
    port map (
            O => \N__10161\,
            I => \N__10151\
        );

    \I__1319\ : IoSpan4Mux
    port map (
            O => \N__10158\,
            I => \N__10148\
        );

    \I__1318\ : CascadeMux
    port map (
            O => \N__10157\,
            I => \N__10145\
        );

    \I__1317\ : LocalMux
    port map (
            O => \N__10154\,
            I => \N__10140\
        );

    \I__1316\ : Span4Mux_v
    port map (
            O => \N__10151\,
            I => \N__10137\
        );

    \I__1315\ : Sp12to4
    port map (
            O => \N__10148\,
            I => \N__10134\
        );

    \I__1314\ : InMux
    port map (
            O => \N__10145\,
            I => \N__10131\
        );

    \I__1313\ : InMux
    port map (
            O => \N__10144\,
            I => \N__10126\
        );

    \I__1312\ : InMux
    port map (
            O => \N__10143\,
            I => \N__10126\
        );

    \I__1311\ : Span4Mux_v
    port map (
            O => \N__10140\,
            I => \N__10123\
        );

    \I__1310\ : Span4Mux_h
    port map (
            O => \N__10137\,
            I => \N__10120\
        );

    \I__1309\ : Span12Mux_v
    port map (
            O => \N__10134\,
            I => \N__10117\
        );

    \I__1308\ : LocalMux
    port map (
            O => \N__10131\,
            I => \b2v_inst.stateZ0Z_2\
        );

    \I__1307\ : LocalMux
    port map (
            O => \N__10126\,
            I => \b2v_inst.stateZ0Z_2\
        );

    \I__1306\ : Odrv4
    port map (
            O => \N__10123\,
            I => \b2v_inst.stateZ0Z_2\
        );

    \I__1305\ : Odrv4
    port map (
            O => \N__10120\,
            I => \b2v_inst.stateZ0Z_2\
        );

    \I__1304\ : Odrv12
    port map (
            O => \N__10117\,
            I => \b2v_inst.stateZ0Z_2\
        );

    \I__1303\ : CascadeMux
    port map (
            O => \N__10106\,
            I => \N__10103\
        );

    \I__1302\ : InMux
    port map (
            O => \N__10103\,
            I => \N__10100\
        );

    \I__1301\ : LocalMux
    port map (
            O => \N__10100\,
            I => \N__10097\
        );

    \I__1300\ : Odrv4
    port map (
            O => \N__10097\,
            I => \b2v_inst.data_a_escribir9_4_and\
        );

    \I__1299\ : InMux
    port map (
            O => \N__10094\,
            I => \N__10091\
        );

    \I__1298\ : LocalMux
    port map (
            O => \N__10091\,
            I => \N__10088\
        );

    \I__1297\ : Span4Mux_v
    port map (
            O => \N__10088\,
            I => \N__10085\
        );

    \I__1296\ : Odrv4
    port map (
            O => \N__10085\,
            I => \SYNTHESIZED_WIRE_3_3\
        );

    \I__1295\ : InMux
    port map (
            O => \N__10082\,
            I => \N__10079\
        );

    \I__1294\ : LocalMux
    port map (
            O => \N__10079\,
            I => \N__10076\
        );

    \I__1293\ : Span4Mux_h
    port map (
            O => \N__10076\,
            I => \N__10073\
        );

    \I__1292\ : Odrv4
    port map (
            O => \N__10073\,
            I => \SYNTHESIZED_WIRE_3_4\
        );

    \I__1291\ : InMux
    port map (
            O => \N__10070\,
            I => \N__10067\
        );

    \I__1290\ : LocalMux
    port map (
            O => \N__10067\,
            I => \N__10064\
        );

    \I__1289\ : Span4Mux_h
    port map (
            O => \N__10064\,
            I => \N__10061\
        );

    \I__1288\ : Odrv4
    port map (
            O => \N__10061\,
            I => \SYNTHESIZED_WIRE_3_5\
        );

    \I__1287\ : CascadeMux
    port map (
            O => \N__10058\,
            I => \N__10055\
        );

    \I__1286\ : InMux
    port map (
            O => \N__10055\,
            I => \N__10052\
        );

    \I__1285\ : LocalMux
    port map (
            O => \N__10052\,
            I => \N__10049\
        );

    \I__1284\ : Span4Mux_h
    port map (
            O => \N__10049\,
            I => \N__10046\
        );

    \I__1283\ : Odrv4
    port map (
            O => \N__10046\,
            I => \SYNTHESIZED_WIRE_3_6\
        );

    \I__1282\ : CascadeMux
    port map (
            O => \N__10043\,
            I => \N__10040\
        );

    \I__1281\ : InMux
    port map (
            O => \N__10040\,
            I => \N__10037\
        );

    \I__1280\ : LocalMux
    port map (
            O => \N__10037\,
            I => \N__10034\
        );

    \I__1279\ : Span4Mux_v
    port map (
            O => \N__10034\,
            I => \N__10031\
        );

    \I__1278\ : Odrv4
    port map (
            O => \N__10031\,
            I => \SYNTHESIZED_WIRE_3_7\
        );

    \I__1277\ : CEMux
    port map (
            O => \N__10028\,
            I => \N__10024\
        );

    \I__1276\ : CascadeMux
    port map (
            O => \N__10027\,
            I => \N__10020\
        );

    \I__1275\ : LocalMux
    port map (
            O => \N__10024\,
            I => \N__10017\
        );

    \I__1274\ : InMux
    port map (
            O => \N__10023\,
            I => \N__10014\
        );

    \I__1273\ : InMux
    port map (
            O => \N__10020\,
            I => \N__10011\
        );

    \I__1272\ : Span4Mux_h
    port map (
            O => \N__10017\,
            I => \N__10008\
        );

    \I__1271\ : LocalMux
    port map (
            O => \N__10014\,
            I => \N__10005\
        );

    \I__1270\ : LocalMux
    port map (
            O => \N__10011\,
            I => \N__10002\
        );

    \I__1269\ : Odrv4
    port map (
            O => \N__10008\,
            I => \b2v_inst4.pix_count_int_0_sqmuxa\
        );

    \I__1268\ : Odrv4
    port map (
            O => \N__10005\,
            I => \b2v_inst4.pix_count_int_0_sqmuxa\
        );

    \I__1267\ : Odrv4
    port map (
            O => \N__10002\,
            I => \b2v_inst4.pix_count_int_0_sqmuxa\
        );

    \I__1266\ : CascadeMux
    port map (
            O => \N__9995\,
            I => \b2v_inst.we_0_a2_0_a2_4_cascade_\
        );

    \I__1265\ : CEMux
    port map (
            O => \N__9992\,
            I => \N__9989\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__9989\,
            I => \N__9986\
        );

    \I__1263\ : Span4Mux_v
    port map (
            O => \N__9986\,
            I => \N__9983\
        );

    \I__1262\ : Odrv4
    port map (
            O => \N__9983\,
            I => \SYNTHESIZED_WIRE_4\
        );

    \I__1261\ : InMux
    port map (
            O => \N__9980\,
            I => \N__9977\
        );

    \I__1260\ : LocalMux
    port map (
            O => \N__9977\,
            I => \b2v_inst.we_0_a2_0_a2_3\
        );

    \I__1259\ : CascadeMux
    port map (
            O => \N__9974\,
            I => \b2v_inst3.un1_m2_0_a2_2_cascade_\
        );

    \I__1258\ : CascadeMux
    port map (
            O => \N__9971\,
            I => \N__9967\
        );

    \I__1257\ : CascadeMux
    port map (
            O => \N__9970\,
            I => \N__9964\
        );

    \I__1256\ : InMux
    port map (
            O => \N__9967\,
            I => \N__9959\
        );

    \I__1255\ : InMux
    port map (
            O => \N__9964\,
            I => \N__9959\
        );

    \I__1254\ : LocalMux
    port map (
            O => \N__9959\,
            I => \b2v_inst3.un1_cycle_counter_5_c5\
        );

    \I__1253\ : CascadeMux
    port map (
            O => \N__9956\,
            I => \b2v_inst3.un1_cycle_counter_5_c5_cascade_\
        );

    \I__1252\ : InMux
    port map (
            O => \N__9953\,
            I => \N__9950\
        );

    \I__1251\ : LocalMux
    port map (
            O => \N__9950\,
            I => \N__9947\
        );

    \I__1250\ : Span4Mux_v
    port map (
            O => \N__9947\,
            I => \N__9943\
        );

    \I__1249\ : InMux
    port map (
            O => \N__9946\,
            I => \N__9940\
        );

    \I__1248\ : Odrv4
    port map (
            O => \N__9943\,
            I => \SYNTHESIZED_WIRE_10_0\
        );

    \I__1247\ : LocalMux
    port map (
            O => \N__9940\,
            I => \SYNTHESIZED_WIRE_10_0\
        );

    \I__1246\ : InMux
    port map (
            O => \N__9935\,
            I => \N__9932\
        );

    \I__1245\ : LocalMux
    port map (
            O => \N__9932\,
            I => \N__9929\
        );

    \I__1244\ : Span4Mux_h
    port map (
            O => \N__9929\,
            I => \N__9926\
        );

    \I__1243\ : Odrv4
    port map (
            O => \N__9926\,
            I => \SYNTHESIZED_WIRE_3_0\
        );

    \I__1242\ : InMux
    port map (
            O => \N__9923\,
            I => \N__9920\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__9920\,
            I => \N__9917\
        );

    \I__1240\ : Span4Mux_h
    port map (
            O => \N__9917\,
            I => \N__9914\
        );

    \I__1239\ : Odrv4
    port map (
            O => \N__9914\,
            I => \SYNTHESIZED_WIRE_3_1\
        );

    \I__1238\ : InMux
    port map (
            O => \N__9911\,
            I => \N__9908\
        );

    \I__1237\ : LocalMux
    port map (
            O => \N__9908\,
            I => \N__9905\
        );

    \I__1236\ : Span4Mux_v
    port map (
            O => \N__9905\,
            I => \N__9902\
        );

    \I__1235\ : Odrv4
    port map (
            O => \N__9902\,
            I => \SYNTHESIZED_WIRE_3_2\
        );

    \I__1234\ : InMux
    port map (
            O => \N__9899\,
            I => \N__9896\
        );

    \I__1233\ : LocalMux
    port map (
            O => \N__9896\,
            I => \b2v_inst.un1_reg_anterior_iv_0_0_2_tz_4\
        );

    \I__1232\ : CascadeMux
    port map (
            O => \N__9893\,
            I => \b2v_inst3.fsm_state_ns_0_0_0_1_cascade_\
        );

    \I__1231\ : CascadeMux
    port map (
            O => \N__9890\,
            I => \N_230_cascade_\
        );

    \I__1230\ : InMux
    port map (
            O => \N__9887\,
            I => \N__9884\
        );

    \I__1229\ : LocalMux
    port map (
            O => \N__9884\,
            I => \b2v_inst3.N_434\
        );

    \I__1228\ : InMux
    port map (
            O => \N__9881\,
            I => \N__9878\
        );

    \I__1227\ : LocalMux
    port map (
            O => \N__9878\,
            I => \b2v_inst3.N_490\
        );

    \I__1226\ : CascadeMux
    port map (
            O => \N__9875\,
            I => \b2v_inst3.fsm_state_ns_i_i_1_0_cascade_\
        );

    \I__1225\ : CascadeMux
    port map (
            O => \N__9872\,
            I => \N__9868\
        );

    \I__1224\ : InMux
    port map (
            O => \N__9871\,
            I => \N__9865\
        );

    \I__1223\ : InMux
    port map (
            O => \N__9868\,
            I => \N__9862\
        );

    \I__1222\ : LocalMux
    port map (
            O => \N__9865\,
            I => \N__9859\
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__9862\,
            I => \b2v_inst.reg_anterior_i_1\
        );

    \I__1220\ : Odrv4
    port map (
            O => \N__9859\,
            I => \b2v_inst.reg_anterior_i_1\
        );

    \I__1219\ : CascadeMux
    port map (
            O => \N__9854\,
            I => \N__9850\
        );

    \I__1218\ : InMux
    port map (
            O => \N__9853\,
            I => \N__9847\
        );

    \I__1217\ : InMux
    port map (
            O => \N__9850\,
            I => \N__9844\
        );

    \I__1216\ : LocalMux
    port map (
            O => \N__9847\,
            I => \N__9841\
        );

    \I__1215\ : LocalMux
    port map (
            O => \N__9844\,
            I => \b2v_inst.reg_anterior_i_2\
        );

    \I__1214\ : Odrv4
    port map (
            O => \N__9841\,
            I => \b2v_inst.reg_anterior_i_2\
        );

    \I__1213\ : CascadeMux
    port map (
            O => \N__9836\,
            I => \N__9832\
        );

    \I__1212\ : InMux
    port map (
            O => \N__9835\,
            I => \N__9829\
        );

    \I__1211\ : InMux
    port map (
            O => \N__9832\,
            I => \N__9826\
        );

    \I__1210\ : LocalMux
    port map (
            O => \N__9829\,
            I => \N__9823\
        );

    \I__1209\ : LocalMux
    port map (
            O => \N__9826\,
            I => \b2v_inst.reg_anterior_i_3\
        );

    \I__1208\ : Odrv4
    port map (
            O => \N__9823\,
            I => \b2v_inst.reg_anterior_i_3\
        );

    \I__1207\ : CascadeMux
    port map (
            O => \N__9818\,
            I => \N__9814\
        );

    \I__1206\ : CascadeMux
    port map (
            O => \N__9817\,
            I => \N__9811\
        );

    \I__1205\ : InMux
    port map (
            O => \N__9814\,
            I => \N__9808\
        );

    \I__1204\ : InMux
    port map (
            O => \N__9811\,
            I => \N__9805\
        );

    \I__1203\ : LocalMux
    port map (
            O => \N__9808\,
            I => \N__9802\
        );

    \I__1202\ : LocalMux
    port map (
            O => \N__9805\,
            I => \b2v_inst.reg_anterior_i_4\
        );

    \I__1201\ : Odrv4
    port map (
            O => \N__9802\,
            I => \b2v_inst.reg_anterior_i_4\
        );

    \I__1200\ : CascadeMux
    port map (
            O => \N__9797\,
            I => \N__9793\
        );

    \I__1199\ : CascadeMux
    port map (
            O => \N__9796\,
            I => \N__9790\
        );

    \I__1198\ : InMux
    port map (
            O => \N__9793\,
            I => \N__9787\
        );

    \I__1197\ : InMux
    port map (
            O => \N__9790\,
            I => \N__9784\
        );

    \I__1196\ : LocalMux
    port map (
            O => \N__9787\,
            I => \N__9781\
        );

    \I__1195\ : LocalMux
    port map (
            O => \N__9784\,
            I => \b2v_inst.reg_anterior_i_5\
        );

    \I__1194\ : Odrv4
    port map (
            O => \N__9781\,
            I => \b2v_inst.reg_anterior_i_5\
        );

    \I__1193\ : CascadeMux
    port map (
            O => \N__9776\,
            I => \N__9772\
        );

    \I__1192\ : CascadeMux
    port map (
            O => \N__9775\,
            I => \N__9769\
        );

    \I__1191\ : InMux
    port map (
            O => \N__9772\,
            I => \N__9766\
        );

    \I__1190\ : InMux
    port map (
            O => \N__9769\,
            I => \N__9763\
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__9766\,
            I => \N__9760\
        );

    \I__1188\ : LocalMux
    port map (
            O => \N__9763\,
            I => \N__9757\
        );

    \I__1187\ : Odrv4
    port map (
            O => \N__9760\,
            I => \b2v_inst.reg_anterior_i_6\
        );

    \I__1186\ : Odrv4
    port map (
            O => \N__9757\,
            I => \b2v_inst.reg_anterior_i_6\
        );

    \I__1185\ : InMux
    port map (
            O => \N__9752\,
            I => \N__9748\
        );

    \I__1184\ : CascadeMux
    port map (
            O => \N__9751\,
            I => \N__9745\
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__9748\,
            I => \N__9742\
        );

    \I__1182\ : InMux
    port map (
            O => \N__9745\,
            I => \N__9739\
        );

    \I__1181\ : Span4Mux_h
    port map (
            O => \N__9742\,
            I => \N__9736\
        );

    \I__1180\ : LocalMux
    port map (
            O => \N__9739\,
            I => \b2v_inst.reg_anterior_i_7\
        );

    \I__1179\ : Odrv4
    port map (
            O => \N__9736\,
            I => \b2v_inst.reg_anterior_i_7\
        );

    \I__1178\ : InMux
    port map (
            O => \N__9731\,
            I => \N__9728\
        );

    \I__1177\ : LocalMux
    port map (
            O => \N__9728\,
            I => \N__9724\
        );

    \I__1176\ : InMux
    port map (
            O => \N__9727\,
            I => \N__9721\
        );

    \I__1175\ : Odrv4
    port map (
            O => \N__9724\,
            I => \b2v_inst.valor_max_final53_THRU_CO\
        );

    \I__1174\ : LocalMux
    port map (
            O => \N__9721\,
            I => \b2v_inst.valor_max_final53_THRU_CO\
        );

    \I__1173\ : CascadeMux
    port map (
            O => \N__9716\,
            I => \N__9713\
        );

    \I__1172\ : InMux
    port map (
            O => \N__9713\,
            I => \N__9710\
        );

    \I__1171\ : LocalMux
    port map (
            O => \N__9710\,
            I => \b2v_inst.un1_m3_0_m3_ns_1\
        );

    \I__1170\ : InMux
    port map (
            O => \N__9707\,
            I => \bfn_3_20_0_\
        );

    \I__1169\ : InMux
    port map (
            O => \N__9704\,
            I => \N__9701\
        );

    \I__1168\ : LocalMux
    port map (
            O => \N__9701\,
            I => \N__9698\
        );

    \I__1167\ : Odrv12
    port map (
            O => \N__9698\,
            I => \b2v_inst.N_497\
        );

    \I__1166\ : InMux
    port map (
            O => \N__9695\,
            I => \N__9692\
        );

    \I__1165\ : LocalMux
    port map (
            O => \N__9692\,
            I => \N__9689\
        );

    \I__1164\ : Odrv4
    port map (
            O => \N__9689\,
            I => \b2v_inst.un1_reg_anterior_iv_0_0_2_tz_2\
        );

    \I__1163\ : CascadeMux
    port map (
            O => \N__9686\,
            I => \b2v_inst.data_a_escribir_RNO_1Z0Z_2_cascade_\
        );

    \I__1162\ : InMux
    port map (
            O => \N__9683\,
            I => \N__9680\
        );

    \I__1161\ : LocalMux
    port map (
            O => \N__9680\,
            I => \b2v_inst.un1_reg_anterior_iv_0_0_1_2\
        );

    \I__1160\ : CascadeMux
    port map (
            O => \N__9677\,
            I => \b2v_inst.data_a_escribir_RNO_4Z0Z_5_cascade_\
        );

    \I__1159\ : CascadeMux
    port map (
            O => \N__9674\,
            I => \b2v_inst.un1_reg_anterior_iv_0_0_2_1_5_cascade_\
        );

    \I__1158\ : InMux
    port map (
            O => \N__9671\,
            I => \N__9663\
        );

    \I__1157\ : InMux
    port map (
            O => \N__9670\,
            I => \N__9663\
        );

    \I__1156\ : InMux
    port map (
            O => \N__9669\,
            I => \N__9660\
        );

    \I__1155\ : InMux
    port map (
            O => \N__9668\,
            I => \N__9657\
        );

    \I__1154\ : LocalMux
    port map (
            O => \N__9663\,
            I => \b2v_inst.un1_reg_anterior_iv_0_0_a2_4_0_1\
        );

    \I__1153\ : LocalMux
    port map (
            O => \N__9660\,
            I => \b2v_inst.un1_reg_anterior_iv_0_0_a2_4_0_1\
        );

    \I__1152\ : LocalMux
    port map (
            O => \N__9657\,
            I => \b2v_inst.un1_reg_anterior_iv_0_0_a2_4_0_1\
        );

    \I__1151\ : InMux
    port map (
            O => \N__9650\,
            I => \N__9647\
        );

    \I__1150\ : LocalMux
    port map (
            O => \N__9647\,
            I => \N__9644\
        );

    \I__1149\ : Span4Mux_h
    port map (
            O => \N__9644\,
            I => \N__9641\
        );

    \I__1148\ : Odrv4
    port map (
            O => \N__9641\,
            I => \b2v_inst.un1_reg_anterior_iv_0_0_0_5\
        );

    \I__1147\ : CascadeMux
    port map (
            O => \N__9638\,
            I => \b2v_inst.data_a_escribir_RNO_0Z0Z_5_cascade_\
        );

    \I__1146\ : InMux
    port map (
            O => \N__9635\,
            I => \N__9632\
        );

    \I__1145\ : LocalMux
    port map (
            O => \N__9632\,
            I => \b2v_inst.data_a_escribir_RNO_1Z0Z_5\
        );

    \I__1144\ : CascadeMux
    port map (
            O => \N__9629\,
            I => \N__9625\
        );

    \I__1143\ : InMux
    port map (
            O => \N__9628\,
            I => \N__9622\
        );

    \I__1142\ : InMux
    port map (
            O => \N__9625\,
            I => \N__9619\
        );

    \I__1141\ : LocalMux
    port map (
            O => \N__9622\,
            I => \N__9616\
        );

    \I__1140\ : LocalMux
    port map (
            O => \N__9619\,
            I => \b2v_inst.reg_anterior_i_0\
        );

    \I__1139\ : Odrv4
    port map (
            O => \N__9616\,
            I => \b2v_inst.reg_anterior_i_0\
        );

    \I__1138\ : InMux
    port map (
            O => \N__9611\,
            I => \N__9608\
        );

    \I__1137\ : LocalMux
    port map (
            O => \N__9608\,
            I => \N__9605\
        );

    \I__1136\ : Span4Mux_h
    port map (
            O => \N__9605\,
            I => \N__9601\
        );

    \I__1135\ : InMux
    port map (
            O => \N__9604\,
            I => \N__9598\
        );

    \I__1134\ : Odrv4
    port map (
            O => \N__9601\,
            I => \b2v_inst.eventosZ0Z_1\
        );

    \I__1133\ : LocalMux
    port map (
            O => \N__9598\,
            I => \b2v_inst.eventosZ0Z_1\
        );

    \I__1132\ : InMux
    port map (
            O => \N__9593\,
            I => \N__9590\
        );

    \I__1131\ : LocalMux
    port map (
            O => \N__9590\,
            I => \N__9586\
        );

    \I__1130\ : InMux
    port map (
            O => \N__9589\,
            I => \N__9583\
        );

    \I__1129\ : Span12Mux_s11_v
    port map (
            O => \N__9586\,
            I => \N__9580\
        );

    \I__1128\ : LocalMux
    port map (
            O => \N__9583\,
            I => \b2v_inst.eventosZ0Z_6\
        );

    \I__1127\ : Odrv12
    port map (
            O => \N__9580\,
            I => \b2v_inst.eventosZ0Z_6\
        );

    \I__1126\ : CascadeMux
    port map (
            O => \N__9575\,
            I => \b2v_inst.un1_reg_anterior_iv_0_0_2_1_1_cascade_\
        );

    \I__1125\ : CascadeMux
    port map (
            O => \N__9572\,
            I => \b2v_inst.data_a_escribir_RNO_4Z0Z_1_cascade_\
        );

    \I__1124\ : InMux
    port map (
            O => \N__9569\,
            I => \N__9566\
        );

    \I__1123\ : LocalMux
    port map (
            O => \N__9566\,
            I => \b2v_inst.un1_reg_anterior_iv_0_0_0_1\
        );

    \I__1122\ : InMux
    port map (
            O => \N__9563\,
            I => \N__9560\
        );

    \I__1121\ : LocalMux
    port map (
            O => \N__9560\,
            I => \b2v_inst.data_a_escribir_RNO_0Z0Z_1\
        );

    \I__1120\ : CascadeMux
    port map (
            O => \N__9557\,
            I => \b2v_inst.data_a_escribir_RNO_1Z0Z_1_cascade_\
        );

    \I__1119\ : InMux
    port map (
            O => \N__9554\,
            I => \N__9551\
        );

    \I__1118\ : LocalMux
    port map (
            O => \N__9551\,
            I => \N__9548\
        );

    \I__1117\ : Span4Mux_h
    port map (
            O => \N__9548\,
            I => \N__9545\
        );

    \I__1116\ : Odrv4
    port map (
            O => \N__9545\,
            I => \b2v_inst.data_a_escribir9_2_and\
        );

    \I__1115\ : InMux
    port map (
            O => \N__9542\,
            I => \N__9539\
        );

    \I__1114\ : LocalMux
    port map (
            O => \N__9539\,
            I => \N__9536\
        );

    \I__1113\ : Odrv4
    port map (
            O => \N__9536\,
            I => \b2v_inst.data_a_escribir9_3_and\
        );

    \I__1112\ : InMux
    port map (
            O => \N__9533\,
            I => \bfn_3_16_0_\
        );

    \I__1111\ : InMux
    port map (
            O => \N__9530\,
            I => \N__9527\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__9527\,
            I => \N__9523\
        );

    \I__1109\ : InMux
    port map (
            O => \N__9526\,
            I => \N__9520\
        );

    \I__1108\ : Span4Mux_h
    port map (
            O => \N__9523\,
            I => \N__9517\
        );

    \I__1107\ : LocalMux
    port map (
            O => \N__9520\,
            I => \b2v_inst.eventosZ0Z_7\
        );

    \I__1106\ : Odrv4
    port map (
            O => \N__9517\,
            I => \b2v_inst.eventosZ0Z_7\
        );

    \I__1105\ : InMux
    port map (
            O => \N__9512\,
            I => \N__9506\
        );

    \I__1104\ : InMux
    port map (
            O => \N__9511\,
            I => \N__9499\
        );

    \I__1103\ : InMux
    port map (
            O => \N__9510\,
            I => \N__9499\
        );

    \I__1102\ : InMux
    port map (
            O => \N__9509\,
            I => \N__9499\
        );

    \I__1101\ : LocalMux
    port map (
            O => \N__9506\,
            I => \SYNTHESIZED_WIRE_2_7\
        );

    \I__1100\ : LocalMux
    port map (
            O => \N__9499\,
            I => \SYNTHESIZED_WIRE_2_7\
        );

    \I__1099\ : InMux
    port map (
            O => \N__9494\,
            I => \N__9491\
        );

    \I__1098\ : LocalMux
    port map (
            O => \N__9491\,
            I => \b2v_inst4.pix_count_int_RNO_0Z0Z_7\
        );

    \I__1097\ : InMux
    port map (
            O => \N__9488\,
            I => \b2v_inst4.un1_pix_count_int_cry_6\
        );

    \I__1096\ : InMux
    port map (
            O => \N__9485\,
            I => \N__9479\
        );

    \I__1095\ : InMux
    port map (
            O => \N__9484\,
            I => \N__9472\
        );

    \I__1094\ : InMux
    port map (
            O => \N__9483\,
            I => \N__9472\
        );

    \I__1093\ : InMux
    port map (
            O => \N__9482\,
            I => \N__9472\
        );

    \I__1092\ : LocalMux
    port map (
            O => \N__9479\,
            I => \SYNTHESIZED_WIRE_2_8\
        );

    \I__1091\ : LocalMux
    port map (
            O => \N__9472\,
            I => \SYNTHESIZED_WIRE_2_8\
        );

    \I__1090\ : InMux
    port map (
            O => \N__9467\,
            I => \N__9464\
        );

    \I__1089\ : LocalMux
    port map (
            O => \N__9464\,
            I => \b2v_inst4.pix_count_int_RNO_0Z0Z_8\
        );

    \I__1088\ : InMux
    port map (
            O => \N__9461\,
            I => \bfn_3_14_0_\
        );

    \I__1087\ : InMux
    port map (
            O => \N__9458\,
            I => \b2v_inst4.un1_pix_count_int_cry_8\
        );

    \I__1086\ : InMux
    port map (
            O => \N__9455\,
            I => \N__9447\
        );

    \I__1085\ : InMux
    port map (
            O => \N__9454\,
            I => \N__9447\
        );

    \I__1084\ : InMux
    port map (
            O => \N__9453\,
            I => \N__9444\
        );

    \I__1083\ : InMux
    port map (
            O => \N__9452\,
            I => \N__9441\
        );

    \I__1082\ : LocalMux
    port map (
            O => \N__9447\,
            I => \N__9436\
        );

    \I__1081\ : LocalMux
    port map (
            O => \N__9444\,
            I => \N__9436\
        );

    \I__1080\ : LocalMux
    port map (
            O => \N__9441\,
            I => \SYNTHESIZED_WIRE_2_10\
        );

    \I__1079\ : Odrv4
    port map (
            O => \N__9436\,
            I => \SYNTHESIZED_WIRE_2_10\
        );

    \I__1078\ : InMux
    port map (
            O => \N__9431\,
            I => \b2v_inst4.un1_pix_count_int_cry_9\
        );

    \I__1077\ : InMux
    port map (
            O => \N__9428\,
            I => \N__9422\
        );

    \I__1076\ : InMux
    port map (
            O => \N__9427\,
            I => \N__9419\
        );

    \I__1075\ : InMux
    port map (
            O => \N__9426\,
            I => \N__9414\
        );

    \I__1074\ : InMux
    port map (
            O => \N__9425\,
            I => \N__9414\
        );

    \I__1073\ : LocalMux
    port map (
            O => \N__9422\,
            I => \SYNTHESIZED_WIRE_2_11\
        );

    \I__1072\ : LocalMux
    port map (
            O => \N__9419\,
            I => \SYNTHESIZED_WIRE_2_11\
        );

    \I__1071\ : LocalMux
    port map (
            O => \N__9414\,
            I => \SYNTHESIZED_WIRE_2_11\
        );

    \I__1070\ : InMux
    port map (
            O => \N__9407\,
            I => \N__9404\
        );

    \I__1069\ : LocalMux
    port map (
            O => \N__9404\,
            I => \b2v_inst4.pix_count_int_RNO_0Z0Z_11\
        );

    \I__1068\ : InMux
    port map (
            O => \N__9401\,
            I => \b2v_inst4.un1_pix_count_int_cry_10\
        );

    \I__1067\ : CascadeMux
    port map (
            O => \N__9398\,
            I => \N__9393\
        );

    \I__1066\ : InMux
    port map (
            O => \N__9397\,
            I => \N__9389\
        );

    \I__1065\ : InMux
    port map (
            O => \N__9396\,
            I => \N__9386\
        );

    \I__1064\ : InMux
    port map (
            O => \N__9393\,
            I => \N__9383\
        );

    \I__1063\ : InMux
    port map (
            O => \N__9392\,
            I => \N__9380\
        );

    \I__1062\ : LocalMux
    port map (
            O => \N__9389\,
            I => \SYNTHESIZED_WIRE_2_12\
        );

    \I__1061\ : LocalMux
    port map (
            O => \N__9386\,
            I => \SYNTHESIZED_WIRE_2_12\
        );

    \I__1060\ : LocalMux
    port map (
            O => \N__9383\,
            I => \SYNTHESIZED_WIRE_2_12\
        );

    \I__1059\ : LocalMux
    port map (
            O => \N__9380\,
            I => \SYNTHESIZED_WIRE_2_12\
        );

    \I__1058\ : InMux
    port map (
            O => \N__9371\,
            I => \b2v_inst4.un1_pix_count_int_cry_11\
        );

    \I__1057\ : InMux
    port map (
            O => \N__9368\,
            I => \N__9365\
        );

    \I__1056\ : LocalMux
    port map (
            O => \N__9365\,
            I => \b2v_inst4.pix_count_int_RNO_0Z0Z_12\
        );

    \I__1055\ : InMux
    port map (
            O => \N__9362\,
            I => \N__9359\
        );

    \I__1054\ : LocalMux
    port map (
            O => \N__9359\,
            I => \b2v_inst.data_a_escribir9_0_and\
        );

    \I__1053\ : InMux
    port map (
            O => \N__9356\,
            I => \N__9353\
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__9353\,
            I => \b2v_inst.data_a_escribir9_1_and\
        );

    \I__1051\ : CascadeMux
    port map (
            O => \N__9350\,
            I => \N__9347\
        );

    \I__1050\ : InMux
    port map (
            O => \N__9347\,
            I => \N__9344\
        );

    \I__1049\ : LocalMux
    port map (
            O => \N__9344\,
            I => \b2v_inst.pix_count_anteriorZ0Z_11\
        );

    \I__1048\ : CEMux
    port map (
            O => \N__9341\,
            I => \N__9323\
        );

    \I__1047\ : CEMux
    port map (
            O => \N__9340\,
            I => \N__9323\
        );

    \I__1046\ : CEMux
    port map (
            O => \N__9339\,
            I => \N__9323\
        );

    \I__1045\ : CEMux
    port map (
            O => \N__9338\,
            I => \N__9323\
        );

    \I__1044\ : CEMux
    port map (
            O => \N__9337\,
            I => \N__9323\
        );

    \I__1043\ : CEMux
    port map (
            O => \N__9336\,
            I => \N__9323\
        );

    \I__1042\ : GlobalMux
    port map (
            O => \N__9323\,
            I => \N__9320\
        );

    \I__1041\ : gio2CtrlBuf
    port map (
            O => \N__9320\,
            I => \b2v_inst.N_254_i_g\
        );

    \I__1040\ : CascadeMux
    port map (
            O => \N__9317\,
            I => \N__9314\
        );

    \I__1039\ : InMux
    port map (
            O => \N__9314\,
            I => \N__9311\
        );

    \I__1038\ : LocalMux
    port map (
            O => \N__9311\,
            I => \N__9305\
        );

    \I__1037\ : InMux
    port map (
            O => \N__9310\,
            I => \N__9302\
        );

    \I__1036\ : InMux
    port map (
            O => \N__9309\,
            I => \N__9297\
        );

    \I__1035\ : InMux
    port map (
            O => \N__9308\,
            I => \N__9297\
        );

    \I__1034\ : Odrv4
    port map (
            O => \N__9305\,
            I => \SYNTHESIZED_WIRE_2_0\
        );

    \I__1033\ : LocalMux
    port map (
            O => \N__9302\,
            I => \SYNTHESIZED_WIRE_2_0\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__9297\,
            I => \SYNTHESIZED_WIRE_2_0\
        );

    \I__1031\ : InMux
    port map (
            O => \N__9290\,
            I => \N__9287\
        );

    \I__1030\ : LocalMux
    port map (
            O => \N__9287\,
            I => \b2v_inst4.pix_count_int_RNO_0Z0Z_0\
        );

    \I__1029\ : InMux
    port map (
            O => \N__9284\,
            I => \N__9278\
        );

    \I__1028\ : InMux
    port map (
            O => \N__9283\,
            I => \N__9271\
        );

    \I__1027\ : InMux
    port map (
            O => \N__9282\,
            I => \N__9271\
        );

    \I__1026\ : InMux
    port map (
            O => \N__9281\,
            I => \N__9271\
        );

    \I__1025\ : LocalMux
    port map (
            O => \N__9278\,
            I => \SYNTHESIZED_WIRE_2_1\
        );

    \I__1024\ : LocalMux
    port map (
            O => \N__9271\,
            I => \SYNTHESIZED_WIRE_2_1\
        );

    \I__1023\ : InMux
    port map (
            O => \N__9266\,
            I => \b2v_inst4.un1_pix_count_int_cry_0\
        );

    \I__1022\ : CascadeMux
    port map (
            O => \N__9263\,
            I => \N__9259\
        );

    \I__1021\ : InMux
    port map (
            O => \N__9262\,
            I => \N__9252\
        );

    \I__1020\ : InMux
    port map (
            O => \N__9259\,
            I => \N__9252\
        );

    \I__1019\ : InMux
    port map (
            O => \N__9258\,
            I => \N__9249\
        );

    \I__1018\ : InMux
    port map (
            O => \N__9257\,
            I => \N__9246\
        );

    \I__1017\ : LocalMux
    port map (
            O => \N__9252\,
            I => \SYNTHESIZED_WIRE_2_2\
        );

    \I__1016\ : LocalMux
    port map (
            O => \N__9249\,
            I => \SYNTHESIZED_WIRE_2_2\
        );

    \I__1015\ : LocalMux
    port map (
            O => \N__9246\,
            I => \SYNTHESIZED_WIRE_2_2\
        );

    \I__1014\ : InMux
    port map (
            O => \N__9239\,
            I => \b2v_inst4.un1_pix_count_int_cry_1\
        );

    \I__1013\ : InMux
    port map (
            O => \N__9236\,
            I => \N__9230\
        );

    \I__1012\ : InMux
    port map (
            O => \N__9235\,
            I => \N__9223\
        );

    \I__1011\ : InMux
    port map (
            O => \N__9234\,
            I => \N__9223\
        );

    \I__1010\ : InMux
    port map (
            O => \N__9233\,
            I => \N__9223\
        );

    \I__1009\ : LocalMux
    port map (
            O => \N__9230\,
            I => \SYNTHESIZED_WIRE_2_3\
        );

    \I__1008\ : LocalMux
    port map (
            O => \N__9223\,
            I => \SYNTHESIZED_WIRE_2_3\
        );

    \I__1007\ : InMux
    port map (
            O => \N__9218\,
            I => \N__9215\
        );

    \I__1006\ : LocalMux
    port map (
            O => \N__9215\,
            I => \b2v_inst4.pix_count_int_RNO_0Z0Z_3\
        );

    \I__1005\ : InMux
    port map (
            O => \N__9212\,
            I => \b2v_inst4.un1_pix_count_int_cry_2\
        );

    \I__1004\ : InMux
    port map (
            O => \N__9209\,
            I => \N__9203\
        );

    \I__1003\ : InMux
    port map (
            O => \N__9208\,
            I => \N__9196\
        );

    \I__1002\ : InMux
    port map (
            O => \N__9207\,
            I => \N__9196\
        );

    \I__1001\ : InMux
    port map (
            O => \N__9206\,
            I => \N__9196\
        );

    \I__1000\ : LocalMux
    port map (
            O => \N__9203\,
            I => \SYNTHESIZED_WIRE_2_4\
        );

    \I__999\ : LocalMux
    port map (
            O => \N__9196\,
            I => \SYNTHESIZED_WIRE_2_4\
        );

    \I__998\ : InMux
    port map (
            O => \N__9191\,
            I => \b2v_inst4.un1_pix_count_int_cry_3\
        );

    \I__997\ : InMux
    port map (
            O => \N__9188\,
            I => \N__9182\
        );

    \I__996\ : InMux
    port map (
            O => \N__9187\,
            I => \N__9179\
        );

    \I__995\ : InMux
    port map (
            O => \N__9186\,
            I => \N__9174\
        );

    \I__994\ : InMux
    port map (
            O => \N__9185\,
            I => \N__9174\
        );

    \I__993\ : LocalMux
    port map (
            O => \N__9182\,
            I => \SYNTHESIZED_WIRE_2_5\
        );

    \I__992\ : LocalMux
    port map (
            O => \N__9179\,
            I => \SYNTHESIZED_WIRE_2_5\
        );

    \I__991\ : LocalMux
    port map (
            O => \N__9174\,
            I => \SYNTHESIZED_WIRE_2_5\
        );

    \I__990\ : InMux
    port map (
            O => \N__9167\,
            I => \N__9164\
        );

    \I__989\ : LocalMux
    port map (
            O => \N__9164\,
            I => \b2v_inst4.pix_count_int_RNO_0Z0Z_5\
        );

    \I__988\ : InMux
    port map (
            O => \N__9161\,
            I => \b2v_inst4.un1_pix_count_int_cry_4\
        );

    \I__987\ : InMux
    port map (
            O => \N__9158\,
            I => \N__9152\
        );

    \I__986\ : InMux
    port map (
            O => \N__9157\,
            I => \N__9149\
        );

    \I__985\ : InMux
    port map (
            O => \N__9156\,
            I => \N__9144\
        );

    \I__984\ : InMux
    port map (
            O => \N__9155\,
            I => \N__9144\
        );

    \I__983\ : LocalMux
    port map (
            O => \N__9152\,
            I => \SYNTHESIZED_WIRE_2_6\
        );

    \I__982\ : LocalMux
    port map (
            O => \N__9149\,
            I => \SYNTHESIZED_WIRE_2_6\
        );

    \I__981\ : LocalMux
    port map (
            O => \N__9144\,
            I => \SYNTHESIZED_WIRE_2_6\
        );

    \I__980\ : InMux
    port map (
            O => \N__9137\,
            I => \b2v_inst4.un1_pix_count_int_cry_5\
        );

    \I__979\ : InMux
    port map (
            O => \N__9134\,
            I => \N__9131\
        );

    \I__978\ : LocalMux
    port map (
            O => \N__9131\,
            I => \N__9128\
        );

    \I__977\ : Odrv4
    port map (
            O => \N__9128\,
            I => \b2v_inst.N_361\
        );

    \I__976\ : InMux
    port map (
            O => \N__9125\,
            I => \N__9119\
        );

    \I__975\ : InMux
    port map (
            O => \N__9124\,
            I => \N__9119\
        );

    \I__974\ : LocalMux
    port map (
            O => \N__9119\,
            I => \b2v_inst.state_ns_i_i_a2_5Z0Z_6\
        );

    \I__973\ : IoInMux
    port map (
            O => \N__9116\,
            I => \N__9113\
        );

    \I__972\ : LocalMux
    port map (
            O => \N__9113\,
            I => \N__9110\
        );

    \I__971\ : Odrv12
    port map (
            O => \N__9110\,
            I => \b2v_inst.N_254_i\
        );

    \I__970\ : InMux
    port map (
            O => \N__9107\,
            I => \N__9104\
        );

    \I__969\ : LocalMux
    port map (
            O => \N__9104\,
            I => \b2v_inst.pix_count_anteriorZ0Z_2\
        );

    \I__968\ : InMux
    port map (
            O => \N__9101\,
            I => \N__9098\
        );

    \I__967\ : LocalMux
    port map (
            O => \N__9098\,
            I => \b2v_inst.un1_pix_count_anterior_0_I_27_c_RNOZ0\
        );

    \I__966\ : CascadeMux
    port map (
            O => \N__9095\,
            I => \N__9092\
        );

    \I__965\ : InMux
    port map (
            O => \N__9092\,
            I => \N__9089\
        );

    \I__964\ : LocalMux
    port map (
            O => \N__9089\,
            I => \b2v_inst.pix_count_anteriorZ0Z_3\
        );

    \I__963\ : InMux
    port map (
            O => \N__9086\,
            I => \N__9083\
        );

    \I__962\ : LocalMux
    port map (
            O => \N__9083\,
            I => \b2v_inst.pix_count_anteriorZ0Z_10\
        );

    \I__961\ : InMux
    port map (
            O => \N__9080\,
            I => \N__9077\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__9077\,
            I => \b2v_inst.un1_pix_count_anterior_0_I_9_c_RNOZ0\
        );

    \I__959\ : InMux
    port map (
            O => \N__9074\,
            I => \N__9071\
        );

    \I__958\ : LocalMux
    port map (
            O => \N__9071\,
            I => \N__9068\
        );

    \I__957\ : Odrv12
    port map (
            O => \N__9068\,
            I => \b2v_inst.data_a_escribir_RNO_0Z0Z_4\
        );

    \I__956\ : CascadeMux
    port map (
            O => \N__9065\,
            I => \N__9062\
        );

    \I__955\ : InMux
    port map (
            O => \N__9062\,
            I => \N__9059\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__9059\,
            I => \N__9056\
        );

    \I__953\ : Span4Mux_h
    port map (
            O => \N__9056\,
            I => \N__9053\
        );

    \I__952\ : Span4Mux_v
    port map (
            O => \N__9053\,
            I => \N__9050\
        );

    \I__951\ : Odrv4
    port map (
            O => \N__9050\,
            I => \b2v_inst.un1_reg_anterior_iv_0_0_0_4\
        );

    \I__950\ : InMux
    port map (
            O => \N__9047\,
            I => \N__9044\
        );

    \I__949\ : LocalMux
    port map (
            O => \N__9044\,
            I => \N__9041\
        );

    \I__948\ : Span4Mux_h
    port map (
            O => \N__9041\,
            I => \N__9038\
        );

    \I__947\ : Odrv4
    port map (
            O => \N__9038\,
            I => \N_211_i\
        );

    \I__946\ : InMux
    port map (
            O => \N__9035\,
            I => \N__9032\
        );

    \I__945\ : LocalMux
    port map (
            O => \N__9032\,
            I => \N__9029\
        );

    \I__944\ : Span4Mux_h
    port map (
            O => \N__9029\,
            I => \N__9026\
        );

    \I__943\ : Span4Mux_h
    port map (
            O => \N__9026\,
            I => \N__9023\
        );

    \I__942\ : Odrv4
    port map (
            O => \N__9023\,
            I => \N_219_i\
        );

    \I__941\ : InMux
    port map (
            O => \N__9020\,
            I => \N__9017\
        );

    \I__940\ : LocalMux
    port map (
            O => \N__9017\,
            I => \N__9014\
        );

    \I__939\ : Span12Mux_v
    port map (
            O => \N__9014\,
            I => \N__9011\
        );

    \I__938\ : Odrv12
    port map (
            O => \N__9011\,
            I => \N_217_i\
        );

    \I__937\ : InMux
    port map (
            O => \N__9008\,
            I => \N__9005\
        );

    \I__936\ : LocalMux
    port map (
            O => \N__9005\,
            I => \N__9002\
        );

    \I__935\ : Span4Mux_h
    port map (
            O => \N__9002\,
            I => \N__8999\
        );

    \I__934\ : Span4Mux_v
    port map (
            O => \N__8999\,
            I => \N__8996\
        );

    \I__933\ : Odrv4
    port map (
            O => \N__8996\,
            I => \N_215_i\
        );

    \I__932\ : CascadeMux
    port map (
            O => \N__8993\,
            I => \N__8990\
        );

    \I__931\ : InMux
    port map (
            O => \N__8990\,
            I => \N__8987\
        );

    \I__930\ : LocalMux
    port map (
            O => \N__8987\,
            I => \b2v_inst.state_ns_i_i_a2_4Z0Z_6\
        );

    \I__929\ : CascadeMux
    port map (
            O => \N__8984\,
            I => \b2v_inst.state_ns_i_i_a2_4Z0Z_6_cascade_\
        );

    \I__928\ : CascadeMux
    port map (
            O => \N__8981\,
            I => \b2v_inst.N_497_cascade_\
        );

    \I__927\ : InMux
    port map (
            O => \N__8978\,
            I => \N__8975\
        );

    \I__926\ : LocalMux
    port map (
            O => \N__8975\,
            I => \b2v_inst.N_317\
        );

    \I__925\ : InMux
    port map (
            O => \N__8972\,
            I => \N__8969\
        );

    \I__924\ : LocalMux
    port map (
            O => \N__8969\,
            I => \b2v_inst.un1_reg_anterior_iv_0_0_a2_4_tz_1_2\
        );

    \I__923\ : InMux
    port map (
            O => \N__8966\,
            I => \N__8963\
        );

    \I__922\ : LocalMux
    port map (
            O => \N__8963\,
            I => \N__8960\
        );

    \I__921\ : Span4Mux_v
    port map (
            O => \N__8960\,
            I => \N__8956\
        );

    \I__920\ : InMux
    port map (
            O => \N__8959\,
            I => \N__8953\
        );

    \I__919\ : Odrv4
    port map (
            O => \N__8956\,
            I => \b2v_inst.eventosZ0Z_2\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__8953\,
            I => \b2v_inst.eventosZ0Z_2\
        );

    \I__917\ : CascadeMux
    port map (
            O => \N__8948\,
            I => \b2v_inst.N_320_tz_cascade_\
        );

    \I__916\ : CascadeMux
    port map (
            O => \N__8945\,
            I => \b2v_inst.un1_m3_0_m3_ns_1_cascade_\
        );

    \I__915\ : InMux
    port map (
            O => \N__8942\,
            I => \N__8939\
        );

    \I__914\ : LocalMux
    port map (
            O => \N__8939\,
            I => \N__8936\
        );

    \I__913\ : Odrv4
    port map (
            O => \N__8936\,
            I => \b2v_inst.N_318\
        );

    \I__912\ : CascadeMux
    port map (
            O => \N__8933\,
            I => \b2v_inst.data_a_escribir_RNO_3Z0Z_4_cascade_\
        );

    \I__911\ : CascadeMux
    port map (
            O => \N__8930\,
            I => \b2v_inst.data_a_escribir_RNO_3Z0Z_0_cascade_\
        );

    \I__910\ : InMux
    port map (
            O => \N__8927\,
            I => \N__8924\
        );

    \I__909\ : LocalMux
    port map (
            O => \N__8924\,
            I => \N__8921\
        );

    \I__908\ : Span4Mux_v
    port map (
            O => \N__8921\,
            I => \N__8918\
        );

    \I__907\ : Odrv4
    port map (
            O => \N__8918\,
            I => \b2v_inst.un1_reg_anterior_iv_0_0_0_0\
        );

    \I__906\ : InMux
    port map (
            O => \N__8915\,
            I => \N__8912\
        );

    \I__905\ : LocalMux
    port map (
            O => \N__8912\,
            I => \b2v_inst.un1_m3_2_0\
        );

    \I__904\ : CascadeMux
    port map (
            O => \N__8909\,
            I => \b2v_inst.data_a_escribir_RNO_1Z0Z_0_cascade_\
        );

    \I__903\ : InMux
    port map (
            O => \N__8906\,
            I => \N__8903\
        );

    \I__902\ : LocalMux
    port map (
            O => \N__8903\,
            I => \N__8900\
        );

    \I__901\ : Odrv4
    port map (
            O => \N__8900\,
            I => \b2v_inst.un1_reg_anterior_iv_0_0_1_1_3\
        );

    \I__900\ : CascadeMux
    port map (
            O => \N__8897\,
            I => \b2v_inst.N_315_cascade_\
        );

    \I__899\ : InMux
    port map (
            O => \N__8894\,
            I => \N__8891\
        );

    \I__898\ : LocalMux
    port map (
            O => \N__8891\,
            I => \b2v_inst.un1_reg_anterior_iv_0_0_1_3\
        );

    \I__897\ : CascadeMux
    port map (
            O => \N__8888\,
            I => \b2v_inst.un1_reg_anterior_iv_0_0_a2_6_0_1_cascade_\
        );

    \I__896\ : InMux
    port map (
            O => \N__8885\,
            I => \N__8873\
        );

    \I__895\ : InMux
    port map (
            O => \N__8884\,
            I => \N__8873\
        );

    \I__894\ : InMux
    port map (
            O => \N__8883\,
            I => \N__8860\
        );

    \I__893\ : InMux
    port map (
            O => \N__8882\,
            I => \N__8860\
        );

    \I__892\ : InMux
    port map (
            O => \N__8881\,
            I => \N__8860\
        );

    \I__891\ : InMux
    port map (
            O => \N__8880\,
            I => \N__8860\
        );

    \I__890\ : InMux
    port map (
            O => \N__8879\,
            I => \N__8860\
        );

    \I__889\ : InMux
    port map (
            O => \N__8878\,
            I => \N__8860\
        );

    \I__888\ : LocalMux
    port map (
            O => \N__8873\,
            I => \N__8855\
        );

    \I__887\ : LocalMux
    port map (
            O => \N__8860\,
            I => \N__8855\
        );

    \I__886\ : Odrv4
    port map (
            O => \N__8855\,
            I => \b2v_inst.ignorar_anchoZ0Z_1\
        );

    \I__885\ : CascadeMux
    port map (
            O => \N__8852\,
            I => \N__8849\
        );

    \I__884\ : InMux
    port map (
            O => \N__8849\,
            I => \N__8846\
        );

    \I__883\ : LocalMux
    port map (
            O => \N__8846\,
            I => \b2v_inst.pix_count_anteriorZ0Z_7\
        );

    \I__882\ : InMux
    port map (
            O => \N__8843\,
            I => \N__8840\
        );

    \I__881\ : LocalMux
    port map (
            O => \N__8840\,
            I => \b2v_inst.pix_count_anteriorZ0Z_8\
        );

    \I__880\ : InMux
    port map (
            O => \N__8837\,
            I => \N__8834\
        );

    \I__879\ : LocalMux
    port map (
            O => \N__8834\,
            I => \N__8831\
        );

    \I__878\ : Odrv12
    port map (
            O => \N__8831\,
            I => \b2v_inst.un1_pix_count_anterior_0_I_51_c_RNOZ0\
        );

    \I__877\ : CascadeMux
    port map (
            O => \N__8828\,
            I => \N__8825\
        );

    \I__876\ : InMux
    port map (
            O => \N__8825\,
            I => \N__8822\
        );

    \I__875\ : LocalMux
    port map (
            O => \N__8822\,
            I => \b2v_inst.pix_count_anteriorZ0Z_9\
        );

    \I__874\ : CEMux
    port map (
            O => \N__8819\,
            I => \N__8816\
        );

    \I__873\ : LocalMux
    port map (
            O => \N__8816\,
            I => \N__8813\
        );

    \I__872\ : Span4Mux_v
    port map (
            O => \N__8813\,
            I => \N__8810\
        );

    \I__871\ : Odrv4
    port map (
            O => \N__8810\,
            I => \b2v_inst.un1_state_17_0\
        );

    \I__870\ : InMux
    port map (
            O => \N__8807\,
            I => \N__8804\
        );

    \I__869\ : LocalMux
    port map (
            O => \N__8804\,
            I => \b2v_inst.pix_count_anteriorZ0Z_12\
        );

    \I__868\ : InMux
    port map (
            O => \N__8801\,
            I => \N__8798\
        );

    \I__867\ : LocalMux
    port map (
            O => \N__8798\,
            I => \N__8795\
        );

    \I__866\ : Odrv4
    port map (
            O => \N__8795\,
            I => \b2v_inst.un1_pix_count_anterior_0_I_39_c_RNOZ0\
        );

    \I__865\ : InMux
    port map (
            O => \N__8792\,
            I => \N__8789\
        );

    \I__864\ : LocalMux
    port map (
            O => \N__8789\,
            I => \N__8786\
        );

    \I__863\ : Odrv4
    port map (
            O => \N__8786\,
            I => \b2v_inst.un1_pix_count_anterior_0_I_21_c_RNOZ0\
        );

    \I__862\ : InMux
    port map (
            O => \N__8783\,
            I => \N__8780\
        );

    \I__861\ : LocalMux
    port map (
            O => \N__8780\,
            I => \b2v_inst.pix_count_anteriorZ0Z_6\
        );

    \I__860\ : CascadeMux
    port map (
            O => \N__8777\,
            I => \b2v_inst4.un1_pix_count_int_0_sqmuxa_8_cascade_\
        );

    \I__859\ : InMux
    port map (
            O => \N__8774\,
            I => \N__8771\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__8771\,
            I => \b2v_inst.pix_count_anteriorZ0Z_4\
        );

    \I__857\ : CascadeMux
    port map (
            O => \N__8768\,
            I => \N__8765\
        );

    \I__856\ : InMux
    port map (
            O => \N__8765\,
            I => \N__8762\
        );

    \I__855\ : LocalMux
    port map (
            O => \N__8762\,
            I => \b2v_inst.pix_count_anteriorZ0Z_5\
        );

    \I__854\ : CascadeMux
    port map (
            O => \N__8759\,
            I => \N__8756\
        );

    \I__853\ : InMux
    port map (
            O => \N__8756\,
            I => \N__8753\
        );

    \I__852\ : LocalMux
    port map (
            O => \N__8753\,
            I => \b2v_inst.pix_count_anteriorZ0Z_1\
        );

    \I__851\ : InMux
    port map (
            O => \N__8750\,
            I => \N__8747\
        );

    \I__850\ : LocalMux
    port map (
            O => \N__8747\,
            I => \b2v_inst.un1_pix_count_anterior_0_I_1_c_RNOZ0\
        );

    \I__849\ : InMux
    port map (
            O => \N__8744\,
            I => \N__8741\
        );

    \I__848\ : LocalMux
    port map (
            O => \N__8741\,
            I => \b2v_inst.pix_count_anteriorZ0Z_0\
        );

    \I__847\ : InMux
    port map (
            O => \N__8738\,
            I => \b2v_inst.un1_pix_count_anterior_0_N_2\
        );

    \I__846\ : InMux
    port map (
            O => \N__8735\,
            I => \N__8732\
        );

    \I__845\ : LocalMux
    port map (
            O => \N__8732\,
            I => \b2v_inst.un1_pix_count_anterior_0_I_15_c_RNOZ0\
        );

    \I__844\ : InMux
    port map (
            O => \N__8729\,
            I => \bfn_1_20_0_\
        );

    \I__843\ : InMux
    port map (
            O => \N__8726\,
            I => \N__8723\
        );

    \I__842\ : LocalMux
    port map (
            O => \N__8723\,
            I => \N__8720\
        );

    \I__841\ : Span12Mux_v
    port map (
            O => \N__8720\,
            I => \N__8717\
        );

    \I__840\ : Odrv12
    port map (
            O => \N__8717\,
            I => \b2v_inst.g0_10_1\
        );

    \I__839\ : InMux
    port map (
            O => \N__8714\,
            I => \N__8711\
        );

    \I__838\ : LocalMux
    port map (
            O => \N__8711\,
            I => \N__8708\
        );

    \I__837\ : Span12Mux_s8_v
    port map (
            O => \N__8708\,
            I => \N__8705\
        );

    \I__836\ : Odrv12
    port map (
            O => \N__8705\,
            I => \b2v_inst.g0_10_a3_7\
        );

    \I__835\ : CascadeMux
    port map (
            O => \N__8702\,
            I => \N__8699\
        );

    \I__834\ : InMux
    port map (
            O => \N__8699\,
            I => \N__8696\
        );

    \I__833\ : LocalMux
    port map (
            O => \N__8696\,
            I => \b2v_inst.reg_ancho_1_i_4\
        );

    \I__832\ : CascadeMux
    port map (
            O => \N__8693\,
            I => \N__8690\
        );

    \I__831\ : InMux
    port map (
            O => \N__8690\,
            I => \N__8687\
        );

    \I__830\ : LocalMux
    port map (
            O => \N__8687\,
            I => \b2v_inst.reg_ancho_1_i_5\
        );

    \I__829\ : CascadeMux
    port map (
            O => \N__8684\,
            I => \N__8681\
        );

    \I__828\ : InMux
    port map (
            O => \N__8681\,
            I => \N__8678\
        );

    \I__827\ : LocalMux
    port map (
            O => \N__8678\,
            I => \b2v_inst.reg_ancho_1_i_6\
        );

    \I__826\ : CascadeMux
    port map (
            O => \N__8675\,
            I => \N__8672\
        );

    \I__825\ : InMux
    port map (
            O => \N__8672\,
            I => \N__8669\
        );

    \I__824\ : LocalMux
    port map (
            O => \N__8669\,
            I => \b2v_inst.reg_ancho_1_i_7\
        );

    \I__823\ : InMux
    port map (
            O => \N__8666\,
            I => \bfn_1_18_0_\
        );

    \I__822\ : CascadeMux
    port map (
            O => \N__8663\,
            I => \N__8659\
        );

    \I__821\ : InMux
    port map (
            O => \N__8662\,
            I => \N__8656\
        );

    \I__820\ : InMux
    port map (
            O => \N__8659\,
            I => \N__8653\
        );

    \I__819\ : LocalMux
    port map (
            O => \N__8656\,
            I => \b2v_inst.eventosZ0Z_3\
        );

    \I__818\ : LocalMux
    port map (
            O => \N__8653\,
            I => \b2v_inst.eventosZ0Z_3\
        );

    \I__817\ : InMux
    port map (
            O => \N__8648\,
            I => \N__8644\
        );

    \I__816\ : InMux
    port map (
            O => \N__8647\,
            I => \N__8641\
        );

    \I__815\ : LocalMux
    port map (
            O => \N__8644\,
            I => \b2v_inst.eventosZ0Z_4\
        );

    \I__814\ : LocalMux
    port map (
            O => \N__8641\,
            I => \b2v_inst.eventosZ0Z_4\
        );

    \I__813\ : InMux
    port map (
            O => \N__8636\,
            I => \N__8632\
        );

    \I__812\ : InMux
    port map (
            O => \N__8635\,
            I => \N__8629\
        );

    \I__811\ : LocalMux
    port map (
            O => \N__8632\,
            I => \b2v_inst.eventosZ0Z_0\
        );

    \I__810\ : LocalMux
    port map (
            O => \N__8629\,
            I => \b2v_inst.eventosZ0Z_0\
        );

    \I__809\ : InMux
    port map (
            O => \N__8624\,
            I => \N__8620\
        );

    \I__808\ : InMux
    port map (
            O => \N__8623\,
            I => \N__8617\
        );

    \I__807\ : LocalMux
    port map (
            O => \N__8620\,
            I => \b2v_inst.eventosZ0Z_5\
        );

    \I__806\ : LocalMux
    port map (
            O => \N__8617\,
            I => \b2v_inst.eventosZ0Z_5\
        );

    \I__805\ : CEMux
    port map (
            O => \N__8612\,
            I => \N__8609\
        );

    \I__804\ : LocalMux
    port map (
            O => \N__8609\,
            I => \N__8606\
        );

    \I__803\ : Odrv4
    port map (
            O => \N__8606\,
            I => \b2v_inst.N_47_i\
        );

    \I__802\ : CascadeMux
    port map (
            O => \N__8603\,
            I => \N__8600\
        );

    \I__801\ : InMux
    port map (
            O => \N__8600\,
            I => \N__8597\
        );

    \I__800\ : LocalMux
    port map (
            O => \N__8597\,
            I => \b2v_inst.reg_ancho_1_i_0\
        );

    \I__799\ : CascadeMux
    port map (
            O => \N__8594\,
            I => \N__8591\
        );

    \I__798\ : InMux
    port map (
            O => \N__8591\,
            I => \N__8588\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__8588\,
            I => \b2v_inst.reg_ancho_1_i_1\
        );

    \I__796\ : CascadeMux
    port map (
            O => \N__8585\,
            I => \N__8582\
        );

    \I__795\ : InMux
    port map (
            O => \N__8582\,
            I => \N__8579\
        );

    \I__794\ : LocalMux
    port map (
            O => \N__8579\,
            I => \b2v_inst.reg_ancho_1_i_2\
        );

    \I__793\ : CascadeMux
    port map (
            O => \N__8576\,
            I => \N__8573\
        );

    \I__792\ : InMux
    port map (
            O => \N__8573\,
            I => \N__8570\
        );

    \I__791\ : LocalMux
    port map (
            O => \N__8570\,
            I => \N__8567\
        );

    \I__790\ : Odrv4
    port map (
            O => \N__8567\,
            I => \b2v_inst.reg_ancho_1_i_3\
        );

    \I__789\ : InMux
    port map (
            O => \N__8564\,
            I => \b2v_inst.eventos_cry_0\
        );

    \I__788\ : InMux
    port map (
            O => \N__8561\,
            I => \b2v_inst.eventos_cry_1\
        );

    \I__787\ : InMux
    port map (
            O => \N__8558\,
            I => \b2v_inst.eventos_cry_2\
        );

    \I__786\ : InMux
    port map (
            O => \N__8555\,
            I => \b2v_inst.eventos_cry_3\
        );

    \I__785\ : InMux
    port map (
            O => \N__8552\,
            I => \b2v_inst.eventos_cry_4\
        );

    \I__784\ : InMux
    port map (
            O => \N__8549\,
            I => \b2v_inst.eventos_cry_5\
        );

    \I__783\ : InMux
    port map (
            O => \N__8546\,
            I => \b2v_inst.eventos_cry_6\
        );

    \I__782\ : CascadeMux
    port map (
            O => \N__8543\,
            I => \N__8539\
        );

    \I__781\ : CascadeMux
    port map (
            O => \N__8542\,
            I => \N__8536\
        );

    \I__780\ : InMux
    port map (
            O => \N__8539\,
            I => \N__8526\
        );

    \I__779\ : InMux
    port map (
            O => \N__8536\,
            I => \N__8526\
        );

    \I__778\ : InMux
    port map (
            O => \N__8535\,
            I => \N__8526\
        );

    \I__777\ : InMux
    port map (
            O => \N__8534\,
            I => \N__8521\
        );

    \I__776\ : InMux
    port map (
            O => \N__8533\,
            I => \N__8521\
        );

    \I__775\ : LocalMux
    port map (
            O => \N__8526\,
            I => \b2v_inst.cuenta_pixelZ0Z_7\
        );

    \I__774\ : LocalMux
    port map (
            O => \N__8521\,
            I => \b2v_inst.cuenta_pixelZ0Z_7\
        );

    \I__773\ : InMux
    port map (
            O => \N__8516\,
            I => \N__8513\
        );

    \I__772\ : LocalMux
    port map (
            O => \N__8513\,
            I => \N__8505\
        );

    \I__771\ : InMux
    port map (
            O => \N__8512\,
            I => \N__8496\
        );

    \I__770\ : InMux
    port map (
            O => \N__8511\,
            I => \N__8496\
        );

    \I__769\ : InMux
    port map (
            O => \N__8510\,
            I => \N__8496\
        );

    \I__768\ : InMux
    port map (
            O => \N__8509\,
            I => \N__8496\
        );

    \I__767\ : InMux
    port map (
            O => \N__8508\,
            I => \N__8493\
        );

    \I__766\ : Odrv4
    port map (
            O => \N__8505\,
            I => \b2v_inst.cuenta_pixelZ0Z_2\
        );

    \I__765\ : LocalMux
    port map (
            O => \N__8496\,
            I => \b2v_inst.cuenta_pixelZ0Z_2\
        );

    \I__764\ : LocalMux
    port map (
            O => \N__8493\,
            I => \b2v_inst.cuenta_pixelZ0Z_2\
        );

    \I__763\ : InMux
    port map (
            O => \N__8486\,
            I => \N__8483\
        );

    \I__762\ : LocalMux
    port map (
            O => \N__8483\,
            I => \b2v_inst.N_6_i\
        );

    \I__761\ : CascadeMux
    port map (
            O => \N__8480\,
            I => \b2v_inst.g0_6_1_cascade_\
        );

    \I__760\ : InMux
    port map (
            O => \N__8477\,
            I => \N__8474\
        );

    \I__759\ : LocalMux
    port map (
            O => \N__8474\,
            I => \N__8471\
        );

    \I__758\ : Odrv4
    port map (
            O => \N__8471\,
            I => \b2v_inst.N_4\
        );

    \I__757\ : CascadeMux
    port map (
            O => \N__8468\,
            I => \b2v_inst.un11_cuenta_pixel_6_cascade_\
        );

    \I__756\ : InMux
    port map (
            O => \N__8465\,
            I => \N__8462\
        );

    \I__755\ : LocalMux
    port map (
            O => \N__8462\,
            I => \N__8457\
        );

    \I__754\ : InMux
    port map (
            O => \N__8461\,
            I => \N__8452\
        );

    \I__753\ : InMux
    port map (
            O => \N__8460\,
            I => \N__8452\
        );

    \I__752\ : Odrv4
    port map (
            O => \N__8457\,
            I => \b2v_inst.un11_cuenta_pixel_6\
        );

    \I__751\ : LocalMux
    port map (
            O => \N__8452\,
            I => \b2v_inst.un11_cuenta_pixel_6\
        );

    \I__750\ : InMux
    port map (
            O => \N__8447\,
            I => \N__8441\
        );

    \I__749\ : InMux
    port map (
            O => \N__8446\,
            I => \N__8436\
        );

    \I__748\ : InMux
    port map (
            O => \N__8445\,
            I => \N__8436\
        );

    \I__747\ : InMux
    port map (
            O => \N__8444\,
            I => \N__8433\
        );

    \I__746\ : LocalMux
    port map (
            O => \N__8441\,
            I => \b2v_inst.cuenta_pixel_RNI3FD32_0Z0Z_5\
        );

    \I__745\ : LocalMux
    port map (
            O => \N__8436\,
            I => \b2v_inst.cuenta_pixel_RNI3FD32_0Z0Z_5\
        );

    \I__744\ : LocalMux
    port map (
            O => \N__8433\,
            I => \b2v_inst.cuenta_pixel_RNI3FD32_0Z0Z_5\
        );

    \I__743\ : InMux
    port map (
            O => \N__8426\,
            I => \N__8420\
        );

    \I__742\ : InMux
    port map (
            O => \N__8425\,
            I => \N__8415\
        );

    \I__741\ : InMux
    port map (
            O => \N__8424\,
            I => \N__8415\
        );

    \I__740\ : InMux
    port map (
            O => \N__8423\,
            I => \N__8408\
        );

    \I__739\ : LocalMux
    port map (
            O => \N__8420\,
            I => \N__8403\
        );

    \I__738\ : LocalMux
    port map (
            O => \N__8415\,
            I => \N__8403\
        );

    \I__737\ : InMux
    port map (
            O => \N__8414\,
            I => \N__8394\
        );

    \I__736\ : InMux
    port map (
            O => \N__8413\,
            I => \N__8394\
        );

    \I__735\ : InMux
    port map (
            O => \N__8412\,
            I => \N__8394\
        );

    \I__734\ : InMux
    port map (
            O => \N__8411\,
            I => \N__8394\
        );

    \I__733\ : LocalMux
    port map (
            O => \N__8408\,
            I => \b2v_inst.cuenta_pixelZ0Z_3\
        );

    \I__732\ : Odrv4
    port map (
            O => \N__8403\,
            I => \b2v_inst.cuenta_pixelZ0Z_3\
        );

    \I__731\ : LocalMux
    port map (
            O => \N__8394\,
            I => \b2v_inst.cuenta_pixelZ0Z_3\
        );

    \I__730\ : InMux
    port map (
            O => \N__8387\,
            I => \N__8383\
        );

    \I__729\ : InMux
    port map (
            O => \N__8386\,
            I => \N__8380\
        );

    \I__728\ : LocalMux
    port map (
            O => \N__8383\,
            I => \N__8373\
        );

    \I__727\ : LocalMux
    port map (
            O => \N__8380\,
            I => \N__8373\
        );

    \I__726\ : InMux
    port map (
            O => \N__8379\,
            I => \N__8368\
        );

    \I__725\ : InMux
    port map (
            O => \N__8378\,
            I => \N__8368\
        );

    \I__724\ : Odrv4
    port map (
            O => \N__8373\,
            I => \b2v_inst.un1_cuenta_pixel_c3\
        );

    \I__723\ : LocalMux
    port map (
            O => \N__8368\,
            I => \b2v_inst.un1_cuenta_pixel_c3\
        );

    \I__722\ : CascadeMux
    port map (
            O => \N__8363\,
            I => \N__8359\
        );

    \I__721\ : CascadeMux
    port map (
            O => \N__8362\,
            I => \N__8356\
        );

    \I__720\ : InMux
    port map (
            O => \N__8359\,
            I => \N__8341\
        );

    \I__719\ : InMux
    port map (
            O => \N__8356\,
            I => \N__8341\
        );

    \I__718\ : InMux
    port map (
            O => \N__8355\,
            I => \N__8341\
        );

    \I__717\ : InMux
    port map (
            O => \N__8354\,
            I => \N__8341\
        );

    \I__716\ : InMux
    port map (
            O => \N__8353\,
            I => \N__8338\
        );

    \I__715\ : InMux
    port map (
            O => \N__8352\,
            I => \N__8331\
        );

    \I__714\ : InMux
    port map (
            O => \N__8351\,
            I => \N__8331\
        );

    \I__713\ : InMux
    port map (
            O => \N__8350\,
            I => \N__8331\
        );

    \I__712\ : LocalMux
    port map (
            O => \N__8341\,
            I => \N__8328\
        );

    \I__711\ : LocalMux
    port map (
            O => \N__8338\,
            I => \b2v_inst.cuenta_pixelZ0Z_4\
        );

    \I__710\ : LocalMux
    port map (
            O => \N__8331\,
            I => \b2v_inst.cuenta_pixelZ0Z_4\
        );

    \I__709\ : Odrv4
    port map (
            O => \N__8328\,
            I => \b2v_inst.cuenta_pixelZ0Z_4\
        );

    \I__708\ : InMux
    port map (
            O => \N__8321\,
            I => \bfn_1_15_0_\
        );

    \I__707\ : CascadeMux
    port map (
            O => \N__8318\,
            I => \b2v_inst.g0_10_a3_0_7_cascade_\
        );

    \I__706\ : InMux
    port map (
            O => \N__8315\,
            I => \N__8312\
        );

    \I__705\ : LocalMux
    port map (
            O => \N__8312\,
            I => \b2v_inst.g0_10_a3_0_5\
        );

    \I__704\ : CascadeMux
    port map (
            O => \N__8309\,
            I => \b2v_inst.g0_10_a3_5_cascade_\
        );

    \I__703\ : InMux
    port map (
            O => \N__8306\,
            I => \N__8303\
        );

    \I__702\ : LocalMux
    port map (
            O => \N__8303\,
            I => \b2v_inst.g0_10_a3_4\
        );

    \I__701\ : InMux
    port map (
            O => \N__8300\,
            I => \N__8297\
        );

    \I__700\ : LocalMux
    port map (
            O => \N__8297\,
            I => \b2v_inst.un1_cuenta_pixel_c6\
        );

    \I__699\ : CascadeMux
    port map (
            O => \N__8294\,
            I => \b2v_inst.un1_cuenta_pixel_c6_cascade_\
        );

    \I__698\ : InMux
    port map (
            O => \N__8291\,
            I => \N__8288\
        );

    \I__697\ : LocalMux
    port map (
            O => \N__8288\,
            I => \b2v_inst.cuenta_pixel_RNO_0Z0Z_1\
        );

    \I__696\ : InMux
    port map (
            O => \N__8285\,
            I => \N__8282\
        );

    \I__695\ : LocalMux
    port map (
            O => \N__8282\,
            I => \b2v_inst.g0_10_a3_0_4\
        );

    \IN_MUX_bfv_2_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_11_0_\
        );

    \IN_MUX_bfv_1_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_19_0_\
        );

    \IN_MUX_bfv_1_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst.valor_max_final53\,
            carryinitout => \bfn_1_20_0_\
        );

    \IN_MUX_bfv_5_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_19_0_\
        );

    \IN_MUX_bfv_5_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst.valor_max_final52\,
            carryinitout => \bfn_5_20_0_\
        );

    \IN_MUX_bfv_6_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_17_0_\
        );

    \IN_MUX_bfv_6_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst.un3_valor_max2\,
            carryinitout => \bfn_6_18_0_\
        );

    \IN_MUX_bfv_10_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_10_0_\
        );

    \IN_MUX_bfv_3_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_15_0_\
        );

    \IN_MUX_bfv_3_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst.data_a_escribir10\,
            carryinitout => \bfn_3_16_0_\
        );

    \IN_MUX_bfv_3_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_13_0_\
        );

    \IN_MUX_bfv_3_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst4.un1_pix_count_int_cry_7\,
            carryinitout => \bfn_3_14_0_\
        );

    \IN_MUX_bfv_1_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_15_0_\
        );

    \IN_MUX_bfv_3_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_19_0_\
        );

    \IN_MUX_bfv_3_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst.valor_max_final51\,
            carryinitout => \bfn_3_20_0_\
        );

    \IN_MUX_bfv_5_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_17_0_\
        );

    \IN_MUX_bfv_5_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst.valor_max_final50\,
            carryinitout => \bfn_5_18_0_\
        );

    \IN_MUX_bfv_1_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_17_0_\
        );

    \IN_MUX_bfv_1_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst.un3_valor_max1\,
            carryinitout => \bfn_1_18_0_\
        );

    \reset_i_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__13151\,
            GLOBALBUFFEROUTPUT => reset_i_g
        );

    \b2v_inst.un1_pix_count_anterior_0_I_39_c_RNIT6R7_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__9116\,
            GLOBALBUFFEROUTPUT => \b2v_inst.N_254_i_g\
        );

    \b2v_inst.state_RNI0PU5_2\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__10171\,
            GLOBALBUFFEROUTPUT => \b2v_inst.state_g_2\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \b2v_inst.cuenta_pixel_1_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010001010101010"
        )
    port map (
            in0 => \N__8291\,
            in1 => \N__8465\,
            in2 => \N__11801\,
            in3 => \N__8447\,
            lcout => \b2v_inst.cuenta_pixelZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22410\,
            ce => \N__9336\,
            sr => \N__22875\
        );

    \b2v_inst.ignorar_ancho_1_RNO_1_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__8509\,
            in1 => \N__12422\,
            in2 => \N__11846\,
            in3 => \N__12493\,
            lcout => \b2v_inst.g0_10_a3_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.cuenta_pixel_2_LC_1_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__12497\,
            in1 => \_gnd_net_\,
            in2 => \N__12438\,
            in3 => \N__8511\,
            lcout => \b2v_inst.cuenta_pixelZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22410\,
            ce => \N__9336\,
            sr => \N__22875\
        );

    \b2v_inst.cuenta_pixel_RNITIM11_2_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__12494\,
            in1 => \_gnd_net_\,
            in2 => \N__12437\,
            in3 => \N__8510\,
            lcout => \b2v_inst.un1_cuenta_pixel_c3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.cuenta_pixel_RNIT0FM_1_LC_1_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12426\,
            in2 => \_gnd_net_\,
            in3 => \N__12495\,
            lcout => \b2v_inst.N_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.cuenta_pixel_3_LC_1_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__12498\,
            in1 => \N__8423\,
            in2 => \N__12439\,
            in3 => \N__8512\,
            lcout => \b2v_inst.cuenta_pixelZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22410\,
            ce => \N__9336\,
            sr => \N__22875\
        );

    \b2v_inst.cuenta_pixel_RNO_0_1_LC_1_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12427\,
            in2 => \_gnd_net_\,
            in3 => \N__12496\,
            lcout => \b2v_inst.cuenta_pixel_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.ignorar_ancho_1_RNO_0_LC_1_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__8315\,
            in1 => \N__8285\,
            in2 => \_gnd_net_\,
            in3 => \N__10210\,
            lcout => OPEN,
            ltout => \b2v_inst.g0_10_a3_0_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.ignorar_ancho_1_RNO_LC_1_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010001000100"
        )
    port map (
            in0 => \N__15677\,
            in1 => \N__10164\,
            in2 => \N__8318\,
            in3 => \N__8444\,
            lcout => \b2v_inst.un1_state_17_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.cuenta_pixel_RNI3FD32_0_5_LC_1_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__8413\,
            in1 => \N__11759\,
            in2 => \N__8362\,
            in3 => \N__8378\,
            lcout => \b2v_inst.cuenta_pixel_RNI3FD32_0Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.ignorar_ancho_1_RNO_2_LC_1_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__8533\,
            in1 => \N__8354\,
            in2 => \N__15685\,
            in3 => \N__8411\,
            lcout => \b2v_inst.g0_10_a3_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.ignorar_anterior_RNO_0_LC_1_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__8414\,
            in1 => \N__11760\,
            in2 => \N__8363\,
            in3 => \N__8379\,
            lcout => \b2v_inst.g0_10_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.ignorar_anterior_RNO_3_LC_1_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__8534\,
            in1 => \N__8355\,
            in2 => \N__15686\,
            in3 => \N__8412\,
            lcout => OPEN,
            ltout => \b2v_inst.g0_10_a3_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.ignorar_anterior_RNO_1_LC_1_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8306\,
            in2 => \N__8309\,
            in3 => \N__10209\,
            lcout => \b2v_inst.g0_10_a3_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.ignorar_anterior_RNO_2_LC_1_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__8508\,
            in1 => \N__12421\,
            in2 => \N__11845\,
            in3 => \N__12473\,
            lcout => \b2v_inst.g0_10_a3_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.cuenta_pixel_7_LC_1_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101101011110000"
        )
    port map (
            in0 => \N__11834\,
            in1 => \_gnd_net_\,
            in2 => \N__8543\,
            in3 => \N__8300\,
            lcout => \b2v_inst.cuenta_pixelZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22562\,
            ce => \N__9337\,
            sr => \N__22876\
        );

    \b2v_inst.cuenta_pixel_RNI3FD32_5_LC_1_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8351\,
            in1 => \N__8386\,
            in2 => \N__11764\,
            in3 => \N__8425\,
            lcout => \b2v_inst.un1_cuenta_pixel_c6\,
            ltout => \b2v_inst.un1_cuenta_pixel_c6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.cuenta_pixel_6_LC_1_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001001001011010"
        )
    port map (
            in0 => \N__11833\,
            in1 => \N__12395\,
            in2 => \N__8294\,
            in3 => \N__8461\,
            lcout => \b2v_inst.cuenta_pixelZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22562\,
            ce => \N__9337\,
            sr => \N__22876\
        );

    \b2v_inst.cuenta_pixel_RNIC2N11_5_LC_1_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100100110011"
        )
    port map (
            in0 => \N__11755\,
            in1 => \N__8535\,
            in2 => \_gnd_net_\,
            in3 => \N__11832\,
            lcout => \b2v_inst.N_6_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.cuenta_pixel_RNI8GUC1_7_LC_1_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011001101"
        )
    port map (
            in0 => \N__8424\,
            in1 => \N__8350\,
            in2 => \N__8542\,
            in3 => \N__8516\,
            lcout => OPEN,
            ltout => \b2v_inst.g0_6_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.cuenta_pixel_RNIJ7CG3_4_LC_1_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000001000"
        )
    port map (
            in0 => \N__8352\,
            in1 => \N__8486\,
            in2 => \N__8480\,
            in3 => \N__8477\,
            lcout => \b2v_inst.un11_cuenta_pixel_6\,
            ltout => \b2v_inst.un11_cuenta_pixel_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.cuenta_pixel_5_LC_1_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000001010"
        )
    port map (
            in0 => \N__8446\,
            in1 => \_gnd_net_\,
            in2 => \N__8468\,
            in3 => \N__11787\,
            lcout => \b2v_inst.cuenta_pixelZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22562\,
            ce => \N__9337\,
            sr => \N__22876\
        );

    \b2v_inst.cuenta_pixel_0_LC_1_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000100011111111"
        )
    port map (
            in0 => \N__8460\,
            in1 => \N__8445\,
            in2 => \N__11794\,
            in3 => \N__12492\,
            lcout => \b2v_inst.cuenta_pixelZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22562\,
            ce => \N__9337\,
            sr => \N__22876\
        );

    \b2v_inst.cuenta_pixel_4_LC_1_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__8353\,
            in1 => \N__8426\,
            in2 => \_gnd_net_\,
            in3 => \N__8387\,
            lcout => \b2v_inst.cuenta_pixelZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22598\,
            ce => \N__9339\,
            sr => \N__22879\
        );

    \b2v_inst.pix_count_anterior_12_LC_1_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9397\,
            lcout => \b2v_inst.pix_count_anteriorZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22598\,
            ce => \N__9339\,
            sr => \N__22879\
        );

    \b2v_inst.eventos_0_LC_1_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1011",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8635\,
            in2 => \_gnd_net_\,
            in3 => \N__8321\,
            lcout => \b2v_inst.eventosZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_1_15_0_\,
            carryout => \b2v_inst.eventos_cry_0\,
            clk => \N__22509\,
            ce => \N__8612\,
            sr => \N__22882\
        );

    \b2v_inst.eventos_1_LC_1_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9604\,
            in2 => \_gnd_net_\,
            in3 => \N__8564\,
            lcout => \b2v_inst.eventosZ0Z_1\,
            ltout => OPEN,
            carryin => \b2v_inst.eventos_cry_0\,
            carryout => \b2v_inst.eventos_cry_1\,
            clk => \N__22509\,
            ce => \N__8612\,
            sr => \N__22882\
        );

    \b2v_inst.eventos_2_LC_1_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8959\,
            in2 => \_gnd_net_\,
            in3 => \N__8561\,
            lcout => \b2v_inst.eventosZ0Z_2\,
            ltout => OPEN,
            carryin => \b2v_inst.eventos_cry_1\,
            carryout => \b2v_inst.eventos_cry_2\,
            clk => \N__22509\,
            ce => \N__8612\,
            sr => \N__22882\
        );

    \b2v_inst.eventos_3_LC_1_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8662\,
            in2 => \_gnd_net_\,
            in3 => \N__8558\,
            lcout => \b2v_inst.eventosZ0Z_3\,
            ltout => OPEN,
            carryin => \b2v_inst.eventos_cry_2\,
            carryout => \b2v_inst.eventos_cry_3\,
            clk => \N__22509\,
            ce => \N__8612\,
            sr => \N__22882\
        );

    \b2v_inst.eventos_4_LC_1_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8647\,
            in2 => \_gnd_net_\,
            in3 => \N__8555\,
            lcout => \b2v_inst.eventosZ0Z_4\,
            ltout => OPEN,
            carryin => \b2v_inst.eventos_cry_3\,
            carryout => \b2v_inst.eventos_cry_4\,
            clk => \N__22509\,
            ce => \N__8612\,
            sr => \N__22882\
        );

    \b2v_inst.eventos_5_LC_1_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8624\,
            in2 => \_gnd_net_\,
            in3 => \N__8552\,
            lcout => \b2v_inst.eventosZ0Z_5\,
            ltout => OPEN,
            carryin => \b2v_inst.eventos_cry_4\,
            carryout => \b2v_inst.eventos_cry_5\,
            clk => \N__22509\,
            ce => \N__8612\,
            sr => \N__22882\
        );

    \b2v_inst.eventos_6_LC_1_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9589\,
            in2 => \_gnd_net_\,
            in3 => \N__8549\,
            lcout => \b2v_inst.eventosZ0Z_6\,
            ltout => OPEN,
            carryin => \b2v_inst.eventos_cry_5\,
            carryout => \b2v_inst.eventos_cry_6\,
            clk => \N__22509\,
            ce => \N__8612\,
            sr => \N__22882\
        );

    \b2v_inst.eventos_7_LC_1_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9526\,
            in2 => \_gnd_net_\,
            in3 => \N__8546\,
            lcout => \b2v_inst.eventosZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22509\,
            ce => \N__8612\,
            sr => \N__22882\
        );

    \b2v_inst.data_a_escribir_RNO_1_7_LC_1_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000010011"
        )
    port map (
            in0 => \N__10695\,
            in1 => \N__10543\,
            in2 => \N__11222\,
            in3 => \N__10793\,
            lcout => \b2v_inst.un1_reg_anterior_iv_0_0_2_0_tz_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.reg_ancho_1_7_LC_1_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8885\,
            in2 => \_gnd_net_\,
            in3 => \N__13638\,
            lcout => \b2v_inst.reg_ancho_1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22570\,
            ce => \N__13913\,
            sr => \N__22886\
        );

    \b2v_inst.reg_ancho_1_6_LC_1_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__8884\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14241\,
            lcout => \b2v_inst.reg_ancho_1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22570\,
            ce => \N__13913\,
            sr => \N__22886\
        );

    \b2v_inst.data_a_escribir_RNO_4_3_LC_1_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000011011"
        )
    port map (
            in0 => \N__10542\,
            in1 => \N__11021\,
            in2 => \N__8663\,
            in3 => \N__10696\,
            lcout => \b2v_inst.un1_reg_anterior_iv_0_0_1_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_1_4_LC_1_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101010101"
        )
    port map (
            in0 => \N__14795\,
            in1 => \N__8648\,
            in2 => \_gnd_net_\,
            in3 => \N__10547\,
            lcout => \b2v_inst.un1_reg_anterior_iv_0_0_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_2_0_LC_1_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011111111"
        )
    port map (
            in0 => \N__10545\,
            in1 => \N__8636\,
            in2 => \_gnd_net_\,
            in3 => \N__14793\,
            lcout => \b2v_inst.un1_reg_anterior_iv_0_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_2_5_LC_1_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101010101"
        )
    port map (
            in0 => \N__14794\,
            in1 => \N__8623\,
            in2 => \_gnd_net_\,
            in3 => \N__10546\,
            lcout => \b2v_inst.un1_reg_anterior_iv_0_0_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNIN3GK_7_LC_1_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__10544\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14792\,
            lcout => \b2v_inst.N_47_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_un3_valor_max1_cry_0_c_inv_LC_1_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__10286\,
            in1 => \N__11511\,
            in2 => \N__8603\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst.reg_ancho_1_i_0\,
            ltout => OPEN,
            carryin => \bfn_1_17_0_\,
            carryout => \b2v_inst.un3_valor_max1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_un3_valor_max1_cry_1_c_inv_LC_1_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11473\,
            in2 => \N__8594\,
            in3 => \N__11155\,
            lcout => \b2v_inst.reg_ancho_1_i_1\,
            ltout => OPEN,
            carryin => \b2v_inst.un3_valor_max1_cry_0\,
            carryout => \b2v_inst.un3_valor_max1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_un3_valor_max1_cry_2_c_inv_LC_1_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11427\,
            in2 => \N__8585\,
            in3 => \N__11056\,
            lcout => \b2v_inst.reg_ancho_1_i_2\,
            ltout => OPEN,
            carryin => \b2v_inst.un3_valor_max1_cry_1\,
            carryout => \b2v_inst.un3_valor_max1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_un3_valor_max1_cry_3_c_inv_LC_1_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11386\,
            in2 => \N__8576\,
            in3 => \N__11011\,
            lcout => \b2v_inst.reg_ancho_1_i_3\,
            ltout => OPEN,
            carryin => \b2v_inst.un3_valor_max1_cry_2\,
            carryout => \b2v_inst.un3_valor_max1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_un3_valor_max1_cry_4_c_inv_LC_1_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11337\,
            in2 => \N__8702\,
            in3 => \N__10942\,
            lcout => \b2v_inst.reg_ancho_1_i_4\,
            ltout => OPEN,
            carryin => \b2v_inst.un3_valor_max1_cry_3\,
            carryout => \b2v_inst.un3_valor_max1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_un3_valor_max1_cry_5_c_inv_LC_1_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11304\,
            in2 => \N__8693\,
            in3 => \N__10870\,
            lcout => \b2v_inst.reg_ancho_1_i_5\,
            ltout => OPEN,
            carryin => \b2v_inst.un3_valor_max1_cry_4\,
            carryout => \b2v_inst.un3_valor_max1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_un3_valor_max1_cry_6_c_inv_LC_1_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11243\,
            in2 => \N__8684\,
            in3 => \N__10828\,
            lcout => \b2v_inst.reg_ancho_1_i_6\,
            ltout => OPEN,
            carryin => \b2v_inst.un3_valor_max1_cry_5\,
            carryout => \b2v_inst.un3_valor_max1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_un3_valor_max1_cry_7_c_inv_LC_1_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11213\,
            in2 => \N__8675\,
            in3 => \N__10783\,
            lcout => \b2v_inst.reg_ancho_1_i_7\,
            ltout => OPEN,
            carryin => \b2v_inst.un3_valor_max1_cry_6\,
            carryout => \b2v_inst.un3_valor_max1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un3_valor_max1_THRU_LUT4_0_LC_1_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8666\,
            lcout => \b2v_inst.un3_valor_max1_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_0_0_LC_1_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111010"
        )
    port map (
            in0 => \N__10287\,
            in1 => \N__11510\,
            in2 => \N__10570\,
            in3 => \N__10681\,
            lcout => \b2v_inst.un1_m3_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_4_2_LC_1_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11426\,
            in2 => \_gnd_net_\,
            in3 => \N__10680\,
            lcout => \b2v_inst.un1_reg_anterior_iv_0_0_a2_4_tz_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst3.reset_i_LC_1_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18933\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => reset_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final5_3_cry_0_c_LC_1_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9628\,
            in2 => \N__11513\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_19_0_\,
            carryout => \b2v_inst.valor_max_final5_3_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final5_3_cry_1_c_LC_1_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9871\,
            in2 => \N__11471\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.valor_max_final5_3_cry_0\,
            carryout => \b2v_inst.valor_max_final5_3_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final5_3_cry_2_c_LC_1_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9853\,
            in2 => \N__11429\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.valor_max_final5_3_cry_1\,
            carryout => \b2v_inst.valor_max_final5_3_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final5_3_cry_3_c_LC_1_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9835\,
            in2 => \N__11389\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.valor_max_final5_3_cry_2\,
            carryout => \b2v_inst.valor_max_final5_3_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final5_3_cry_4_c_LC_1_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11345\,
            in2 => \N__9818\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.valor_max_final5_3_cry_3\,
            carryout => \b2v_inst.valor_max_final5_3_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final5_3_cry_5_c_LC_1_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11308\,
            in2 => \N__9797\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.valor_max_final5_3_cry_4\,
            carryout => \b2v_inst.valor_max_final5_3_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final5_3_cry_6_c_LC_1_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11263\,
            in2 => \N__9775\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.valor_max_final5_3_cry_5\,
            carryout => \b2v_inst.valor_max_final5_3_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final5_3_cry_7_c_LC_1_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9752\,
            in2 => \N__11217\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.valor_max_final5_3_cry_6\,
            carryout => \b2v_inst.valor_max_final53\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.valor_max_final53_THRU_LUT4_0_LC_1_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8729\,
            lcout => \b2v_inst.valor_max_final53_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.ignorar_anterior_RNO_LC_1_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110001010000"
        )
    port map (
            in0 => \N__15683\,
            in1 => \N__8726\,
            in2 => \N__10172\,
            in3 => \N__8714\,
            lcout => \b2v_inst.un1_state_19_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un1_pix_count_anterior_0_I_1_c_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8750\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_11_0_\,
            carryout => \b2v_inst.un1_pix_count_anterior_0_data_tmp_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un1_pix_count_anterior_0_I_27_c_LC_2_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9101\,
            in2 => \N__18605\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.un1_pix_count_anterior_0_data_tmp_0\,
            carryout => \b2v_inst.un1_pix_count_anterior_0_data_tmp_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un1_pix_count_anterior_0_I_15_c_LC_2_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8735\,
            in2 => \N__18601\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.un1_pix_count_anterior_0_data_tmp_1\,
            carryout => \b2v_inst.un1_pix_count_anterior_0_data_tmp_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un1_pix_count_anterior_0_I_21_c_LC_2_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8792\,
            in2 => \N__18604\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.un1_pix_count_anterior_0_data_tmp_2\,
            carryout => \b2v_inst.un1_pix_count_anterior_0_data_tmp_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un1_pix_count_anterior_0_I_51_c_LC_2_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8837\,
            in2 => \N__18603\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.un1_pix_count_anterior_0_data_tmp_3\,
            carryout => \b2v_inst.un1_pix_count_anterior_0_data_tmp_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un1_pix_count_anterior_0_I_9_c_LC_2_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9080\,
            in2 => \N__18606\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.un1_pix_count_anterior_0_data_tmp_4\,
            carryout => \b2v_inst.un1_pix_count_anterior_0_data_tmp_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un1_pix_count_anterior_0_I_39_c_LC_2_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8801\,
            in2 => \N__18602\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.un1_pix_count_anterior_0_data_tmp_5\,
            carryout => \b2v_inst.un1_pix_count_anterior_0_N_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un1_pix_count_anterior_0_N_2_THRU_LUT4_0_LC_2_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8738\,
            lcout => \b2v_inst.un1_pix_count_anterior_0_N_2_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un1_pix_count_anterior_0_I_15_c_RNO_LC_2_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__9206\,
            in1 => \N__8774\,
            in2 => \N__8768\,
            in3 => \N__9185\,
            lcout => \b2v_inst.un1_pix_count_anterior_0_I_15_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.pix_count_anterior_4_LC_2_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9208\,
            lcout => \b2v_inst.pix_count_anteriorZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22587\,
            ce => \N__9338\,
            sr => \N__22877\
        );

    \b2v_inst.pix_count_anterior_5_LC_2_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9186\,
            lcout => \b2v_inst.pix_count_anteriorZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22587\,
            ce => \N__9338\,
            sr => \N__22877\
        );

    \b2v_inst4.pix_count_int_RNITN3K1_1_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__9158\,
            in1 => \N__9282\,
            in2 => \N__9263\,
            in3 => \N__9207\,
            lcout => \b2v_inst4.un1_pix_count_int_0_sqmuxa_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.pix_count_anterior_1_LC_2_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__9283\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst.pix_count_anteriorZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22587\,
            ce => \N__9338\,
            sr => \N__22877\
        );

    \b2v_inst.un1_pix_count_anterior_0_I_1_c_RNO_LC_2_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__8744\,
            in1 => \N__9308\,
            in2 => \N__8759\,
            in3 => \N__9281\,
            lcout => \b2v_inst.un1_pix_count_anterior_0_I_1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.pix_count_anterior_0_LC_2_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__9309\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst.pix_count_anteriorZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22587\,
            ce => \N__9338\,
            sr => \N__22877\
        );

    \b2v_inst.pix_count_anterior_2_LC_2_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__9262\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst.pix_count_anteriorZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22587\,
            ce => \N__9338\,
            sr => \N__22877\
        );

    \b2v_inst4.pix_count_int_0_LC_2_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__12007\,
            in1 => \N__11971\,
            in2 => \N__11944\,
            in3 => \N__9290\,
            lcout => \SYNTHESIZED_WIRE_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22496\,
            ce => 'H',
            sr => \N__22880\
        );

    \b2v_inst4.pix_count_int_11_LC_2_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__11972\,
            in1 => \N__12008\,
            in2 => \N__11923\,
            in3 => \N__9407\,
            lcout => \SYNTHESIZED_WIRE_2_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22496\,
            ce => 'H',
            sr => \N__22880\
        );

    \b2v_inst4.pix_count_int_12_LC_2_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__12009\,
            in1 => \N__11973\,
            in2 => \N__11945\,
            in3 => \N__9368\,
            lcout => \SYNTHESIZED_WIRE_2_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22496\,
            ce => 'H',
            sr => \N__22880\
        );

    \b2v_inst.un1_pix_count_anterior_0_I_39_c_RNO_LC_2_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8807\,
            in2 => \_gnd_net_\,
            in3 => \N__9392\,
            lcout => \b2v_inst.un1_pix_count_anterior_0_I_39_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst4.pix_count_int_3_LC_2_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__12010\,
            in1 => \N__11974\,
            in2 => \N__11946\,
            in3 => \N__9218\,
            lcout => \SYNTHESIZED_WIRE_2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22496\,
            ce => 'H',
            sr => \N__22880\
        );

    \b2v_inst4.pix_count_int_5_LC_2_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__11975\,
            in1 => \N__12011\,
            in2 => \N__11924\,
            in3 => \N__9167\,
            lcout => \SYNTHESIZED_WIRE_2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22496\,
            ce => 'H',
            sr => \N__22880\
        );

    \b2v_inst4.pix_count_int_7_LC_2_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__12012\,
            in1 => \N__11976\,
            in2 => \N__11947\,
            in3 => \N__9494\,
            lcout => \SYNTHESIZED_WIRE_2_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22496\,
            ce => 'H',
            sr => \N__22880\
        );

    \b2v_inst4.pix_count_int_8_LC_2_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__11977\,
            in1 => \N__12013\,
            in2 => \N__11925\,
            in3 => \N__9467\,
            lcout => \SYNTHESIZED_WIRE_2_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22496\,
            ce => 'H',
            sr => \N__22880\
        );

    \b2v_inst.un1_pix_count_anterior_0_I_21_c_RNO_LC_2_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__9509\,
            in1 => \N__8783\,
            in2 => \N__8852\,
            in3 => \N__9155\,
            lcout => \b2v_inst.un1_pix_count_anterior_0_I_21_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.pix_count_anterior_6_LC_2_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__9156\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst.pix_count_anteriorZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22588\,
            ce => \N__9341\,
            sr => \N__22883\
        );

    \b2v_inst4.pix_count_int_RNI6KOL1_12_LC_2_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9428\,
            in1 => \N__11868\,
            in2 => \N__9398\,
            in3 => \N__9483\,
            lcout => OPEN,
            ltout => \b2v_inst4.un1_pix_count_int_0_sqmuxa_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst4.state_RNIC9UM2_0_LC_2_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__11714\,
            in1 => \N__9510\,
            in2 => \N__8777\,
            in3 => \N__9188\,
            lcout => \b2v_inst4.un1_pix_count_int_0_sqmuxa_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.pix_count_anterior_7_LC_2_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__9511\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst.pix_count_anteriorZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22588\,
            ce => \N__9341\,
            sr => \N__22883\
        );

    \b2v_inst.pix_count_anterior_8_LC_2_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__9484\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst.pix_count_anteriorZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22588\,
            ce => \N__9341\,
            sr => \N__22883\
        );

    \b2v_inst.un1_pix_count_anterior_0_I_51_c_RNO_LC_2_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__8843\,
            in1 => \N__11867\,
            in2 => \N__8828\,
            in3 => \N__9482\,
            lcout => \b2v_inst.un1_pix_count_anterior_0_I_51_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.pix_count_anterior_9_LC_2_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__11869\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst.pix_count_anteriorZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22588\,
            ce => \N__9341\,
            sr => \N__22883\
        );

    \b2v_inst.ignorar_ancho_1_LC_2_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15678\,
            lcout => \b2v_inst.ignorar_anchoZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22578\,
            ce => \N__8819\,
            sr => \N__22887\
        );

    \b2v_inst.data_a_escribir9_0_c_RNO_LC_2_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__11060\,
            in1 => \N__11156\,
            in2 => \N__11022\,
            in3 => \N__10282\,
            lcout => \b2v_inst.data_a_escribir9_0_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.reg_ancho_1_0_LC_2_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__13095\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8878\,
            lcout => \b2v_inst.reg_ancho_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22606\,
            ce => \N__13912\,
            sr => \N__22892\
        );

    \b2v_inst.reg_ancho_1_1_LC_2_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__8879\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13020\,
            lcout => \b2v_inst.reg_ancho_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22606\,
            ce => \N__13912\,
            sr => \N__22892\
        );

    \b2v_inst.reg_ancho_1_2_LC_2_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8880\,
            in2 => \_gnd_net_\,
            in3 => \N__12951\,
            lcout => \b2v_inst.reg_ancho_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22606\,
            ce => \N__13912\,
            sr => \N__22892\
        );

    \b2v_inst.reg_ancho_1_3_LC_2_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__8881\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12879\,
            lcout => \b2v_inst.reg_ancho_1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22606\,
            ce => \N__13912\,
            sr => \N__22892\
        );

    \b2v_inst.reg_ancho_1_4_LC_2_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__13545\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8882\,
            lcout => \b2v_inst.reg_ancho_1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22606\,
            ce => \N__13912\,
            sr => \N__22892\
        );

    \b2v_inst.data_a_escribir9_1_c_RNO_LC_2_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__10829\,
            in1 => \N__10871\,
            in2 => \N__10794\,
            in3 => \N__10946\,
            lcout => \b2v_inst.data_a_escribir9_1_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.reg_ancho_1_5_LC_2_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14693\,
            in2 => \_gnd_net_\,
            in3 => \N__8883\,
            lcout => \b2v_inst.reg_ancho_1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22606\,
            ce => \N__13912\,
            sr => \N__22892\
        );

    \b2v_inst.data_a_escribir9_3_c_RNO_LC_2_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__11242\,
            in1 => \N__11293\,
            in2 => \N__11203\,
            in3 => \N__11326\,
            lcout => \b2v_inst.data_a_escribir9_3_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.reg_ancho_2_4_LC_2_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13553\,
            lcout => \b2v_inst.reg_ancho_2Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22564\,
            ce => \N__15490\,
            sr => \N__22897\
        );

    \b2v_inst.reg_ancho_2_5_LC_2_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14704\,
            lcout => \b2v_inst.reg_ancho_2Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22564\,
            ce => \N__15490\,
            sr => \N__22897\
        );

    \b2v_inst.reg_ancho_2_6_LC_2_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14243\,
            lcout => \b2v_inst.reg_ancho_2Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22564\,
            ce => \N__15490\,
            sr => \N__22897\
        );

    \b2v_inst.reg_ancho_2_7_LC_2_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13642\,
            lcout => \b2v_inst.reg_ancho_2Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22564\,
            ce => \N__15490\,
            sr => \N__22897\
        );

    \b2v_inst.data_a_escribir_RNO_3_4_LC_2_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__11327\,
            in1 => \N__10516\,
            in2 => \_gnd_net_\,
            in3 => \N__10679\,
            lcout => OPEN,
            ltout => \b2v_inst.data_a_escribir_RNO_3Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_0_4_LC_2_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9668\,
            in2 => \N__8933\,
            in3 => \N__10950\,
            lcout => \b2v_inst.data_a_escribir_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_un3_valor_max1_cry_7_c_RNIV45S_LC_2_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10515\,
            in2 => \_gnd_net_\,
            in3 => \N__10678\,
            lcout => \b2v_inst.un1_reg_anterior_iv_0_0_a2_4_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_3_0_LC_2_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__10250\,
            in1 => \N__10557\,
            in2 => \_gnd_net_\,
            in3 => \N__13219\,
            lcout => OPEN,
            ltout => \b2v_inst.data_a_escribir_RNO_3Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_1_0_LC_2_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10611\,
            in2 => \N__8930\,
            in3 => \N__13067\,
            lcout => OPEN,
            ltout => \b2v_inst.data_a_escribir_RNO_1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_0_LC_2_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001010000"
        )
    port map (
            in0 => \N__8927\,
            in1 => \N__8915\,
            in2 => \N__8909\,
            in3 => \N__10431\,
            lcout => b2v_inst_data_a_escribir_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22607\,
            ce => \N__10350\,
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_3_3_LC_2_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100011111111"
        )
    port map (
            in0 => \N__8906\,
            in1 => \N__10426\,
            in2 => \N__10569\,
            in3 => \N__14797\,
            lcout => \b2v_inst.un1_reg_anterior_iv_0_0_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_0_3_LC_2_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__10706\,
            in1 => \N__10558\,
            in2 => \N__11390\,
            in3 => \N__10430\,
            lcout => OPEN,
            ltout => \b2v_inst.N_315_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_3_LC_2_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__8978\,
            in1 => \N__8942\,
            in2 => \N__8897\,
            in3 => \N__8894\,
            lcout => b2v_inst_data_a_escribir_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22607\,
            ce => \N__10350\,
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_un3_valor_max2_cry_7_c_RNI0D1L_LC_2_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10553\,
            in2 => \_gnd_net_\,
            in3 => \N__13218\,
            lcout => \b2v_inst.un1_reg_anterior_iv_0_0_a2_6_0_1\,
            ltout => \b2v_inst.un1_reg_anterior_iv_0_0_a2_6_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_1_3_LC_2_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10425\,
            in2 => \N__8888\,
            in3 => \N__12851\,
            lcout => \b2v_inst.N_317\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir9_2_c_RNO_LC_2_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__11419\,
            in1 => \N__11458\,
            in2 => \N__11387\,
            in3 => \N__11506\,
            lcout => \b2v_inst.data_a_escribir9_2_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.reg_ancho_2_0_LC_2_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13103\,
            lcout => \b2v_inst.reg_ancho_2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22597\,
            ce => \N__15491\,
            sr => \N__22907\
        );

    \b2v_inst.reg_ancho_2_1_LC_2_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13031\,
            lcout => \b2v_inst.reg_ancho_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22597\,
            ce => \N__15491\,
            sr => \N__22907\
        );

    \b2v_inst.reg_ancho_2_2_LC_2_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12959\,
            lcout => \b2v_inst.reg_ancho_2Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22597\,
            ce => \N__15491\,
            sr => \N__22907\
        );

    \b2v_inst.reg_ancho_2_3_LC_2_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12887\,
            lcout => \b2v_inst.reg_ancho_2Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22597\,
            ce => \N__15491\,
            sr => \N__22907\
        );

    \b2v_inst.data_a_escribir_RNO_2_2_LC_2_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000000000"
        )
    port map (
            in0 => \N__11635\,
            in1 => \N__9727\,
            in2 => \N__13238\,
            in3 => \N__8972\,
            lcout => OPEN,
            ltout => \b2v_inst.N_320_tz_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_0_2_LC_2_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111110011"
        )
    port map (
            in0 => \N__8966\,
            in1 => \N__14798\,
            in2 => \N__8948\,
            in3 => \N__10563\,
            lcout => \b2v_inst.un1_reg_anterior_iv_0_0_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final5_0_cry_7_c_RNI5KAH1_LC_2_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100011011"
        )
    port map (
            in0 => \N__10688\,
            in1 => \N__10727\,
            in2 => \N__11636\,
            in3 => \N__13227\,
            lcout => \b2v_inst.un1_m3_0_m3_ns_1\,
            ltout => \b2v_inst.un1_m3_0_m3_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_2_3_LC_2_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__13228\,
            in1 => \N__10562\,
            in2 => \N__8945\,
            in3 => \N__10988\,
            lcout => \b2v_inst.N_318\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_4_LC_2_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000000101"
        )
    port map (
            in0 => \N__9899\,
            in1 => \N__9074\,
            in2 => \N__9065\,
            in3 => \N__10419\,
            lcout => b2v_inst_data_a_escribir_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22596\,
            ce => \N__10349\,
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNIA6JL_4_LC_2_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__17717\,
            in1 => \N__17033\,
            in2 => \_gnd_net_\,
            in3 => \N__14509\,
            lcout => \N_211_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNI62JL_0_LC_2_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010100000"
        )
    port map (
            in0 => \N__17031\,
            in1 => \_gnd_net_\,
            in2 => \N__13459\,
            in3 => \N__17716\,
            lcout => \N_219_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNI73JL_1_LC_2_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17032\,
            in2 => \N__13480\,
            in3 => \N__17714\,
            lcout => \N_217_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNI84JL_2_LC_2_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__17030\,
            in1 => \N__13411\,
            in2 => \_gnd_net_\,
            in3 => \N__17715\,
            lcout => \N_215_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_11_LC_3_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010101000000000"
        )
    port map (
            in0 => \N__15682\,
            in1 => \N__9125\,
            in2 => \N__8993\,
            in3 => \N__10208\,
            lcout => \b2v_inst.stateZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22481\,
            ce => 'H',
            sr => \N__22878\
        );

    \b2v_inst.state_ns_i_i_a2_4_6_LC_3_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__10070\,
            in1 => \N__10082\,
            in2 => \N__10058\,
            in3 => \N__10094\,
            lcout => \b2v_inst.state_ns_i_i_a2_4Z0Z_6\,
            ltout => \b2v_inst.state_ns_i_i_a2_4Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un1_pix_count_anterior_0_I_39_c_RNIP5QR3_LC_3_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__15681\,
            in1 => \N__9124\,
            in2 => \N__8984\,
            in3 => \N__10207\,
            lcout => \b2v_inst.N_497\,
            ltout => \b2v_inst.N_497_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_6_LC_3_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__9134\,
            in1 => \N__14791\,
            in2 => \N__8981\,
            in3 => \N__14873\,
            lcout => \b2v_inst.stateZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22481\,
            ce => 'H',
            sr => \N__22878\
        );

    \b2v_inst.state_RNO_0_6_LC_3_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17702\,
            in2 => \_gnd_net_\,
            in3 => \N__15680\,
            lcout => \b2v_inst.N_361\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_ns_i_i_a2_5_6_LC_3_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__9911\,
            in1 => \N__9923\,
            in2 => \N__10043\,
            in3 => \N__9935\,
            lcout => \b2v_inst.state_ns_i_i_a2_5Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un1_pix_count_anterior_0_I_39_c_RNIT6R7_LC_3_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15679\,
            in2 => \_gnd_net_\,
            in3 => \N__10206\,
            lcout => \b2v_inst.N_254_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.borrado_LC_3_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__17703\,
            in1 => \N__15901\,
            in2 => \_gnd_net_\,
            in3 => \N__18776\,
            lcout => \b2v_inst.borradoZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22481\,
            ce => 'H',
            sr => \N__22878\
        );

    \b2v_inst.un1_pix_count_anterior_0_I_27_c_RNO_LC_3_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__9107\,
            in1 => \N__9233\,
            in2 => \N__9095\,
            in3 => \N__9257\,
            lcout => \b2v_inst.un1_pix_count_anterior_0_I_27_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.pix_count_anterior_3_LC_3_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__9235\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst.pix_count_anteriorZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22380\,
            ce => \N__9340\,
            sr => \N__22881\
        );

    \b2v_inst4.pix_count_int_RNIATHH1_0_LC_3_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__9454\,
            in1 => \N__9234\,
            in2 => \N__9317\,
            in3 => \N__15721\,
            lcout => \b2v_inst4.un1_pix_count_int_0_sqmuxa_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.pix_count_anterior_10_LC_3_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9455\,
            lcout => \b2v_inst.pix_count_anteriorZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22380\,
            ce => \N__9340\,
            sr => \N__22881\
        );

    \b2v_inst.un1_pix_count_anterior_0_I_9_c_RNO_LC_3_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__9086\,
            in1 => \N__9425\,
            in2 => \N__9350\,
            in3 => \N__9453\,
            lcout => \b2v_inst.un1_pix_count_anterior_0_I_9_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.pix_count_anterior_11_LC_3_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__9426\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst.pix_count_anteriorZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22380\,
            ce => \N__9340\,
            sr => \N__22881\
        );

    \b2v_inst4.state_RNICJOG_0_LC_3_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11713\,
            in2 => \_gnd_net_\,
            in3 => \N__15720\,
            lcout => \b2v_inst4.pix_count_int_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst4.pix_count_int_RNO_0_0_LC_3_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9310\,
            in2 => \N__10027\,
            in3 => \N__10023\,
            lcout => \b2v_inst4.pix_count_int_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \bfn_3_13_0_\,
            carryout => \b2v_inst4.un1_pix_count_int_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst4.pix_count_int_1_LC_3_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9284\,
            in2 => \_gnd_net_\,
            in3 => \N__9266\,
            lcout => \SYNTHESIZED_WIRE_2_1\,
            ltout => OPEN,
            carryin => \b2v_inst4.un1_pix_count_int_cry_0\,
            carryout => \b2v_inst4.un1_pix_count_int_cry_1\,
            clk => \N__22482\,
            ce => 'H',
            sr => \N__22884\
        );

    \b2v_inst4.pix_count_int_2_LC_3_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9258\,
            in2 => \_gnd_net_\,
            in3 => \N__9239\,
            lcout => \SYNTHESIZED_WIRE_2_2\,
            ltout => OPEN,
            carryin => \b2v_inst4.un1_pix_count_int_cry_1\,
            carryout => \b2v_inst4.un1_pix_count_int_cry_2\,
            clk => \N__22482\,
            ce => 'H',
            sr => \N__22884\
        );

    \b2v_inst4.pix_count_int_RNO_0_3_LC_3_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9236\,
            in2 => \_gnd_net_\,
            in3 => \N__9212\,
            lcout => \b2v_inst4.pix_count_int_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \b2v_inst4.un1_pix_count_int_cry_2\,
            carryout => \b2v_inst4.un1_pix_count_int_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst4.pix_count_int_4_LC_3_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9209\,
            in2 => \_gnd_net_\,
            in3 => \N__9191\,
            lcout => \SYNTHESIZED_WIRE_2_4\,
            ltout => OPEN,
            carryin => \b2v_inst4.un1_pix_count_int_cry_3\,
            carryout => \b2v_inst4.un1_pix_count_int_cry_4\,
            clk => \N__22482\,
            ce => 'H',
            sr => \N__22884\
        );

    \b2v_inst4.pix_count_int_RNO_0_5_LC_3_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9187\,
            in2 => \_gnd_net_\,
            in3 => \N__9161\,
            lcout => \b2v_inst4.pix_count_int_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \b2v_inst4.un1_pix_count_int_cry_4\,
            carryout => \b2v_inst4.un1_pix_count_int_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst4.pix_count_int_6_LC_3_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9157\,
            in2 => \_gnd_net_\,
            in3 => \N__9137\,
            lcout => \SYNTHESIZED_WIRE_2_6\,
            ltout => OPEN,
            carryin => \b2v_inst4.un1_pix_count_int_cry_5\,
            carryout => \b2v_inst4.un1_pix_count_int_cry_6\,
            clk => \N__22482\,
            ce => 'H',
            sr => \N__22884\
        );

    \b2v_inst4.pix_count_int_RNO_0_7_LC_3_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9512\,
            in2 => \_gnd_net_\,
            in3 => \N__9488\,
            lcout => \b2v_inst4.pix_count_int_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \b2v_inst4.un1_pix_count_int_cry_6\,
            carryout => \b2v_inst4.un1_pix_count_int_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst4.pix_count_int_RNO_0_8_LC_3_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9485\,
            in2 => \_gnd_net_\,
            in3 => \N__9461\,
            lcout => \b2v_inst4.pix_count_int_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \bfn_3_14_0_\,
            carryout => \b2v_inst4.un1_pix_count_int_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst4.pix_count_int_RNO_0_9_LC_3_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11870\,
            in2 => \_gnd_net_\,
            in3 => \N__9458\,
            lcout => \b2v_inst4.pix_count_int_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \b2v_inst4.un1_pix_count_int_cry_8\,
            carryout => \b2v_inst4.un1_pix_count_int_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst4.pix_count_int_10_LC_3_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9452\,
            in2 => \_gnd_net_\,
            in3 => \N__9431\,
            lcout => \SYNTHESIZED_WIRE_2_10\,
            ltout => OPEN,
            carryin => \b2v_inst4.un1_pix_count_int_cry_9\,
            carryout => \b2v_inst4.un1_pix_count_int_cry_10\,
            clk => \N__22381\,
            ce => 'H',
            sr => \N__22888\
        );

    \b2v_inst4.pix_count_int_RNO_0_11_LC_3_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9427\,
            in2 => \_gnd_net_\,
            in3 => \N__9401\,
            lcout => \b2v_inst4.pix_count_int_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \b2v_inst4.un1_pix_count_int_cry_10\,
            carryout => \b2v_inst4.un1_pix_count_int_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst4.pix_count_int_RNO_0_12_LC_3_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9396\,
            in2 => \_gnd_net_\,
            in3 => \N__9371\,
            lcout => \b2v_inst4.pix_count_int_RNO_0Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir9_0_c_LC_3_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9362\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_3_15_0_\,
            carryout => \b2v_inst.data_a_escribir9_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir9_1_c_LC_3_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9356\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.data_a_escribir9_0\,
            carryout => \b2v_inst.data_a_escribir9_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir9_2_c_LC_3_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9554\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.data_a_escribir9_1\,
            carryout => \b2v_inst.data_a_escribir9_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir9_3_c_LC_3_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9542\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.data_a_escribir9_2\,
            carryout => \b2v_inst.data_a_escribir9_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir9_4_c_LC_3_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10106\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.data_a_escribir9_3\,
            carryout => \b2v_inst.data_a_escribir9_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir9_5_c_LC_3_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10715\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.data_a_escribir9_4\,
            carryout => \b2v_inst.data_a_escribir9_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir9_6_c_LC_3_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11525\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.data_a_escribir9_5\,
            carryout => \b2v_inst.data_a_escribir9_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir9_7_c_LC_3_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13568\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.data_a_escribir9_6\,
            carryout => \b2v_inst.data_a_escribir10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir10_THRU_LUT4_0_LC_3_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9533\,
            lcout => \b2v_inst.data_a_escribir10_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_RX_Byte_0_LC_3_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__17126\,
            in1 => \N__9946\,
            in2 => \N__22751\,
            in3 => \N__17177\,
            lcout => \SYNTHESIZED_WIRE_10_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22605\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_0_7_LC_3_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011111111"
        )
    port map (
            in0 => \N__10511\,
            in1 => \N__9530\,
            in2 => \_gnd_net_\,
            in3 => \N__14785\,
            lcout => \b2v_inst.un1_reg_anterior_iv_0_0_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_2_1_LC_3_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101010101"
        )
    port map (
            in0 => \N__14787\,
            in1 => \N__9611\,
            in2 => \_gnd_net_\,
            in3 => \N__10514\,
            lcout => \b2v_inst.un1_reg_anterior_iv_0_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_3_2_LC_3_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100010001"
        )
    port map (
            in0 => \N__10513\,
            in1 => \N__11102\,
            in2 => \N__12923\,
            in3 => \N__13232\,
            lcout => \b2v_inst.un1_reg_anterior_iv_0_0_2_tz_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_3_6_LC_3_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__13231\,
            in1 => \N__10510\,
            in2 => \_gnd_net_\,
            in3 => \N__12812\,
            lcout => \b2v_inst.data_a_escribir_RNO_3Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_2_6_LC_3_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011111111"
        )
    port map (
            in0 => \N__10512\,
            in1 => \N__9593\,
            in2 => \_gnd_net_\,
            in3 => \N__14786\,
            lcout => \b2v_inst.un1_reg_anterior_iv_0_0_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_3_1_LC_3_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__11472\,
            in1 => \N__10517\,
            in2 => \_gnd_net_\,
            in3 => \N__10705\,
            lcout => OPEN,
            ltout => \b2v_inst.un1_reg_anterior_iv_0_0_2_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_0_1_LC_3_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9669\,
            in2 => \N__9575\,
            in3 => \N__11163\,
            lcout => \b2v_inst.data_a_escribir_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_4_1_LC_3_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__11129\,
            in1 => \N__10518\,
            in2 => \_gnd_net_\,
            in3 => \N__13237\,
            lcout => OPEN,
            ltout => \b2v_inst.data_a_escribir_RNO_4Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_1_1_LC_3_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12992\,
            in2 => \N__9572\,
            in3 => \N__10612\,
            lcout => OPEN,
            ltout => \b2v_inst.data_a_escribir_RNO_1Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_1_LC_3_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001010000"
        )
    port map (
            in0 => \N__9569\,
            in1 => \N__9563\,
            in2 => \N__9557\,
            in3 => \N__10429\,
            lcout => b2v_inst_data_a_escribir_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22563\,
            ce => \N__10352\,
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNI9HNM5_7_LC_3_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010110000"
        )
    port map (
            in0 => \N__14781\,
            in1 => \N__14872\,
            in2 => \N__18941\,
            in3 => \N__9704\,
            lcout => \b2v_inst.un1_reset_inv_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_1_2_LC_3_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001101010101"
        )
    port map (
            in0 => \N__9695\,
            in1 => \N__9670\,
            in2 => \N__11075\,
            in3 => \N__10427\,
            lcout => OPEN,
            ltout => \b2v_inst.data_a_escribir_RNO_1Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_2_LC_3_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9686\,
            in3 => \N__9683\,
            lcout => b2v_inst_data_a_escribir_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22565\,
            ce => \N__10333\,
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_4_5_LC_3_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__10540\,
            in1 => \N__12791\,
            in2 => \_gnd_net_\,
            in3 => \N__13223\,
            lcout => OPEN,
            ltout => \b2v_inst.data_a_escribir_RNO_4Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_1_5_LC_3_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14663\,
            in2 => \N__9677\,
            in3 => \N__10610\,
            lcout => \b2v_inst.data_a_escribir_RNO_1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_3_5_LC_3_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__10541\,
            in1 => \N__11303\,
            in2 => \_gnd_net_\,
            in3 => \N__10700\,
            lcout => OPEN,
            ltout => \b2v_inst.un1_reg_anterior_iv_0_0_2_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_0_5_LC_3_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10885\,
            in2 => \N__9674\,
            in3 => \N__9671\,
            lcout => OPEN,
            ltout => \b2v_inst.data_a_escribir_RNO_0Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_5_LC_3_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__10428\,
            in1 => \N__9650\,
            in2 => \N__9638\,
            in3 => \N__9635\,
            lcout => b2v_inst_data_a_escribir_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22565\,
            ce => \N__10333\,
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final5_1_cry_0_c_inv_LC_3_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10295\,
            in2 => \N__9629\,
            in3 => \N__13059\,
            lcout => \b2v_inst.reg_anterior_i_0\,
            ltout => OPEN,
            carryin => \bfn_3_19_0_\,
            carryout => \b2v_inst.valor_max_final5_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final5_1_cry_1_c_inv_LC_3_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11167\,
            in2 => \N__9872\,
            in3 => \N__12987\,
            lcout => \b2v_inst.reg_anterior_i_1\,
            ltout => OPEN,
            carryin => \b2v_inst.valor_max_final5_1_cry_0\,
            carryout => \b2v_inst.valor_max_final5_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final5_1_cry_2_c_inv_LC_3_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11070\,
            in2 => \N__9854\,
            in3 => \N__12915\,
            lcout => \b2v_inst.reg_anterior_i_2\,
            ltout => OPEN,
            carryin => \b2v_inst.valor_max_final5_1_cry_1\,
            carryout => \b2v_inst.valor_max_final5_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final5_1_cry_3_c_inv_LC_3_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11032\,
            in2 => \N__9836\,
            in3 => \N__12845\,
            lcout => \b2v_inst.reg_anterior_i_3\,
            ltout => OPEN,
            carryin => \b2v_inst.valor_max_final5_1_cry_2\,
            carryout => \b2v_inst.valor_max_final5_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final5_1_cry_4_c_inv_LC_3_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__13509\,
            in1 => \N__10954\,
            in2 => \N__9817\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst.reg_anterior_i_4\,
            ltout => OPEN,
            carryin => \b2v_inst.valor_max_final5_1_cry_3\,
            carryout => \b2v_inst.valor_max_final5_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final5_1_cry_5_c_inv_LC_3_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10884\,
            in2 => \N__9796\,
            in3 => \N__14658\,
            lcout => \b2v_inst.reg_anterior_i_5\,
            ltout => OPEN,
            carryin => \b2v_inst.valor_max_final5_1_cry_4\,
            carryout => \b2v_inst.valor_max_final5_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final5_1_cry_6_c_inv_LC_3_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10847\,
            in2 => \N__9776\,
            in3 => \N__14199\,
            lcout => \b2v_inst.reg_anterior_i_6\,
            ltout => OPEN,
            carryin => \b2v_inst.valor_max_final5_1_cry_5\,
            carryout => \b2v_inst.valor_max_final5_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final5_1_cry_7_c_inv_LC_3_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10802\,
            in2 => \N__9751\,
            in3 => \N__13604\,
            lcout => \b2v_inst.reg_anterior_i_7\,
            ltout => OPEN,
            carryin => \b2v_inst.valor_max_final5_1_cry_6\,
            carryout => \b2v_inst.valor_max_final51\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final5_1_cry_7_c_RNIVOP62_LC_3_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__13229\,
            in1 => \N__9731\,
            in2 => \N__9716\,
            in3 => \N__9707\,
            lcout => \b2v_inst.N_264\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_2_4_LC_3_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000111"
        )
    port map (
            in0 => \N__13230\,
            in1 => \N__13514\,
            in2 => \N__10571\,
            in3 => \N__10916\,
            lcout => \b2v_inst.un1_reg_anterior_iv_0_0_2_tz_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst3.fsm_state_RNO_2_0_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__12157\,
            in1 => \N__12234\,
            in2 => \_gnd_net_\,
            in3 => \N__11600\,
            lcout => \b2v_inst3.N_434\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst3.fsm_state_RNO_0_1_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__12235\,
            in1 => \N__12158\,
            in2 => \_gnd_net_\,
            in3 => \N__11536\,
            lcout => OPEN,
            ltout => \b2v_inst3.fsm_state_ns_0_0_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst3.fsm_state_1_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000001000"
        )
    port map (
            in0 => \N__12159\,
            in1 => \N__18863\,
            in2 => \N__9893\,
            in3 => \N__13357\,
            lcout => \b2v_inst3.fsm_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22447\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst3.fsm_state_RNO_0_0_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001010"
        )
    port map (
            in0 => \N__12233\,
            in1 => \_gnd_net_\,
            in2 => \N__12166\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst3.N_490\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst3.fsm_state_RNIDA67_0_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12153\,
            in2 => \_gnd_net_\,
            in3 => \N__12232\,
            lcout => \N_230\,
            ltout => \N_230_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst3.fsm_state_RNO_1_0_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001101"
        )
    port map (
            in0 => \N__12265\,
            in1 => \N__11537\,
            in2 => \N__9890\,
            in3 => \N__9887\,
            lcout => OPEN,
            ltout => \b2v_inst3.fsm_state_ns_i_i_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst3.fsm_state_0_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001000001010"
        )
    port map (
            in0 => \N__18915\,
            in1 => \N__9881\,
            in2 => \N__9875\,
            in3 => \N__13351\,
            lcout => \b2v_inst3.fsm_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22267\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNIAJF6_9_LC_5_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__18914\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13970\,
            lcout => \b2v_inst.N_138_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst3.cycle_counter_6_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010001000100"
        )
    port map (
            in0 => \N__13349\,
            in1 => \N__11690\,
            in2 => \N__9970\,
            in3 => \N__11672\,
            lcout => \b2v_inst3.cycle_counterZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22515\,
            ce => 'H',
            sr => \N__22889\
        );

    \b2v_inst3.cycle_counter_7_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__11653\,
            in1 => \N__11689\,
            in2 => \N__9971\,
            in3 => \N__11670\,
            lcout => \b2v_inst3.cycle_counterZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22515\,
            ce => 'H',
            sr => \N__22889\
        );

    \b2v_inst3.cycle_counter_RNI4OAT_4_LC_5_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__12058\,
            in1 => \N__12035\,
            in2 => \_gnd_net_\,
            in3 => \N__12118\,
            lcout => OPEN,
            ltout => \b2v_inst3.un1_m2_0_a2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst3.cycle_counter_RNIIR2O1_1_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__14298\,
            in1 => \N__12081\,
            in2 => \N__9974\,
            in3 => \N__12198\,
            lcout => \b2v_inst3.un1_cycle_counter_5_c5\,
            ltout => \b2v_inst3.un1_cycle_counter_5_c5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst3.cycle_counter_5_LC_5_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001011010"
        )
    port map (
            in0 => \N__11671\,
            in1 => \_gnd_net_\,
            in2 => \N__9956\,
            in3 => \N__13348\,
            lcout => \b2v_inst3.cycle_counterZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22515\,
            ce => 'H',
            sr => \N__22889\
        );

    \b2v_inst3.cycle_counter_3_LC_5_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001101010"
        )
    port map (
            in0 => \N__12059\,
            in1 => \N__12095\,
            in2 => \N__12089\,
            in3 => \N__13347\,
            lcout => \b2v_inst3.cycle_counterZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22515\,
            ce => 'H',
            sr => \N__22889\
        );

    \b2v_inst3.cycle_counter_2_LC_5_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__12199\,
            in1 => \N__14299\,
            in2 => \N__12088\,
            in3 => \N__12119\,
            lcout => \b2v_inst3.cycle_counterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22515\,
            ce => 'H',
            sr => \N__22889\
        );

    \b2v_inst4.reg_data_0_LC_5_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9953\,
            lcout => \SYNTHESIZED_WIRE_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22405\,
            ce => \N__10028\,
            sr => \N__22893\
        );

    \b2v_inst4.reg_data_1_LC_5_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15749\,
            lcout => \SYNTHESIZED_WIRE_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22405\,
            ce => \N__10028\,
            sr => \N__22893\
        );

    \b2v_inst4.reg_data_2_LC_5_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12350\,
            lcout => \SYNTHESIZED_WIRE_3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22405\,
            ce => \N__10028\,
            sr => \N__22893\
        );

    \b2v_inst4.reg_data_3_LC_5_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12338\,
            lcout => \SYNTHESIZED_WIRE_3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22405\,
            ce => \N__10028\,
            sr => \N__22893\
        );

    \b2v_inst4.reg_data_4_LC_5_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12326\,
            lcout => \SYNTHESIZED_WIRE_3_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22405\,
            ce => \N__10028\,
            sr => \N__22893\
        );

    \b2v_inst4.reg_data_5_LC_5_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12314\,
            lcout => \SYNTHESIZED_WIRE_3_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22405\,
            ce => \N__10028\,
            sr => \N__22893\
        );

    \b2v_inst4.reg_data_6_LC_5_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12301\,
            lcout => \SYNTHESIZED_WIRE_3_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22405\,
            ce => \N__10028\,
            sr => \N__22893\
        );

    \b2v_inst4.reg_data_7_LC_5_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12557\,
            lcout => \SYNTHESIZED_WIRE_3_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22405\,
            ce => \N__10028\,
            sr => \N__22893\
        );

    \b2v_inst.state_RNINUTP_2_LC_5_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__10143\,
            in1 => \N__16481\,
            in2 => \N__14796\,
            in3 => \N__15234\,
            lcout => OPEN,
            ltout => \b2v_inst.we_0_a2_0_a2_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNIJHF42_2_LC_5_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__9980\,
            in1 => \N__16958\,
            in2 => \N__9995\,
            in3 => \N__15380\,
            lcout => \SYNTHESIZED_WIRE_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNICN8L_3_LC_5_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__10182\,
            in1 => \N__15632\,
            in2 => \N__12278\,
            in3 => \N__18998\,
            lcout => \b2v_inst.we_0_a2_0_a2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNI3LTB_3_LC_5_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12276\,
            in2 => \_gnd_net_\,
            in3 => \N__10183\,
            lcout => \N_458\,
            ltout => \N_458_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_3_LC_5_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111100001010"
        )
    port map (
            in0 => \N__12277\,
            in1 => \_gnd_net_\,
            in2 => \N__10223\,
            in3 => \N__14322\,
            lcout => \b2v_inst.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22517\,
            ce => 'H',
            sr => \N__22898\
        );

    \b2v_inst.state_RNO_0_16_LC_5_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000101"
        )
    port map (
            in0 => \N__15633\,
            in1 => \N__17698\,
            in2 => \N__10157\,
            in3 => \N__18774\,
            lcout => OPEN,
            ltout => \b2v_inst.N_429_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_16_LC_5_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101100001111"
        )
    port map (
            in0 => \N__10144\,
            in1 => \N__13709\,
            in2 => \N__10220\,
            in3 => \N__10217\,
            lcout => \b2v_inst.stateZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22517\,
            ce => 'H',
            sr => \N__22898\
        );

    \b2v_inst.state_2_LC_5_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__14321\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10184\,
            lcout => \b2v_inst.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22517\,
            ce => 'H',
            sr => \N__22898\
        );

    \b2v_inst.data_a_escribir9_4_c_RNO_LC_5_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__11094\,
            in1 => \N__11121\,
            in2 => \N__10984\,
            in3 => \N__10242\,
            lcout => \b2v_inst.data_a_escribir9_4_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.reg_ancho_3_0_LC_5_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15594\,
            in2 => \_gnd_net_\,
            in3 => \N__13085\,
            lcout => \b2v_inst.reg_ancho_3Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22406\,
            ce => \N__16045\,
            sr => \N__22902\
        );

    \b2v_inst.reg_ancho_3_1_LC_5_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__15595\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13010\,
            lcout => \b2v_inst.reg_ancho_3Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22406\,
            ce => \N__16045\,
            sr => \N__22902\
        );

    \b2v_inst.reg_ancho_3_2_LC_5_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15596\,
            in2 => \_gnd_net_\,
            in3 => \N__12941\,
            lcout => \b2v_inst.reg_ancho_3Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22406\,
            ce => \N__16045\,
            sr => \N__22902\
        );

    \b2v_inst.reg_ancho_3_3_LC_5_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__15597\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12869\,
            lcout => \b2v_inst.reg_ancho_3Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22406\,
            ce => \N__16045\,
            sr => \N__22902\
        );

    \b2v_inst.reg_ancho_3_7_LC_5_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15599\,
            in2 => \_gnd_net_\,
            in3 => \N__13619\,
            lcout => \b2v_inst.reg_ancho_3Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22406\,
            ce => \N__16045\,
            sr => \N__22902\
        );

    \b2v_inst.data_a_escribir9_5_c_RNO_LC_5_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__12784\,
            in1 => \N__12808\,
            in2 => \N__10756\,
            in3 => \N__10905\,
            lcout => \b2v_inst.data_a_escribir9_5_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.reg_ancho_3_4_LC_5_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15598\,
            in2 => \_gnd_net_\,
            in3 => \N__13535\,
            lcout => \b2v_inst.reg_ancho_3Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22406\,
            ce => \N__16045\,
            sr => \N__22902\
        );

    \b2v_inst.data_a_escribir_RNO_0_6_LC_5_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011101110"
        )
    port map (
            in0 => \N__10567\,
            in1 => \N__10845\,
            in2 => \N__11267\,
            in3 => \N__10701\,
            lcout => \b2v_inst.un1_m3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_1_6_LC_5_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001010101"
        )
    port map (
            in0 => \N__10628\,
            in1 => \N__14204\,
            in2 => \_gnd_net_\,
            in3 => \N__10619\,
            lcout => OPEN,
            ltout => \b2v_inst.data_a_escribir_RNO_1Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_6_LC_5_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__10589\,
            in1 => \N__10583\,
            in2 => \N__10574\,
            in3 => \N__10433\,
            lcout => b2v_inst_data_a_escribir_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22573\,
            ce => \N__10351\,
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNO_2_7_LC_5_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100100011"
        )
    port map (
            in0 => \N__13233\,
            in1 => \N__10568\,
            in2 => \N__10757\,
            in3 => \N__13602\,
            lcout => OPEN,
            ltout => \b2v_inst.un1_reg_anterior_iv_0_0_3_0_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_7_LC_5_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100100011"
        )
    port map (
            in0 => \N__10432\,
            in1 => \N__10376\,
            in2 => \N__10367\,
            in3 => \N__10364\,
            lcout => b2v_inst_data_a_escribir_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22573\,
            ce => \N__10351\,
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final5_0_cry_0_c_inv_LC_5_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10294\,
            in2 => \N__12763\,
            in3 => \N__10246\,
            lcout => \b2v_inst.reg_ancho_3_i_0\,
            ltout => OPEN,
            carryin => \bfn_5_17_0_\,
            carryout => \b2v_inst.valor_max_final5_0_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final5_0_cry_1_c_inv_LC_5_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11168\,
            in2 => \N__12736\,
            in3 => \N__11125\,
            lcout => \b2v_inst.reg_ancho_3_i_1\,
            ltout => OPEN,
            carryin => \b2v_inst.valor_max_final5_0_cry_0\,
            carryout => \b2v_inst.valor_max_final5_0_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final5_0_cry_2_c_inv_LC_5_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__11098\,
            in1 => \N__11074\,
            in2 => \N__12703\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst.reg_ancho_3_i_2\,
            ltout => OPEN,
            carryin => \b2v_inst.valor_max_final5_0_cry_1\,
            carryout => \b2v_inst.valor_max_final5_0_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final5_0_cry_3_c_inv_LC_5_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11033\,
            in2 => \N__12676\,
            in3 => \N__10980\,
            lcout => \b2v_inst.reg_ancho_3_i_3\,
            ltout => OPEN,
            carryin => \b2v_inst.valor_max_final5_0_cry_2\,
            carryout => \b2v_inst.valor_max_final5_0_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final5_0_cry_4_c_inv_LC_5_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10958\,
            in2 => \N__12643\,
            in3 => \N__10909\,
            lcout => \b2v_inst.reg_ancho_3_i_4\,
            ltout => OPEN,
            carryin => \b2v_inst.valor_max_final5_0_cry_3\,
            carryout => \b2v_inst.valor_max_final5_0_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final5_0_cry_5_c_inv_LC_5_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10886\,
            in2 => \N__12613\,
            in3 => \N__12783\,
            lcout => \b2v_inst.reg_ancho_3_i_5\,
            ltout => OPEN,
            carryin => \b2v_inst.valor_max_final5_0_cry_4\,
            carryout => \b2v_inst.valor_max_final5_0_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final5_0_cry_6_c_inv_LC_5_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10846\,
            in2 => \N__12583\,
            in3 => \N__12807\,
            lcout => \b2v_inst.reg_ancho_3_i_6\,
            ltout => OPEN,
            carryin => \b2v_inst.valor_max_final5_0_cry_5\,
            carryout => \b2v_inst.valor_max_final5_0_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final5_0_cry_7_c_inv_LC_5_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10801\,
            in2 => \N__13267\,
            in3 => \N__10752\,
            lcout => \b2v_inst.reg_ancho_3_i_7\,
            ltout => OPEN,
            carryin => \b2v_inst.valor_max_final5_0_cry_6\,
            carryout => \b2v_inst.valor_max_final50\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.valor_max_final50_THRU_LUT4_0_LC_5_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10730\,
            lcout => \b2v_inst.valor_max_final50_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir9_6_c_RNO_LC_5_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__12914\,
            in1 => \N__12986\,
            in2 => \N__12847\,
            in3 => \N__13058\,
            lcout => \b2v_inst.data_a_escribir9_6_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final5_2_cry_0_c_LC_5_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11512\,
            in2 => \N__12767\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_19_0_\,
            carryout => \b2v_inst.valor_max_final5_2_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final5_2_cry_1_c_LC_5_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11474\,
            in2 => \N__12737\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.valor_max_final5_2_cry_0\,
            carryout => \b2v_inst.valor_max_final5_2_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final5_2_cry_2_c_LC_5_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11428\,
            in2 => \N__12707\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.valor_max_final5_2_cry_1\,
            carryout => \b2v_inst.valor_max_final5_2_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final5_2_cry_3_c_LC_5_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11388\,
            in2 => \N__12677\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.valor_max_final5_2_cry_2\,
            carryout => \b2v_inst.valor_max_final5_2_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final5_2_cry_4_c_LC_5_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11344\,
            in2 => \N__12647\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.valor_max_final5_2_cry_3\,
            carryout => \b2v_inst.valor_max_final5_2_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final5_2_cry_5_c_LC_5_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11309\,
            in2 => \N__12617\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.valor_max_final5_2_cry_4\,
            carryout => \b2v_inst.valor_max_final5_2_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final5_2_cry_6_c_LC_5_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11262\,
            in2 => \N__12587\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.valor_max_final5_2_cry_5\,
            carryout => \b2v_inst.valor_max_final5_2_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_valor_max_final5_2_cry_7_c_LC_5_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11221\,
            in2 => \N__13271\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.valor_max_final5_2_cry_6\,
            carryout => \b2v_inst.valor_max_final52\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.valor_max_final52_THRU_LUT4_0_LC_5_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11639\,
            lcout => \b2v_inst.valor_max_final52_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst3.bit_counter_2_LC_6_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__13380\,
            in1 => \N__11589\,
            in2 => \_gnd_net_\,
            in3 => \N__11609\,
            lcout => \b2v_inst3.bit_counterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22419\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst3.bit_counter_1_LC_6_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011000001100"
        )
    port map (
            in0 => \N__13356\,
            in1 => \N__11573\,
            in2 => \N__13382\,
            in3 => \N__13304\,
            lcout => \b2v_inst3.bit_counterZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22419\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst3.bit_counter_RNIHGA63_1_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__11572\,
            in1 => \N__13302\,
            in2 => \_gnd_net_\,
            in3 => \N__13355\,
            lcout => \b2v_inst3.un1_bit_counter_3_c2\,
            ltout => \b2v_inst3.un1_bit_counter_3_c2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst3.bit_counter_3_LC_6_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010101000000"
        )
    port map (
            in0 => \N__13379\,
            in1 => \N__11591\,
            in2 => \N__11603\,
            in3 => \N__11551\,
            lcout => \b2v_inst3.bit_counterZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22419\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst3.bit_counter_RNIUR5G1_3_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__11590\,
            in1 => \N__11571\,
            in2 => \N__11552\,
            in3 => \N__13300\,
            lcout => \b2v_inst3.N_258\,
            ltout => \b2v_inst3.N_258_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst3.fsm_state_RNIEPSN1_0_LC_6_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101111111"
        )
    port map (
            in0 => \N__18841\,
            in1 => \N__12161\,
            in2 => \N__11594\,
            in3 => \N__12242\,
            lcout => \b2v_inst3.fsm_state_RNIEPSN1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst3.bit_counter_RNIVT2O_1_LC_6_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11588\,
            in2 => \_gnd_net_\,
            in3 => \N__11570\,
            lcout => OPEN,
            ltout => \b2v_inst3.N_102_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst3.bit_counter_RNIL1PJ1_3_LC_6_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__13301\,
            in1 => \N__12160\,
            in2 => \N__11555\,
            in3 => \N__11550\,
            lcout => \b2v_inst3.N_436\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst3.txd_reg_LC_6_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110010111011"
        )
    port map (
            in0 => \N__13427\,
            in1 => \N__12165\,
            in2 => \_gnd_net_\,
            in3 => \N__12241\,
            lcout => uart_tx_o,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22263\,
            ce => 'H',
            sr => \N__22885\
        );

    \b2v_inst.state_4_LC_6_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15902\,
            in2 => \_gnd_net_\,
            in3 => \N__15866\,
            lcout => \SYNTHESIZED_WIRE_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22263\,
            ce => 'H',
            sr => \N__22885\
        );

    \b2v_inst.state_fast_17_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__15867\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15903\,
            lcout => \b2v_inst.state_fastZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22263\,
            ce => 'H',
            sr => \N__22885\
        );

    \b2v_inst.state_13_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15080\,
            lcout => \b2v_inst.stateZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22263\,
            ce => 'H',
            sr => \N__22885\
        );

    \b2v_inst4.state_0_LC_6_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11706\,
            in2 => \_gnd_net_\,
            in3 => \N__15725\,
            lcout => \b2v_inst4.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22263\,
            ce => 'H',
            sr => \N__22885\
        );

    \b2v_inst3.cycle_counter_0_LC_6_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__14342\,
            in1 => \N__13350\,
            in2 => \_gnd_net_\,
            in3 => \N__12117\,
            lcout => \b2v_inst3.cycle_counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22514\,
            ce => 'H',
            sr => \N__22890\
        );

    \b2v_inst3.cycle_counter_1_LC_6_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101011110000"
        )
    port map (
            in0 => \N__12116\,
            in1 => \_gnd_net_\,
            in2 => \N__12200\,
            in3 => \N__14343\,
            lcout => \b2v_inst3.cycle_counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22514\,
            ce => 'H',
            sr => \N__22890\
        );

    \b2v_inst3.cycle_counter_RNIVMHJ_1_LC_6_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12193\,
            in2 => \_gnd_net_\,
            in3 => \N__12114\,
            lcout => \b2v_inst3.next_bit_0_a3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst3.cycle_counter_RNII2471_7_LC_6_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__11688\,
            in1 => \N__11669\,
            in2 => \N__11654\,
            in3 => \N__12033\,
            lcout => OPEN,
            ltout => \b2v_inst3.next_bit_0_a3_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst3.cycle_counter_RNIKK7E2_3_LC_6_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__12056\,
            in1 => \N__12079\,
            in2 => \N__12287\,
            in3 => \N__12284\,
            lcout => \b2v_inst3.N_105_7\,
            ltout => \b2v_inst3.N_105_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst3.fsm_state_RNI3QCR2_0_LC_6_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011100010"
        )
    port map (
            in0 => \N__12264\,
            in1 => \N__12172\,
            in2 => \N__12245\,
            in3 => \N__12236\,
            lcout => \b2v_inst3.un2_n_fsm_state_0_sqmuxa_2_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst3.cycle_counter_RNIC1OQ_1_LC_6_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000000000"
        )
    port map (
            in0 => \N__12237\,
            in1 => \N__12194\,
            in2 => \N__12176\,
            in3 => \N__12115\,
            lcout => \b2v_inst3.un1_cycle_counter_5_c2\,
            ltout => \b2v_inst3.un1_cycle_counter_5_c2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst3.cycle_counter_4_LC_6_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__12080\,
            in1 => \N__12057\,
            in2 => \N__12038\,
            in3 => \N__12034\,
            lcout => \b2v_inst3.cycle_counterZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22514\,
            ce => 'H',
            sr => \N__22890\
        );

    \b2v_inst4.pix_count_int_9_LC_6_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__12020\,
            in1 => \N__11984\,
            in2 => \N__11948\,
            in3 => \N__11882\,
            lcout => \SYNTHESIZED_WIRE_2_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22230\,
            ce => 'H',
            sr => \N__22894\
        );

    \b2v_inst.cuenta_RNIQI4F_2_LC_6_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__13757\,
            in1 => \N__13670\,
            in2 => \_gnd_net_\,
            in3 => \N__13804\,
            lcout => \b2v_inst.cuenta_RNIQI4FZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.cuenta_RNIR03A_1_LC_6_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13803\,
            in2 => \_gnd_net_\,
            in3 => \N__13758\,
            lcout => \b2v_inst.cuenta_RNIR03AZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.cuenta_pixel_RNI1NM11_6_LC_6_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111111111"
        )
    port map (
            in0 => \N__12500\,
            in1 => \_gnd_net_\,
            in2 => \N__12452\,
            in3 => \N__11844\,
            lcout => \b2v_inst.un11_cuenta_pixel_i_0_o2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.cuenta_pixel_RNO_0_6_LC_6_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__11768\,
            in1 => \N__12499\,
            in2 => \_gnd_net_\,
            in3 => \N__12448\,
            lcout => \b2v_inst.cuenta_pixel_4_i_a2_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNI95JL_3_LC_6_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__14549\,
            in1 => \N__17666\,
            in2 => \_gnd_net_\,
            in3 => \N__17018\,
            lcout => \N_213_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNIB7JL_5_LC_6_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__17019\,
            in1 => \N__14489\,
            in2 => \_gnd_net_\,
            in3 => \N__17668\,
            lcout => \N_209_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNIC8JL_6_LC_6_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__14456\,
            in1 => \N__17667\,
            in2 => \_gnd_net_\,
            in3 => \N__17020\,
            lcout => \N_207_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNIJV55_11_LC_6_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18937\,
            in2 => \_gnd_net_\,
            in3 => \N__14094\,
            lcout => \b2v_inst.N_136_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_RX_Byte_2_LC_6_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__17189\,
            in1 => \N__12349\,
            in2 => \N__22746\,
            in3 => \N__17171\,
            lcout => \SYNTHESIZED_WIRE_10_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22516\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_RX_Byte_3_LC_6_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__17172\,
            in1 => \N__12337\,
            in2 => \N__22748\,
            in3 => \N__14573\,
            lcout => \SYNTHESIZED_WIRE_10_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22516\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_RX_Byte_4_LC_6_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__14561\,
            in1 => \N__12325\,
            in2 => \N__22747\,
            in3 => \N__17173\,
            lcout => \SYNTHESIZED_WIRE_10_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22516\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_RX_Byte_5_LC_6_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__17174\,
            in1 => \N__12313\,
            in2 => \N__22749\,
            in3 => \N__15251\,
            lcout => \SYNTHESIZED_WIRE_10_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22516\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_RX_Byte_6_LC_6_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__13115\,
            in1 => \N__22733\,
            in2 => \N__12302\,
            in3 => \N__17175\,
            lcout => \SYNTHESIZED_WIRE_10_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22516\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_RX_Byte_7_LC_6_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__17176\,
            in1 => \N__12556\,
            in2 => \N__22750\,
            in3 => \N__18278\,
            lcout => \SYNTHESIZED_WIRE_10_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22516\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_3_RNIGC1F1_5_LC_6_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111011101"
        )
    port map (
            in0 => \N__15146\,
            in1 => \N__12509\,
            in2 => \N__14150\,
            in3 => \N__16951\,
            lcout => OPEN,
            ltout => \b2v_inst.addr_ram_1_iv_i_2_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_RNIBUK83_5_LC_6_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__16409\,
            in1 => \N__12515\,
            in2 => \N__12545\,
            in3 => \N__19264\,
            lcout => \N_54\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_1_RNI1SAQ_5_LC_6_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__19979\,
            in1 => \N__16473\,
            in2 => \N__16697\,
            in3 => \N__15375\,
            lcout => \b2v_inst.addr_ram_1_iv_i_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNILLMH_6_LC_6_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__15181\,
            in1 => \N__15846\,
            in2 => \_gnd_net_\,
            in3 => \N__20478\,
            lcout => \b2v_inst.N_341\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_5_LC_6_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15183\,
            lcout => \b2v_inst.stateZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22454\,
            ce => 'H',
            sr => \N__22903\
        );

    \b2v_inst.state_RNI7PTB_6_LC_6_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__15180\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15844\,
            lcout => \b2v_inst.N_238\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNIEG2F_6_LC_6_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__15845\,
            in1 => \N__15182\,
            in2 => \_gnd_net_\,
            in3 => \N__17882\,
            lcout => OPEN,
            ltout => \b2v_inst.N_404_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_3_RNI42DC1_0_LC_6_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011111111"
        )
    port map (
            in0 => \N__16950\,
            in1 => \N__14156\,
            in2 => \N__12503\,
            in3 => \N__15145\,
            lcout => \b2v_inst.addr_ram_1_iv_i_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.reg_ancho_3_6_LC_6_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__15577\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14231\,
            lcout => \b2v_inst.reg_ancho_3Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22572\,
            ce => \N__16046\,
            sr => \N__22908\
        );

    \b2v_inst.reg_ancho_3_5_LC_6_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14694\,
            in2 => \_gnd_net_\,
            in3 => \N__15576\,
            lcout => \b2v_inst.reg_ancho_3Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22572\,
            ce => \N__16046\,
            sr => \N__22908\
        );

    \b2v_inst.encontrar_maximo_un3_valor_max2_cry_0_c_LC_6_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13060\,
            in2 => \N__12762\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_17_0_\,
            carryout => \b2v_inst.un3_valor_max2_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_un3_valor_max2_cry_1_c_LC_6_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12991\,
            in2 => \N__12735\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.un3_valor_max2_cry_0\,
            carryout => \b2v_inst.un3_valor_max2_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_un3_valor_max2_cry_2_c_LC_6_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12919\,
            in2 => \N__12702\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.un3_valor_max2_cry_1\,
            carryout => \b2v_inst.un3_valor_max2_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_un3_valor_max2_cry_3_c_LC_6_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12846\,
            in2 => \N__12675\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.un3_valor_max2_cry_2\,
            carryout => \b2v_inst.un3_valor_max2_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_un3_valor_max2_cry_4_c_LC_6_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13513\,
            in2 => \N__12642\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.un3_valor_max2_cry_3\,
            carryout => \b2v_inst.un3_valor_max2_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_un3_valor_max2_cry_5_c_LC_6_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14659\,
            in2 => \N__12612\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.un3_valor_max2_cry_4\,
            carryout => \b2v_inst.un3_valor_max2_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_un3_valor_max2_cry_6_c_LC_6_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14200\,
            in2 => \N__12582\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.un3_valor_max2_cry_5\,
            carryout => \b2v_inst.un3_valor_max2_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.encontrar_maximo_un3_valor_max2_cry_7_c_LC_6_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13601\,
            in2 => \N__13266\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst.un3_valor_max2_cry_6\,
            carryout => \b2v_inst.un3_valor_max2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.un3_valor_max2_THRU_LUT4_0_LC_6_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13241\,
            lcout => \b2v_inst.un3_valor_max2_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst3.fsm_state_RNI6DTR2_0_LC_6_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13141\,
            in2 => \_gnd_net_\,
            in3 => \N__13127\,
            lcout => \b2v_inst3.un2_n_fsm_state_0_sqmuxa_2_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_RX_Byte_RNO_0_6_LC_6_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__18260\,
            in1 => \N__18184\,
            in2 => \_gnd_net_\,
            in3 => \N__18125\,
            lcout => \b2v_inst1.r_RX_Bytece_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.reg_anterior_0_LC_6_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15559\,
            in2 => \_gnd_net_\,
            in3 => \N__13102\,
            lcout => \b2v_inst.reg_anteriorZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22244\,
            ce => \N__15239\,
            sr => \N__22914\
        );

    \b2v_inst.reg_anterior_1_LC_6_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101000001010"
        )
    port map (
            in0 => \N__13027\,
            in1 => \_gnd_net_\,
            in2 => \N__15575\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst.reg_anteriorZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22244\,
            ce => \N__15239\,
            sr => \N__22914\
        );

    \b2v_inst.reg_anterior_2_LC_6_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15563\,
            in2 => \_gnd_net_\,
            in3 => \N__12958\,
            lcout => \b2v_inst.reg_anteriorZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22244\,
            ce => \N__15239\,
            sr => \N__22914\
        );

    \b2v_inst.reg_anterior_3_LC_6_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__15564\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12886\,
            lcout => \b2v_inst.reg_anteriorZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22244\,
            ce => \N__15239\,
            sr => \N__22914\
        );

    \b2v_inst.reg_anterior_7_LC_6_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15566\,
            in2 => \_gnd_net_\,
            in3 => \N__13643\,
            lcout => \b2v_inst.reg_anteriorZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22244\,
            ce => \N__15239\,
            sr => \N__22914\
        );

    \b2v_inst.data_a_escribir9_7_c_RNO_LC_6_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__14198\,
            in1 => \N__14648\,
            in2 => \N__13603\,
            in3 => \N__13508\,
            lcout => \b2v_inst.data_a_escribir9_7_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.reg_anterior_4_LC_6_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__13552\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15565\,
            lcout => \b2v_inst.reg_anteriorZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22244\,
            ce => \N__15239\,
            sr => \N__22914\
        );

    \b2v_inst3.data_to_send_esr_1_LC_6_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000000100010"
        )
    port map (
            in0 => \N__13481\,
            in1 => \N__14419\,
            in2 => \N__13391\,
            in3 => \N__14341\,
            lcout => \b2v_inst3.data_to_sendZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22571\,
            ce => \N__14258\,
            sr => \N__22918\
        );

    \b2v_inst3.data_to_send_esr_0_LC_6_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000000100010"
        )
    port map (
            in0 => \N__13460\,
            in1 => \N__14418\,
            in2 => \N__13436\,
            in3 => \N__14340\,
            lcout => \b2v_inst3.data_to_sendZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22571\,
            ce => \N__14258\,
            sr => \N__22918\
        );

    \b2v_inst3.data_to_send_esr_2_LC_6_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011011000"
        )
    port map (
            in0 => \N__14339\,
            in1 => \N__14525\,
            in2 => \N__13415\,
            in3 => \N__14420\,
            lcout => \b2v_inst3.data_to_sendZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22571\,
            ce => \N__14258\,
            sr => \N__22918\
        );

    \b2v_inst3.bit_counter_0_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__13381\,
            in1 => \N__13303\,
            in2 => \_gnd_net_\,
            in3 => \N__13358\,
            lcout => \b2v_inst3.bit_counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22083\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.cuenta_RNIFIIS1_4_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001111101100"
        )
    port map (
            in0 => \N__13852\,
            in1 => \N__15020\,
            in2 => \N__13280\,
            in3 => \N__14988\,
            lcout => \b2v_inst.state_ns_a2_0_o2_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.cuenta_RNIQI4F_0_2_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__13668\,
            in1 => \N__13801\,
            in2 => \_gnd_net_\,
            in3 => \N__13743\,
            lcout => \b2v_inst.state_ns_a2_0_a2_0_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.cuenta_RNIQ56K_0_3_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__13742\,
            in1 => \N__13666\,
            in2 => \N__13805\,
            in3 => \N__13686\,
            lcout => \b2v_inst.cuenta_RNIQ56K_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.cuenta_RNO_0_0_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100110011"
        )
    port map (
            in0 => \N__18707\,
            in1 => \N__13745\,
            in2 => \N__17700\,
            in3 => \N__14606\,
            lcout => OPEN,
            ltout => \b2v_inst.cuenta_5_i_a2_2_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.cuenta_0_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101011111000"
        )
    port map (
            in0 => \N__14859\,
            in1 => \N__16217\,
            in2 => \N__13694\,
            in3 => \N__16168\,
            lcout => \b2v_inst.cuentaZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21947\,
            ce => \N__14905\,
            sr => \N__22891\
        );

    \b2v_inst.cuenta_RNIQ56K_3_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__13665\,
            in1 => \N__13796\,
            in2 => \N__13688\,
            in3 => \N__13741\,
            lcout => \b2v_inst.un4_cuenta_c4\,
            ltout => \b2v_inst.un4_cuenta_c4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.cuenta_4_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000101000"
        )
    port map (
            in0 => \N__17683\,
            in1 => \N__15021\,
            in2 => \N__13691\,
            in3 => \N__18708\,
            lcout => \b2v_inst.cuentaZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21947\,
            ce => \N__14905\,
            sr => \N__22891\
        );

    \b2v_inst.cuenta_RNO_1_3_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__13667\,
            in1 => \N__13800\,
            in2 => \_gnd_net_\,
            in3 => \N__13744\,
            lcout => \b2v_inst.cuenta_5_i_a2_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.cuenta_3_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__13853\,
            in1 => \N__13718\,
            in2 => \_gnd_net_\,
            in3 => \N__14585\,
            lcout => \b2v_inst.cuentaZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22084\,
            ce => \N__14898\,
            sr => \N__22895\
        );

    \b2v_inst.cuenta_2_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010001000100"
        )
    port map (
            in0 => \N__14584\,
            in1 => \N__13829\,
            in2 => \N__13820\,
            in3 => \N__13835\,
            lcout => \b2v_inst.cuentaZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22084\,
            ce => \N__14898\,
            sr => \N__22895\
        );

    \b2v_inst.cuenta_fast_RNIBDJQ_4_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__13687\,
            in1 => \N__13669\,
            in2 => \N__13868\,
            in3 => \N__13802\,
            lcout => \b2v_inst.un2_cuentalto7_3\,
            ltout => \b2v_inst.un2_cuentalto7_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.cuenta_RNIKFO91_7_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__14925\,
            in1 => \N__14953\,
            in2 => \N__13874\,
            in3 => \N__15058\,
            lcout => \b2v_inst.N_351_0\,
            ltout => \b2v_inst.N_351_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.cuenta_fast_4_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000001000001000"
        )
    port map (
            in0 => \N__17669\,
            in1 => \N__13867\,
            in2 => \N__13871\,
            in3 => \N__14989\,
            lcout => \b2v_inst.cuenta_fastZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22084\,
            ce => \N__14898\,
            sr => \N__22895\
        );

    \b2v_inst.cuenta_RNI1OL72_0_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001010"
        )
    port map (
            in0 => \N__13851\,
            in1 => \N__18709\,
            in2 => \N__17701\,
            in3 => \N__13760\,
            lcout => \b2v_inst.N_376_1\,
            ltout => \b2v_inst.N_376_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.cuenta_1_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001001100"
        )
    port map (
            in0 => \N__13828\,
            in1 => \N__13816\,
            in2 => \N__13808\,
            in3 => \N__14583\,
            lcout => \b2v_inst.cuentaZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22084\,
            ce => \N__14898\,
            sr => \N__22895\
        );

    \b2v_inst.cuenta_RNO_0_3_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001010"
        )
    port map (
            in0 => \N__13769\,
            in1 => \N__18703\,
            in2 => \N__17692\,
            in3 => \N__13759\,
            lcout => \b2v_inst.N_377\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNIP7VJ_10_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__13892\,
            in1 => \N__15477\,
            in2 => \N__15224\,
            in3 => \N__16024\,
            lcout => \b2v_inst.N_491\,
            ltout => \b2v_inst.N_491_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNIFQKO_17_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13712\,
            in3 => \N__17639\,
            lcout => \b2v_inst.state_RNIFQKOZ0Z_17\,
            ltout => \b2v_inst.state_RNIFQKOZ0Z_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNIFQKO_0_17_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13697\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst.N_399_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNIDVTB_9_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16023\,
            in2 => \_gnd_net_\,
            in3 => \N__13962\,
            lcout => \b2v_inst.N_236\,
            ltout => \b2v_inst.N_236_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_8_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010000010110000"
        )
    port map (
            in0 => \N__13963\,
            in1 => \N__16077\,
            in2 => \N__13973\,
            in3 => \N__14824\,
            lcout => \b2v_inst.stateZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22554\,
            ce => 'H',
            sr => \N__22899\
        );

    \b2v_inst.state_17_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__15865\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15910\,
            lcout => \b2v_inst.stateZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22554\,
            ce => 'H',
            sr => \N__22899\
        );

    \b2v_inst.state_9_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101000"
        )
    port map (
            in0 => \N__13893\,
            in1 => \N__16076\,
            in2 => \N__16229\,
            in3 => \N__16173\,
            lcout => \b2v_inst.stateZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22554\,
            ce => 'H',
            sr => \N__22899\
        );

    \b2v_inst.dir_mem_1_RNI3UAQ_6_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__16286\,
            in1 => \N__16465\,
            in2 => \N__14111\,
            in3 => \N__15369\,
            lcout => \b2v_inst.addr_ram_1_iv_i_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNIMMMH_6_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__15184\,
            in1 => \N__15847\,
            in2 => \_gnd_net_\,
            in3 => \N__20631\,
            lcout => OPEN,
            ltout => \b2v_inst.N_399_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_3_RNIIE1F1_6_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111110011"
        )
    port map (
            in0 => \N__14135\,
            in1 => \N__15139\,
            in2 => \N__13949\,
            in3 => \N__16936\,
            lcout => OPEN,
            ltout => \b2v_inst.addr_ram_1_iv_i_2_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_RNIG3L83_6_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__16395\,
            in1 => \N__13946\,
            in2 => \N__13940\,
            in3 => \N__19127\,
            lcout => \N_165\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_12_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100010001100"
        )
    port map (
            in0 => \N__15946\,
            in1 => \N__15370\,
            in2 => \N__16115\,
            in3 => \N__14820\,
            lcout => \b2v_inst.stateZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22589\,
            ce => 'H',
            sr => \N__22904\
        );

    \b2v_inst.state_RNI3SA9_13_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15945\,
            in2 => \_gnd_net_\,
            in3 => \N__13894\,
            lcout => \b2v_inst.N_235\,
            ltout => \b2v_inst.N_235_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_1_RNIKA1U_7_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__15287\,
            in1 => \N__18041\,
            in2 => \N__14099\,
            in3 => \N__16935\,
            lcout => \b2v_inst.addr_ram_1_0_iv_i_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_10_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000000010000"
        )
    port map (
            in0 => \N__14825\,
            in1 => \N__16111\,
            in2 => \N__16480\,
            in3 => \N__14096\,
            lcout => \b2v_inst.stateZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22352\,
            ce => 'H',
            sr => \N__22909\
        );

    \b2v_inst.dir_mem_1_RNIPJAQ_1_LC_7_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__19949\,
            in1 => \N__16466\,
            in2 => \N__16526\,
            in3 => \N__15371\,
            lcout => \b2v_inst.addr_ram_1_0_iv_i_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNIVNA9_11_LC_7_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14095\,
            in2 => \_gnd_net_\,
            in3 => \N__15469\,
            lcout => \b2v_inst.N_237\,
            ltout => \b2v_inst.N_237_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_1_RNINHAQ_0_LC_7_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__16493\,
            in1 => \N__20162\,
            in2 => \N__14072\,
            in3 => \N__15372\,
            lcout => OPEN,
            ltout => \b2v_inst.addr_ram_1_iv_i_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_RNIG4063_0_LC_7_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__19895\,
            in1 => \N__14069\,
            in2 => \N__14063\,
            in3 => \N__16396\,
            lcout => \N_167\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_RNIQQMS2_1_LC_7_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011101110"
        )
    port map (
            in0 => \N__14162\,
            in1 => \N__14033\,
            in2 => \N__16405\,
            in3 => \N__19817\,
            lcout => \N_60\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_1_RNIRLAQ_2_LC_7_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__15373\,
            in1 => \N__16508\,
            in2 => \N__16479\,
            in3 => \N__20000\,
            lcout => OPEN,
            ltout => \b2v_inst.addr_ram_1_0_iv_i_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_RNIVVMS2_2_LC_7_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__16400\,
            in1 => \N__16880\,
            in2 => \N__14003\,
            in3 => \N__19217\,
            lcout => \N_56\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_RNI88AO1_7_LC_7_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111110101"
        )
    port map (
            in0 => \N__20936\,
            in1 => \N__20632\,
            in2 => \N__17900\,
            in3 => \N__20503\,
            lcout => \b2v_inst.dir_mem_315_0\,
            ltout => \b2v_inst.dir_mem_315_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_3_1_LC_7_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110100101"
        )
    port map (
            in0 => \N__23027\,
            in1 => \_gnd_net_\,
            in2 => \N__14171\,
            in3 => \N__23211\,
            lcout => \b2v_inst.dir_mem_3Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22595\,
            ce => \N__15274\,
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_3_2_LC_7_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101010011001"
        )
    port map (
            in0 => \N__20147\,
            in1 => \N__23028\,
            in2 => \N__23219\,
            in3 => \N__15316\,
            lcout => \b2v_inst.dir_mem_3Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22595\,
            ce => \N__15274\,
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_3_RNIBL331_1_LC_7_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__16952\,
            in1 => \N__14168\,
            in2 => \N__23054\,
            in3 => \N__17000\,
            lcout => \b2v_inst.addr_ram_1_0_iv_i_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_3_0_LC_7_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__23210\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15315\,
            lcout => \b2v_inst.dir_mem_3Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22595\,
            ce => \N__15274\,
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_3_5_LC_7_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001010110101001"
        )
    port map (
            in0 => \N__20504\,
            in1 => \N__16247\,
            in2 => \N__15325\,
            in3 => \N__18027\,
            lcout => \b2v_inst.dir_mem_3Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22595\,
            ce => \N__15274\,
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_3_4_LC_7_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011001011010"
        )
    port map (
            in0 => \N__18026\,
            in1 => \N__20825\,
            in2 => \N__15980\,
            in3 => \N__15317\,
            lcout => \b2v_inst.dir_mem_3Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22595\,
            ce => \N__15274\,
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_3_6_LC_7_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101011010100110"
        )
    port map (
            in0 => \N__20633\,
            in1 => \N__16274\,
            in2 => \N__15326\,
            in3 => \N__16553\,
            lcout => \b2v_inst.dir_mem_3Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22595\,
            ce => \N__15274\,
            sr => \_gnd_net_\
        );

    \b2v_inst.data_a_escribir_RNID9JL_7_LC_7_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__17679\,
            in1 => \N__14371\,
            in2 => \_gnd_net_\,
            in3 => \N__17017\,
            lcout => \N_205_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_2_6_LC_7_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__20354\,
            in1 => \N__16732\,
            in2 => \_gnd_net_\,
            in3 => \N__15731\,
            lcout => \b2v_inst.dir_mem_2Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22354\,
            ce => \N__16682\,
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_RX_Byte_RNO_0_3_LC_7_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__18163\,
            in1 => \N__18251\,
            in2 => \_gnd_net_\,
            in3 => \N__18123\,
            lcout => \b2v_inst1.r_RX_Bytece_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_RX_Byte_RNO_0_4_LC_7_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__18124\,
            in1 => \_gnd_net_\,
            in2 => \N__18259\,
            in3 => \N__18164\,
            lcout => \b2v_inst1.r_RX_Bytece_0_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst3.data_to_send_esr_3_LC_7_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__14413\,
            in1 => \N__14545\,
            in2 => \N__14498\,
            in3 => \N__14346\,
            lcout => \b2v_inst3.data_to_sendZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22242\,
            ce => \N__14254\,
            sr => \N__22915\
        );

    \b2v_inst3.data_to_send_esr_4_LC_7_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011100100"
        )
    port map (
            in0 => \N__14344\,
            in1 => \N__14516\,
            in2 => \N__14465\,
            in3 => \N__14414\,
            lcout => \b2v_inst3.data_to_sendZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22242\,
            ce => \N__14254\,
            sr => \N__22915\
        );

    \b2v_inst3.data_to_send_esr_5_LC_7_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__14415\,
            in1 => \N__14485\,
            in2 => \N__14429\,
            in3 => \N__14347\,
            lcout => \b2v_inst3.data_to_sendZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22242\,
            ce => \N__14254\,
            sr => \N__22915\
        );

    \b2v_inst3.data_to_send_esr_6_LC_7_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011100100"
        )
    port map (
            in0 => \N__14345\,
            in1 => \N__14455\,
            in2 => \N__14270\,
            in3 => \N__14416\,
            lcout => \b2v_inst3.data_to_sendZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22242\,
            ce => \N__14254\,
            sr => \N__22915\
        );

    \b2v_inst3.data_to_send_esr_7_LC_7_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110001010000"
        )
    port map (
            in0 => \N__14417\,
            in1 => \N__14269\,
            in2 => \N__14375\,
            in3 => \N__14348\,
            lcout => \b2v_inst3.data_to_sendZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22242\,
            ce => \N__14254\,
            sr => \N__22915\
        );

    \b2v_inst.reg_anterior_6_LC_7_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__15535\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14242\,
            lcout => \b2v_inst.reg_anteriorZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22243\,
            ce => \N__15235\,
            sr => \N__22919\
        );

    \b2v_inst.reg_anterior_5_LC_7_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15534\,
            in2 => \_gnd_net_\,
            in3 => \N__14705\,
            lcout => \b2v_inst.reg_anteriorZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22243\,
            ce => \N__15235\,
            sr => \N__22919\
        );

    \b2v_inst.cuenta_RNI5B3A_6_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14952\,
            in2 => \_gnd_net_\,
            in3 => \N__15053\,
            lcout => OPEN,
            ltout => \b2v_inst.un4_cuenta_ac0_11_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.cuenta_RNI4SC81_7_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__14985\,
            in1 => \N__14924\,
            in2 => \N__14624\,
            in3 => \N__15022\,
            lcout => \b2v_inst.cuenta_RNI4SC81Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.cuenta_RNIK17D1_4_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101100110"
        )
    port map (
            in0 => \N__15026\,
            in1 => \N__14984\,
            in2 => \_gnd_net_\,
            in3 => \N__14621\,
            lcout => \b2v_inst.cuenta_5_i_o2_0_0_1\,
            ltout => \b2v_inst.cuenta_5_i_o2_0_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.cuenta_RNIO2VO3_4_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16202\,
            in2 => \N__14612\,
            in3 => \N__16150\,
            lcout => \b2v_inst.cuenta_RNIO2VO3Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.cuenta_RNI05B31_6_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111011101110"
        )
    port map (
            in0 => \N__14957\,
            in1 => \N__15054\,
            in2 => \N__15029\,
            in3 => \N__14986\,
            lcout => \b2v_inst.state_ns_a2_0_o2_1_0_2\,
            ltout => \b2v_inst.state_ns_a2_0_o2_1_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_17_rep1_RNICDK34_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010100"
        )
    port map (
            in0 => \N__19080\,
            in1 => \N__16151\,
            in2 => \N__14609\,
            in3 => \N__14605\,
            lcout => OPEN,
            ltout => \b2v_inst.state_17_rep1_RNICDKZ0Z34_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_17_rep1_RNIOVB69_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18749\,
            in2 => \N__14594\,
            in3 => \N__14591\,
            lcout => \b2v_inst.N_374\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.cuenta_5_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001111000"
        )
    port map (
            in0 => \N__14987\,
            in1 => \N__15027\,
            in2 => \N__15062\,
            in3 => \N__14858\,
            lcout => \b2v_inst.cuentaZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21971\,
            ce => \N__14906\,
            sr => \N__22896\
        );

    \b2v_inst.dir_mem_RNO_3_0_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__14927\,
            in1 => \N__14955\,
            in2 => \N__17572\,
            in3 => \N__15060\,
            lcout => \b2v_inst.un2_indice_3_0_iv_0_a2_5_sx_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.cuenta_RNI925F_7_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__14926\,
            in1 => \N__14954\,
            in2 => \_gnd_net_\,
            in3 => \N__15059\,
            lcout => \b2v_inst.cuenta_RNI925FZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.cuenta_RNO_0_6_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__15061\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15028\,
            lcout => OPEN,
            ltout => \b2v_inst.un4_cuenta_ac0_9_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.cuenta_6_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001010001000100"
        )
    port map (
            in0 => \N__14856\,
            in1 => \N__14956\,
            in2 => \N__14993\,
            in3 => \N__14990\,
            lcout => \b2v_inst.cuentaZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22187\,
            ce => \N__14897\,
            sr => \N__22900\
        );

    \b2v_inst.cuenta_7_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14857\,
            in2 => \_gnd_net_\,
            in3 => \N__16169\,
            lcout => \b2v_inst.cuentaZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22187\,
            ce => \N__14897\,
            sr => \N__22900\
        );

    \b2v_inst.state_17_rep1_RNI8QDK1_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19052\,
            in2 => \_gnd_net_\,
            in3 => \N__18699\,
            lcout => \b2v_inst.N_227\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.cuenta_RNI41OB2_6_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16221\,
            in2 => \_gnd_net_\,
            in3 => \N__16170\,
            lcout => \b2v_inst.N_232\,
            ltout => \b2v_inst.N_232_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_14_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000010"
        )
    port map (
            in0 => \N__15214\,
            in1 => \N__16101\,
            in2 => \N__14801\,
            in3 => \N__18985\,
            lcout => \b2v_inst.stateZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22468\,
            ce => 'H',
            sr => \N__22905\
        );

    \b2v_inst.state_7_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__16222\,
            in1 => \N__15215\,
            in2 => \N__16112\,
            in3 => \N__16171\,
            lcout => \b2v_inst.stateZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22468\,
            ce => 'H',
            sr => \N__22905\
        );

    \b2v_inst.state_fast_15_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__16172\,
            in1 => \N__16223\,
            in2 => \N__16044\,
            in3 => \N__16100\,
            lcout => \b2v_inst.state_fastZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22468\,
            ce => 'H',
            sr => \N__22905\
        );

    \b2v_inst.state_RNIRA0K_15_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__18984\,
            in1 => \N__19062\,
            in2 => \_gnd_net_\,
            in3 => \N__15213\,
            lcout => \b2v_inst.N_239\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_RNO_2_6_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__18918\,
            in1 => \N__19076\,
            in2 => \_gnd_net_\,
            in3 => \N__18983\,
            lcout => \b2v_inst.N_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNITETB_0_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__15073\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15439\,
            lcout => \b2v_inst.state_RNITETBZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_1_RNITNAQ_3_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__15374\,
            in1 => \N__15989\,
            in2 => \N__20210\,
            in3 => \N__16458\,
            lcout => \b2v_inst.addr_ram_1_iv_i_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNIHV0E_6_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__15185\,
            in1 => \N__15871\,
            in2 => \_gnd_net_\,
            in3 => \N__17115\,
            lcout => OPEN,
            ltout => \b2v_inst.N_351_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_3_RNIAKBB1_3_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111110011"
        )
    port map (
            in0 => \N__15296\,
            in1 => \N__15138\,
            in2 => \N__15119\,
            in3 => \N__16946\,
            lcout => OPEN,
            ltout => \b2v_inst.addr_ram_1_iv_i_2_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_RNIVVU43_3_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__16374\,
            in1 => \N__15116\,
            in2 => \N__15110\,
            in3 => \N__19322\,
            lcout => \N_58\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_0_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__15440\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22355\,
            ce => 'H',
            sr => \N__22910\
        );

    \b2v_inst.state_1_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111000000000"
        )
    port map (
            in0 => \N__16224\,
            in1 => \N__16174\,
            in2 => \N__16114\,
            in3 => \N__15470\,
            lcout => \b2v_inst.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22355\,
            ce => 'H',
            sr => \N__22910\
        );

    \b2v_inst.dir_mem_3_RNIHR331_4_LC_8_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__17012\,
            in1 => \N__16953\,
            in2 => \N__15431\,
            in3 => \N__18005\,
            lcout => OPEN,
            ltout => \b2v_inst.addr_ram_1_0_iv_i_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_RNI9ANS2_4_LC_8_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__16394\,
            in1 => \N__15332\,
            in2 => \N__15419\,
            in3 => \N__19373\,
            lcout => \N_163\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_1_RNO_1_4_LC_8_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100010001"
        )
    port map (
            in0 => \N__20492\,
            in1 => \N__20687\,
            in2 => \_gnd_net_\,
            in3 => \N__18006\,
            lcout => OPEN,
            ltout => \b2v_inst.g0_11_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_1_4_LC_8_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001101010011001"
        )
    port map (
            in0 => \N__18007\,
            in1 => \N__17912\,
            in2 => \N__15389\,
            in3 => \N__20610\,
            lcout => \b2v_inst.dir_mem_1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22351\,
            ce => \N__19920\,
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_1_RNIVPAQ_4_LC_8_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__16474\,
            in1 => \N__15386\,
            in2 => \N__16541\,
            in3 => \N__15376\,
            lcout => \b2v_inst.addr_ram_1_0_iv_i_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_3_3_LC_8_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__15761\,
            in1 => \N__17045\,
            in2 => \_gnd_net_\,
            in3 => \N__15324\,
            lcout => \b2v_inst.dir_mem_3Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22594\,
            ce => \N__15275\,
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_3_7_LC_8_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__20639\,
            in1 => \N__16270\,
            in2 => \_gnd_net_\,
            in3 => \N__20934\,
            lcout => \b2v_inst.dir_mem_3Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22594\,
            ce => \N__15275\,
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_RX_Byte_RNO_0_5_LC_8_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__18191\,
            in1 => \N__18104\,
            in2 => \_gnd_net_\,
            in3 => \N__18239\,
            lcout => \b2v_inst1.r_RX_Bytece_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_SM_Main_RNIC98H_2_LC_8_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__23483\,
            in1 => \N__23753\,
            in2 => \_gnd_net_\,
            in3 => \N__23629\,
            lcout => \b2v_inst1.r_SM_Main_d_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_3_RNO_0_3_LC_8_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010011001"
        )
    port map (
            in0 => \N__23081\,
            in1 => \N__20332\,
            in2 => \_gnd_net_\,
            in3 => \N__20140\,
            lcout => \b2v_inst.dir_mem_3_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_RX_Byte_RNO_0_1_LC_8_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__18119\,
            in1 => \N__18165\,
            in2 => \_gnd_net_\,
            in3 => \N__18255\,
            lcout => OPEN,
            ltout => \b2v_inst1.r_RX_Bytece_0_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_RX_Byte_1_LC_8_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__15742\,
            in1 => \N__22708\,
            in2 => \N__15752\,
            in3 => \N__17170\,
            lcout => \SYNTHESIZED_WIRE_10_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22353\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_2_RNO_0_6_LC_8_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011011001100"
        )
    port map (
            in0 => \N__18028\,
            in1 => \N__20636\,
            in2 => \N__17060\,
            in3 => \N__20501\,
            lcout => \b2v_inst.dir_mem_2_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_Bit_Index_0_LC_8_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011010010"
        )
    port map (
            in0 => \N__16633\,
            in1 => \N__23494\,
            in2 => \N__18185\,
            in3 => \N__23754\,
            lcout => \b2v_inst1.r_Bit_IndexZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22593\,
            ce => 'H',
            sr => \N__24063\
        );

    \b2v_inst1.r_RX_DV_LC_8_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110100011100000"
        )
    port map (
            in0 => \N__23755\,
            in1 => \N__23630\,
            in2 => \N__15719\,
            in3 => \N__16634\,
            lcout => \SYNTHESIZED_WIRE_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22593\,
            ce => 'H',
            sr => \N__24063\
        );

    \b2v_inst.ignorar_anterior_LC_8_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15684\,
            lcout => \b2v_inst.ignorar_anteriorZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22480\,
            ce => \N__15521\,
            sr => \N__22921\
        );

    \b2v_inst.dir_mem_RNO_0_6_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001010"
        )
    port map (
            in0 => \N__15797\,
            in1 => \N__15803\,
            in2 => \N__15506\,
            in3 => \N__18775\,
            lcout => OPEN,
            ltout => \b2v_inst.N_7_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_6_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__17828\,
            in1 => \N__16808\,
            in2 => \N__15809\,
            in3 => \N__16574\,
            lcout => \b2v_inst.dir_memZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22392\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_RNO_5_6_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19320\,
            in2 => \_gnd_net_\,
            in3 => \N__19213\,
            lcout => OPEN,
            ltout => \b2v_inst.g2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_RNO_3_6_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001101010"
        )
    port map (
            in0 => \N__19112\,
            in1 => \N__15926\,
            in2 => \N__15806\,
            in3 => \N__19727\,
            lcout => \b2v_inst.g1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_RNO_4_6_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010011010"
        )
    port map (
            in0 => \N__20635\,
            in1 => \N__21145\,
            in2 => \N__16829\,
            in3 => \N__21059\,
            lcout => \b2v_inst.un2_indice_21_s0_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_RNITB3H1_6_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110010011001"
        )
    port map (
            in0 => \N__20634\,
            in1 => \N__17782\,
            in2 => \N__19119\,
            in3 => \N__19726\,
            lcout => \b2v_inst.dir_mem_RNITB3H1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_3_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__20139\,
            in1 => \N__23134\,
            in2 => \N__20276\,
            in3 => \N__23084\,
            lcout => \b2v_inst.indiceZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22114\,
            ce => \N__22952\,
            sr => \N__22901\
        );

    \b2v_inst.state_fast_RNI711G_0_15_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101110111"
        )
    port map (
            in0 => \N__18916\,
            in1 => \N__15776\,
            in2 => \_gnd_net_\,
            in3 => \N__15787\,
            lcout => \b2v_inst.N_253\,
            ltout => \b2v_inst.N_253_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_RNIGVEE1_0_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__19862\,
            in1 => \N__21038\,
            in2 => \N__15791\,
            in3 => \N__17768\,
            lcout => \b2v_inst.dir_mem_RNIGVEE1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_fast_RNI711G_15_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__18917\,
            in1 => \N__15788\,
            in2 => \_gnd_net_\,
            in3 => \N__15775\,
            lcout => \b2v_inst.N_253_i\,
            ltout => \b2v_inst.N_253_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_RNII5PO1_1_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110010100101"
        )
    port map (
            in0 => \N__21146\,
            in1 => \N__19816\,
            in2 => \N__15764\,
            in3 => \N__19721\,
            lcout => \b2v_inst.dir_mem_RNII5PO1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_RNIN53H1_3_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100101111100001"
        )
    port map (
            in0 => \N__19723\,
            in1 => \N__20242\,
            in2 => \N__17790\,
            in3 => \N__19319\,
            lcout => \b2v_inst.dir_mem_RNIN53H1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_RNIL33H1_2_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011000011"
        )
    port map (
            in0 => \N__19205\,
            in1 => \N__17764\,
            in2 => \N__20146\,
            in3 => \N__19722\,
            lcout => \b2v_inst.dir_mem_RNIL33H1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_17_rep1_RNIBDUK1_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__18922\,
            in1 => \N__19066\,
            in2 => \_gnd_net_\,
            in3 => \N__18745\,
            lcout => \b2v_inst.N_467\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_RNO_0_0_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15959\,
            in2 => \_gnd_net_\,
            in3 => \N__17391\,
            lcout => OPEN,
            ltout => \b2v_inst.N_452_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_0_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001001100"
        )
    port map (
            in0 => \N__23152\,
            in1 => \N__16235\,
            in2 => \N__15953\,
            in3 => \N__17585\,
            lcout => \b2v_inst.dir_memZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22501\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNIL165_13_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18923\,
            in2 => \_gnd_net_\,
            in3 => \N__15950\,
            lcout => \b2v_inst.N_134_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_RNO_6_6_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__19372\,
            in1 => \N__19815\,
            in2 => \N__19260\,
            in3 => \N__19869\,
            lcout => \b2v_inst.g2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_17_rep1_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15914\,
            in2 => \_gnd_net_\,
            in3 => \N__15872\,
            lcout => \b2v_inst.state_17_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22318\,
            ce => 'H',
            sr => \N__22911\
        );

    \b2v_inst.dir_mem_RNO_7_0_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111111100000"
        )
    port map (
            in0 => \N__19070\,
            in1 => \N__18982\,
            in2 => \N__18939\,
            in3 => \N__19873\,
            lcout => OPEN,
            ltout => \b2v_inst.g4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_RNO_2_0_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001011111010"
        )
    port map (
            in0 => \N__18773\,
            in1 => \N__16814\,
            in2 => \N__16238\,
            in3 => \N__16301\,
            lcout => \b2v_inst.g0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNIBERF_15_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__18927\,
            in1 => \N__19048\,
            in2 => \_gnd_net_\,
            in3 => \N__18981\,
            lcout => \b2v_inst.N_451\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_15_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111000000000"
        )
    port map (
            in0 => \N__16228\,
            in1 => \N__16175\,
            in2 => \N__16113\,
            in3 => \N__16037\,
            lcout => \b2v_inst.stateZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22318\,
            ce => 'H',
            sr => \N__22911\
        );

    \b2v_inst.indice_0_rep1_RNI3OC22_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__19667\,
            in1 => \N__17486\,
            in2 => \N__17398\,
            in3 => \N__17507\,
            lcout => \b2v_inst.N_410\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_2_RNO_0_3_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__23083\,
            in1 => \N__20298\,
            in2 => \_gnd_net_\,
            in3 => \N__20117\,
            lcout => OPEN,
            ltout => \b2v_inst.dir_mem_2_RNO_0Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_2_3_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17341\,
            in2 => \N__15992\,
            in3 => \N__16733\,
            lcout => \b2v_inst.dir_mem_2Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22502\,
            ce => \N__16673\,
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_3_RNO_0_4_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__23082\,
            in1 => \N__20297\,
            in2 => \_gnd_net_\,
            in3 => \N__20116\,
            lcout => \b2v_inst.un1_dir_mem_3_ns_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_2_7_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__20604\,
            in1 => \N__20914\,
            in2 => \N__20500\,
            in3 => \N__15965\,
            lcout => \b2v_inst.dir_mem_2Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22319\,
            ce => \N__16677\,
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_2_RNO_0_7_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__18391\,
            in1 => \N__17872\,
            in2 => \N__20768\,
            in3 => \N__19673\,
            lcout => \b2v_inst.dir_mem_2_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_2_RNI8NDV_7_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__17013\,
            in1 => \N__16478\,
            in2 => \N__16418\,
            in3 => \N__20913\,
            lcout => OPEN,
            ltout => \b2v_inst.addr_ram_1_0_iv_i_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_RNIOPNS2_7_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__16401\,
            in1 => \N__19160\,
            in2 => \N__16349\,
            in3 => \N__16346\,
            lcout => \N_50\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_RNO_8_0_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__17871\,
            in1 => \N__20912\,
            in2 => \N__18395\,
            in3 => \N__18336\,
            lcout => OPEN,
            ltout => \b2v_inst.g0_2_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_RNO_6_0_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__18938\,
            in1 => \N__19082\,
            in2 => \N__16304\,
            in3 => \N__20603\,
            lcout => \b2v_inst.g0_2_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_1_RNO_0_6_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000001000"
        )
    port map (
            in0 => \N__20296\,
            in1 => \N__18004\,
            in2 => \N__16565\,
            in3 => \N__20637\,
            lcout => OPEN,
            ltout => \b2v_inst.i4_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_1_6_LC_9_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011100100"
        )
    port map (
            in0 => \N__20494\,
            in1 => \N__20638\,
            in2 => \N__16289\,
            in3 => \N__20933\,
            lcout => \b2v_inst.dir_mem_1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22569\,
            ce => \N__19926\,
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_RNI3ML81_3_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000000"
        )
    port map (
            in0 => \N__20294\,
            in1 => \N__18002\,
            in2 => \N__16259\,
            in3 => \N__20493\,
            lcout => \b2v_inst.un2_dir_mem_3_c5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_3_rep1_RNIS3BN_LC_9_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__17116\,
            in1 => \N__19514\,
            in2 => \_gnd_net_\,
            in3 => \N__21174\,
            lcout => \b2v_inst.un2_dir_mem_3_ac0_3\,
            ltout => \b2v_inst.un2_dir_mem_3_ac0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_3_RNO_0_5_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000101"
        )
    port map (
            in0 => \N__20295\,
            in1 => \N__20797\,
            in2 => \N__16250\,
            in3 => \N__18003\,
            lcout => \b2v_inst.un1_dir_mem_3_ns_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_1_RNO_1_6_LC_9_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000001110001"
        )
    port map (
            in0 => \N__21092\,
            in1 => \N__20115\,
            in2 => \N__18019\,
            in3 => \N__21176\,
            lcout => \b2v_inst.m7_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_0_rep2_RNI875S_LC_9_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21175\,
            in1 => \N__20093\,
            in2 => \N__20324\,
            in3 => \N__21091\,
            lcout => \b2v_inst.un8_dir_mem_3_c4\,
            ltout => \b2v_inst.un8_dir_mem_3_c4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_3_RNO_0_6_LC_9_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16556\,
            in3 => \N__20957\,
            lcout => \b2v_inst.un8_dir_mem_3_c6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_2_RNO_0_4_LC_9_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110001001101"
        )
    port map (
            in0 => \N__20123\,
            in1 => \N__20330\,
            in2 => \N__23077\,
            in3 => \N__21094\,
            lcout => OPEN,
            ltout => \b2v_inst.un2_indice_1_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_2_4_LC_9_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110011100011000"
        )
    port map (
            in0 => \N__20331\,
            in1 => \N__16725\,
            in2 => \N__16544\,
            in3 => \N__18029\,
            lcout => \b2v_inst.dir_mem_2Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22412\,
            ce => \N__16678\,
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_2_1_LC_9_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110011001"
        )
    port map (
            in0 => \N__23063\,
            in1 => \N__23202\,
            in2 => \_gnd_net_\,
            in3 => \N__16724\,
            lcout => \b2v_inst.dir_mem_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22412\,
            ce => \N__16678\,
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_2_2_LC_9_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001011011000"
        )
    port map (
            in0 => \N__16722\,
            in1 => \N__20124\,
            in2 => \N__17471\,
            in3 => \N__23064\,
            lcout => \b2v_inst.dir_mem_2Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22412\,
            ce => \N__16678\,
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_RNI6V1O2_7_LC_9_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010011"
        )
    port map (
            in0 => \N__19615\,
            in1 => \N__18299\,
            in2 => \N__20666\,
            in3 => \N__20932\,
            lcout => \b2v_inst.dir_mem_215_0\,
            ltout => \b2v_inst.dir_mem_215_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_2_0_LC_9_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010110100101"
        )
    port map (
            in0 => \N__23201\,
            in1 => \_gnd_net_\,
            in2 => \N__16496\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst.dir_mem_2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22412\,
            ce => \N__16678\,
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_2_5_LC_9_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100011110111000"
        )
    port map (
            in0 => \N__20664\,
            in1 => \N__16723\,
            in2 => \N__17930\,
            in3 => \N__20502\,
            lcout => \b2v_inst.dir_mem_2Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22412\,
            ce => \N__16678\,
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_SM_Main_ns_2_0__m13_LC_9_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21359\,
            in2 => \_gnd_net_\,
            in3 => \N__24020\,
            lcout => \b2v_inst1.N_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_RNIN0GU1_0_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17773\,
            in2 => \N__16625\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_10_10_0_\,
            carryout => \b2v_inst.un2_indice_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_RNO_4_1_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16616\,
            in2 => \N__17792\,
            in3 => \N__16610\,
            lcout => \b2v_inst.un2_indice_20_1\,
            ltout => OPEN,
            carryin => \b2v_inst.un2_indice_cry_0\,
            carryout => \b2v_inst.un2_indice_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_RNO_2_2_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16607\,
            in2 => \N__17794\,
            in3 => \N__16601\,
            lcout => \b2v_inst.un2_indice_20_2\,
            ltout => OPEN,
            carryin => \b2v_inst.un2_indice_cry_1\,
            carryout => \b2v_inst.un2_indice_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_RNO_2_3_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16598\,
            in2 => \N__17793\,
            in3 => \N__16592\,
            lcout => \b2v_inst.un2_indice_20_3\,
            ltout => OPEN,
            carryin => \b2v_inst.un2_indice_cry_2\,
            carryout => \b2v_inst.un2_indice_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_RNO_1_4_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17780\,
            in2 => \N__16745\,
            in3 => \N__16589\,
            lcout => \b2v_inst.un2_indice_20_4\,
            ltout => OPEN,
            carryin => \b2v_inst.un2_indice_cry_3\,
            carryout => \b2v_inst.un2_indice_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_RNO_2_5_LC_10_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17786\,
            in2 => \N__16841\,
            in3 => \N__16586\,
            lcout => \b2v_inst.un2_indice_20_5\,
            ltout => OPEN,
            carryin => \b2v_inst.un2_indice_cry_4\,
            carryout => \b2v_inst.un2_indice_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_RNO_1_6_LC_10_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17781\,
            in2 => \N__16583\,
            in3 => \N__16568\,
            lcout => \b2v_inst.un2_indice_20_6\,
            ltout => OPEN,
            carryin => \b2v_inst.un2_indice_cry_5\,
            carryout => \b2v_inst.un2_indice_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_RNO_3_7_LC_10_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111011010001"
        )
    port map (
            in0 => \N__20935\,
            in1 => \N__19740\,
            in2 => \N__19159\,
            in3 => \N__16775\,
            lcout => \b2v_inst.un2_indice_20_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_1_rep2_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__21134\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23166\,
            lcout => \b2v_inst.indice_1_repZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21964\,
            ce => \N__22951\,
            sr => \N__22906\
        );

    \b2v_inst.indice_0_rep2_RNIHJJG_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21133\,
            in2 => \_gnd_net_\,
            in3 => \N__21058\,
            lcout => \b2v_inst.un2_indice_21_s0_1\,
            ltout => \b2v_inst.un2_indice_21_s0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_RNO_2_1_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18766\,
            in2 => \N__16772\,
            in3 => \N__17399\,
            lcout => \b2v_inst.dir_mem_RNO_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_0_rep2_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1000111100001111"
        )
    port map (
            in0 => \N__19671\,
            in1 => \N__21005\,
            in2 => \N__21085\,
            in3 => \N__19613\,
            lcout => \b2v_inst.indice_0_repZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21964\,
            ce => \N__22951\,
            sr => \N__22906\
        );

    \b2v_inst.dir_mem_RNO_3_1_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100000"
        )
    port map (
            in0 => \N__17400\,
            in1 => \N__18767\,
            in2 => \N__16769\,
            in3 => \N__16760\,
            lcout => OPEN,
            ltout => \b2v_inst.dir_mem_RNO_3Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_RNO_0_1_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16754\,
            in2 => \N__16748\,
            in3 => \N__16803\,
            lcout => \b2v_inst.un2_indice_3_iv_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_0_LC_10_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1000000011111111"
        )
    port map (
            in0 => \N__21004\,
            in1 => \N__19672\,
            in2 => \N__19616\,
            in3 => \N__23167\,
            lcout => \b2v_inst.indiceZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21964\,
            ce => \N__22951\,
            sr => \N__22906\
        );

    \b2v_inst.dir_mem_RNIP73H1_4_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011000011"
        )
    port map (
            in0 => \N__19357\,
            in1 => \N__17769\,
            in2 => \N__17973\,
            in3 => \N__19724\,
            lcout => \b2v_inst.dir_mem_RNIP73H1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_4_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20822\,
            in2 => \_gnd_net_\,
            in3 => \N__17958\,
            lcout => \b2v_inst.indiceZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22280\,
            ce => \N__22950\,
            sr => \N__22912\
        );

    \b2v_inst.indice_5_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101010"
        )
    port map (
            in0 => \N__20407\,
            in1 => \N__20824\,
            in2 => \N__17974\,
            in3 => \N__21265\,
            lcout => \b2v_inst.indiceZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22280\,
            ce => \N__22950\,
            sr => \N__22912\
        );

    \b2v_inst.indice_4_rep1_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__20823\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21222\,
            lcout => \b2v_inst.indice_4_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22280\,
            ce => \N__22950\,
            sr => \N__22912\
        );

    \b2v_inst.dir_mem_RNIR93H1_5_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100000101101"
        )
    port map (
            in0 => \N__19725\,
            in1 => \N__19256\,
            in2 => \N__17791\,
            in3 => \N__20404\,
            lcout => \b2v_inst.dir_mem_RNIR93H1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_RNO_7_6_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__20405\,
            in1 => \N__17108\,
            in2 => \N__19519\,
            in3 => \N__21220\,
            lcout => \b2v_inst.g1_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_RNO_5_0_LC_10_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__21221\,
            in1 => \N__18986\,
            in2 => \N__17117\,
            in3 => \N__20406\,
            lcout => \b2v_inst.g0_2_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_RNO_0_5_LC_10_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16868\,
            in2 => \_gnd_net_\,
            in3 => \N__18764\,
            lcout => OPEN,
            ltout => \b2v_inst.N_411_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_5_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110111110101"
        )
    port map (
            in0 => \N__17303\,
            in1 => \N__16804\,
            in2 => \N__16787\,
            in3 => \N__16784\,
            lcout => \b2v_inst.dir_memZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21945\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_4_rep1_RNI93E71_LC_10_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__20277\,
            in1 => \N__21206\,
            in2 => \N__19517\,
            in3 => \N__21155\,
            lcout => \b2v_inst.un8_dir_mem_2_c4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_3_rep1_RNI4RFQ_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000001"
        )
    port map (
            in0 => \N__21157\,
            in1 => \N__21084\,
            in2 => \N__19518\,
            in3 => \N__17088\,
            lcout => \b2v_inst.un2_indice_21_s0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_RNO_3_5_LC_10_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011011111111"
        )
    port map (
            in0 => \N__20403\,
            in1 => \N__17962\,
            in2 => \N__16862\,
            in3 => \N__17380\,
            lcout => \b2v_inst.un2_indice_3_iv_0_a2_2_sx_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_2_rep1_RNIQKCO_LC_10_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000010001"
        )
    port map (
            in0 => \N__21156\,
            in1 => \N__21083\,
            in2 => \_gnd_net_\,
            in3 => \N__19504\,
            lcout => \b2v_inst.un2_indice_21_s0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_4_rep1_RNIP76I_0_LC_10_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__20402\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21204\,
            lcout => \b2v_inst.un2_indice_3_0_iv_0_a2_0_8_2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_fast_RNIDAJG_2_LC_10_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__21205\,
            in1 => \N__17087\,
            in2 => \_gnd_net_\,
            in3 => \N__18338\,
            lcout => \b2v_inst.indice_fast_RNIDAJGZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_3_rep1_RNI2RFQ_LC_10_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__17112\,
            in1 => \N__18389\,
            in2 => \N__19515\,
            in3 => \N__17873\,
            lcout => \b2v_inst.un2_indice_0_d0_c4_d\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_RNO_5_7_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20630\,
            in2 => \_gnd_net_\,
            in3 => \N__20441\,
            lcout => OPEN,
            ltout => \b2v_inst.un2_m1_e_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_RNO_2_7_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111100010000"
        )
    port map (
            in0 => \N__21225\,
            in1 => \N__16855\,
            in2 => \N__16844\,
            in3 => \N__20928\,
            lcout => \b2v_inst.dir_mem_RNO_2Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_0_rep1_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1101010101010101"
        )
    port map (
            in0 => \N__17875\,
            in1 => \N__21003\,
            in2 => \N__19614\,
            in3 => \N__19665\,
            lcout => \b2v_inst.indice_0_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22281\,
            ce => \N__22949\,
            sr => \N__22913\
        );

    \b2v_inst.dir_mem_RNO_4_4_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__17113\,
            in1 => \N__18390\,
            in2 => \N__19516\,
            in3 => \N__17874\,
            lcout => OPEN,
            ltout => \b2v_inst.dir_mem_RNO_4Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_RNO_2_4_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111111110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17390\,
            in2 => \N__17048\,
            in3 => \N__21224\,
            lcout => \b2v_inst.dir_mem_RNO_2Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_3_rep1_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__20113\,
            in1 => \N__23036\,
            in2 => \N__20333\,
            in3 => \N__23195\,
            lcout => \b2v_inst.indice_3_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22281\,
            ce => \N__22949\,
            sr => \N__22913\
        );

    \b2v_inst.indice_RNIA33N_1_LC_10_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__23037\,
            in1 => \N__20323\,
            in2 => \N__23215\,
            in3 => \N__20114\,
            lcout => \b2v_inst.indice_RNIA33NZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_3_RNIDN331_2_LC_10_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__17011\,
            in1 => \N__16957\,
            in2 => \N__16895\,
            in3 => \N__20094\,
            lcout => \b2v_inst.addr_ram_1_0_iv_i_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_2_LC_10_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101010"
        )
    port map (
            in0 => \N__20095\,
            in1 => \N__23174\,
            in2 => \N__23076\,
            in3 => \N__21251\,
            lcout => \b2v_inst.indiceZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21946\,
            ce => \N__22947\,
            sr => \N__22916\
        );

    \b2v_inst.indice_4_rep1_RNIQ9HI1_LC_10_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__20990\,
            in1 => \N__19603\,
            in2 => \_gnd_net_\,
            in3 => \N__19656\,
            lcout => \b2v_inst.un10_indice\,
            ltout => \b2v_inst.un10_indice_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_fast_2_LC_10_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000011000001100"
        )
    port map (
            in0 => \N__23058\,
            in1 => \N__18337\,
            in2 => \N__16871\,
            in3 => \N__23175\,
            lcout => \b2v_inst.indice_fastZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21946\,
            ce => \N__22947\,
            sr => \N__22916\
        );

    \b2v_inst.indice_fast_3_LC_10_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__23059\,
            in1 => \N__20106\,
            in2 => \N__20329\,
            in3 => \N__23176\,
            lcout => \b2v_inst.indice_fastZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21946\,
            ce => \N__22947\,
            sr => \N__22916\
        );

    \b2v_inst.indice_1_rep1_LC_10_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__23173\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18392\,
            lcout => \b2v_inst.indice_1_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21946\,
            ce => \N__22947\,
            sr => \N__22916\
        );

    \b2v_inst1.r_RX_Byte_RNO_0_2_LC_10_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__18090\,
            in1 => \N__18227\,
            in2 => \_gnd_net_\,
            in3 => \N__18193\,
            lcout => \b2v_inst1.r_RX_Bytece_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_Clk_Count_RNO_10_5_LC_10_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__23591\,
            in1 => \N__21467\,
            in2 => \N__23474\,
            in3 => \N__21563\,
            lcout => \b2v_inst1.g0_0_i_a6_3_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_Clk_Count_RNI9O3K3_6_LC_10_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__24018\,
            in1 => \N__23749\,
            in2 => \N__21354\,
            in3 => \N__23593\,
            lcout => \b2v_inst1.r_RX_Byte_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_Clk_Count_RNO_1_6_LC_10_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001100000101"
        )
    port map (
            in0 => \N__23592\,
            in1 => \N__23445\,
            in2 => \N__23756\,
            in3 => \N__24019\,
            lcout => \b2v_inst1.g0_7_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_RX_Byte_RNO_0_0_LC_10_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__18089\,
            in1 => \N__18226\,
            in2 => \_gnd_net_\,
            in3 => \N__18192\,
            lcout => \b2v_inst1.r_RX_Bytece_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_SM_Main_2_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__23989\,
            in1 => \N__23738\,
            in2 => \N__23623\,
            in3 => \N__21353\,
            lcout => \b2v_inst1.r_SM_MainZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22411\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_Clk_Count_RNO_6_4_LC_10_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__23910\,
            in1 => \N__23594\,
            in2 => \_gnd_net_\,
            in3 => \N__23988\,
            lcout => \b2v_inst1.g0_0_i_a6_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_2_RNO_2_6_LC_10_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__17114\,
            in1 => \N__21158\,
            in2 => \N__19520\,
            in3 => \N__21093\,
            lcout => \b2v_inst.un2_dir_mem_2_c4_d\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_Clk_Count_RNO_11_5_LC_10_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__23987\,
            in1 => \N__23603\,
            in2 => \N__23475\,
            in3 => \N__23911\,
            lcout => \b2v_inst1.g0_0_i_a6_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_Clk_Count_RNO_3_5_LC_10_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__19411\,
            in1 => \N__22694\,
            in2 => \N__23625\,
            in3 => \N__21725\,
            lcout => \b2v_inst1.N_11_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_Clk_Count_1_LC_10_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110011101110"
        )
    port map (
            in0 => \N__21395\,
            in1 => \N__17204\,
            in2 => \N__23496\,
            in3 => \N__18461\,
            lcout => \b2v_inst1.r_Clk_CountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22453\,
            ce => 'H',
            sr => \N__24082\
        );

    \b2v_inst1.r_Clk_Count_RNO_3_6_LC_10_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__23837\,
            in1 => \N__21456\,
            in2 => \N__21562\,
            in3 => \N__23918\,
            lcout => OPEN,
            ltout => \b2v_inst1.N_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_Clk_Count_RNO_0_6_LC_10_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111110001111"
        )
    port map (
            in0 => \N__21694\,
            in1 => \N__23919\,
            in2 => \N__17237\,
            in3 => \N__23343\,
            lcout => \b2v_inst1.N_11_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_Clk_Count_RNO_7_5_LC_10_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__19418\,
            in1 => \N__22690\,
            in2 => \_gnd_net_\,
            in3 => \N__21724\,
            lcout => \b2v_inst1.N_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_Clk_Count_RNI64771_1_LC_10_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__21455\,
            in1 => \N__21552\,
            in2 => \_gnd_net_\,
            in3 => \N__23836\,
            lcout => \b2v_inst1.N_9\,
            ltout => \b2v_inst1.N_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_Clk_Count_RNO_8_5_LC_10_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001010"
        )
    port map (
            in0 => \N__17234\,
            in1 => \N__23342\,
            in2 => \N__17228\,
            in3 => \N__21693\,
            lcout => OPEN,
            ltout => \b2v_inst1.N_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_Clk_Count_RNO_2_5_LC_10_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__18287\,
            in1 => \N__17225\,
            in2 => \N__17216\,
            in3 => \N__17213\,
            lcout => \b2v_inst1.g0_0_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_Clk_Count_RNO_2_1_LC_10_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__21734\,
            in1 => \N__23729\,
            in2 => \N__17198\,
            in3 => \N__23620\,
            lcout => \b2v_inst1.r_SM_Main_1_sqmuxa_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_Clk_Count_RNO_5_1_LC_10_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__19416\,
            in1 => \N__23316\,
            in2 => \N__22698\,
            in3 => \N__21689\,
            lcout => \b2v_inst1.g0_3_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_Clk_Count_RNO_6_5_LC_10_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__21690\,
            in1 => \N__23728\,
            in2 => \N__23341\,
            in3 => \N__23619\,
            lcout => OPEN,
            ltout => \b2v_inst1.g0_0_i_a6_2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_Clk_Count_RNO_1_5_LC_10_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101100"
        )
    port map (
            in0 => \N__17294\,
            in1 => \N__17288\,
            in2 => \N__17297\,
            in3 => \N__18449\,
            lcout => \b2v_inst1.g0_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_Clk_Count_RNO_5_5_LC_10_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010101010"
        )
    port map (
            in0 => \N__23915\,
            in1 => \N__23618\,
            in2 => \_gnd_net_\,
            in3 => \N__24003\,
            lcout => \b2v_inst1.g0_0_i_a6_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_Clk_Count_RNO_4_5_LC_10_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100010001"
        )
    port map (
            in0 => \N__23617\,
            in1 => \N__23705\,
            in2 => \N__23495\,
            in3 => \N__23916\,
            lcout => \b2v_inst1.N_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_RNO_0_4_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111101001100"
        )
    port map (
            in0 => \N__17535\,
            in1 => \N__17282\,
            in2 => \N__17429\,
            in3 => \N__18770\,
            lcout => OPEN,
            ltout => \b2v_inst.un2_indice_3_0_i_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_4_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000000010000"
        )
    port map (
            in0 => \N__18530\,
            in1 => \N__18771\,
            in2 => \N__17270\,
            in3 => \N__17267\,
            lcout => \b2v_inst.dir_memZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21874\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_RNO_1_2_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011010011110000"
        )
    port map (
            in0 => \N__19755\,
            in1 => \N__19808\,
            in2 => \N__19212\,
            in3 => \N__19890\,
            lcout => \b2v_inst.un2_indice_21_s1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_RNO_0_7_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010010101110"
        )
    port map (
            in0 => \N__18769\,
            in1 => \N__17411\,
            in2 => \N__17258\,
            in3 => \N__17246\,
            lcout => OPEN,
            ltout => \b2v_inst.un2_indice_3_0_iv_0_0_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_7_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001101"
        )
    port map (
            in0 => \N__17537\,
            in1 => \N__19091\,
            in2 => \N__17240\,
            in3 => \N__18529\,
            lcout => \b2v_inst.dir_memZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21874\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_RNO_0_2_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010010101110"
        )
    port map (
            in0 => \N__18768\,
            in1 => \N__17410\,
            in2 => \N__17467\,
            in3 => \N__17444\,
            lcout => OPEN,
            ltout => \b2v_inst.un2_indice_3_0_iv_0_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_2_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001101"
        )
    port map (
            in0 => \N__17536\,
            in1 => \N__17438\,
            in2 => \N__17432\,
            in3 => \N__18528\,
            lcout => \b2v_inst.dir_memZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21874\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_RNO_3_4_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101100110"
        )
    port map (
            in0 => \N__17309\,
            in1 => \N__19362\,
            in2 => \_gnd_net_\,
            in3 => \N__19754\,
            lcout => \b2v_inst.dir_mem_RNO_3Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_RNO_1_3_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__19315\,
            in1 => \N__17417\,
            in2 => \_gnd_net_\,
            in3 => \N__19199\,
            lcout => \b2v_inst.un2_indice_21_s1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_RNO_3_3_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000001000000"
        )
    port map (
            in0 => \N__19760\,
            in1 => \N__19805\,
            in2 => \N__19889\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst.un2_indice_0_d1_c2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_RNO_0_3_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001011001110"
        )
    port map (
            in0 => \N__17409\,
            in1 => \N__18772\,
            in2 => \N__17342\,
            in3 => \N__17327\,
            lcout => OPEN,
            ltout => \b2v_inst.un2_indice_3_0_iv_0_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_3_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010000000101"
        )
    port map (
            in0 => \N__18527\,
            in1 => \N__17318\,
            in2 => \N__17312\,
            in3 => \N__17534\,
            lcout => \b2v_inst.dir_memZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22081\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_RNO_5_4_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__19804\,
            in1 => \N__19198\,
            in2 => \N__19321\,
            in3 => \N__19876\,
            lcout => \b2v_inst.dir_mem_RNO_5Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_RNO_1_5_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000100010101"
        )
    port map (
            in0 => \N__17823\,
            in1 => \N__17525\,
            in2 => \N__19385\,
            in3 => \N__19255\,
            lcout => \b2v_inst.un2_indice_3_iv_0_1_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_1_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__17526\,
            in1 => \N__17824\,
            in2 => \N__19685\,
            in3 => \N__17804\,
            lcout => \b2v_inst.dir_memZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22081\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_RNO_4_0_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011000111100"
        )
    port map (
            in0 => \N__19894\,
            in1 => \N__17798\,
            in2 => \N__21095\,
            in3 => \N__19756\,
            lcout => OPEN,
            ltout => \b2v_inst.un2_indice_20_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_RNO_1_0_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100000000"
        )
    port map (
            in0 => \N__18931\,
            in1 => \N__17699\,
            in2 => \N__17588\,
            in3 => \N__18763\,
            lcout => \b2v_inst.N_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNIN365_15_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18932\,
            in2 => \_gnd_net_\,
            in3 => \N__18990\,
            lcout => \b2v_inst.N_228\,
            ltout => \b2v_inst.N_228_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_17_rep1_RNIVTJP1_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010011111100"
        )
    port map (
            in0 => \N__17573\,
            in1 => \N__19075\,
            in2 => \N__17552\,
            in3 => \N__17549\,
            lcout => \b2v_inst.N_234\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_0_rep1_RNIO9HI1_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__19655\,
            in1 => \N__17482\,
            in2 => \_gnd_net_\,
            in3 => \N__17506\,
            lcout => OPEN,
            ltout => \b2v_inst.N_383_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_17_rep1_RNIN75C3_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000010000"
        )
    port map (
            in0 => \N__19071\,
            in1 => \N__17495\,
            in2 => \N__17489\,
            in3 => \N__18762\,
            lcout => \b2v_inst.state_17_rep1_RNIN75CZ0Z3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_0_rep1_RNIEF5S_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__20867\,
            in1 => \N__17868\,
            in2 => \N__18393\,
            in3 => \N__20557\,
            lcout => \b2v_inst.un2_indice_3_0_iv_0_a2_0_8_3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_fast_RNIHI54_3_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20710\,
            in2 => \_gnd_net_\,
            in3 => \N__18330\,
            lcout => \b2v_inst.un10_indice_2\,
            ltout => \b2v_inst.un10_indice_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_fast_RNI7BF71_4_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111110001100"
        )
    port map (
            in0 => \N__20756\,
            in1 => \N__17834\,
            in2 => \N__18056\,
            in3 => \N__18053\,
            lcout => \b2v_inst.dir_mem_115lto6_1\,
            ltout => \b2v_inst.dir_mem_115lto6_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_1_RNO_0_7_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18047\,
            in3 => \N__20192\,
            lcout => OPEN,
            ltout => \b2v_inst.un1_dir_mem_1_mb_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_1_7_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101001010100"
        )
    port map (
            in0 => \N__19588\,
            in1 => \N__20180\,
            in2 => \N__18044\,
            in3 => \N__20868\,
            lcout => \b2v_inst.dir_mem_1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22082\,
            ce => \N__19933\,
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_2_RNO_0_5_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__18018\,
            in1 => \N__20096\,
            in2 => \N__20027\,
            in3 => \N__20325\,
            lcout => \b2v_inst.un2_dir_mem_2_c5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_1_RNO_2_4_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21172\,
            in2 => \_gnd_net_\,
            in3 => \N__21090\,
            lcout => OPEN,
            ltout => \b2v_inst.N_4_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_1_RNO_0_4_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111111111111"
        )
    port map (
            in0 => \N__20898\,
            in1 => \N__20097\,
            in2 => \N__17915\,
            in3 => \N__20326\,
            lcout => \b2v_inst.N_8_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_0_rep1_RNIATP21_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010011"
        )
    port map (
            in0 => \N__17870\,
            in1 => \N__20897\,
            in2 => \N__18394\,
            in3 => \N__21223\,
            lcout => OPEN,
            ltout => \b2v_inst.dir_mem_315lto8_a0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_fast_RNIRFV61_3_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20712\,
            in2 => \N__17903\,
            in3 => \N__18332\,
            lcout => \b2v_inst.indice_fast_RNIRFV61Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_0_rep1_RNIFJJG_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__17869\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18381\,
            lcout => \b2v_inst.indice_0_rep1_RNIFJJGZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_fast_RNIJ9NJ_3_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000001"
        )
    port map (
            in0 => \N__18382\,
            in1 => \N__20711\,
            in2 => \N__20763\,
            in3 => \N__18331\,
            lcout => OPEN,
            ltout => \b2v_inst.dir_mem_215lt6_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_RNIG39V_6_LC_11_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20453\,
            in2 => \N__18302\,
            in3 => \N__20561\,
            lcout => \b2v_inst.dir_mem_215lt8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_Clk_Count_RNO_9_5_LC_11_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__21657\,
            in1 => \N__24016\,
            in2 => \N__23344\,
            in3 => \N__23832\,
            lcout => \b2v_inst1.g0_0_i_a6_3_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_Clk_Count_RNO_0_3_LC_11_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__21560\,
            in1 => \_gnd_net_\,
            in2 => \N__21476\,
            in3 => \N__23833\,
            lcout => \b2v_inst1.un1_r_Clk_Count_ac0_3_out\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_SM_Main_ns_2_0__m16_e_LC_11_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__18224\,
            in1 => \N__18088\,
            in2 => \_gnd_net_\,
            in3 => \N__18186\,
            lcout => \b2v_inst1.r_rx_byteZ0Z_7\,
            ltout => \b2v_inst1.r_rx_byteZ0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_SM_Main_ns_2_0__m17_LC_11_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100011001100"
        )
    port map (
            in0 => \N__21351\,
            in1 => \N__23741\,
            in2 => \N__18263\,
            in3 => \N__24017\,
            lcout => \b2v_inst1.N_32_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_Clk_Count_RNO_4_6_LC_11_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111111111"
        )
    port map (
            in0 => \N__20339\,
            in1 => \N__21463\,
            in2 => \_gnd_net_\,
            in3 => \N__21559\,
            lcout => \b2v_inst1.N_10_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_Bit_Index_2_LC_11_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__21311\,
            in1 => \N__18225\,
            in2 => \N__18194\,
            in3 => \N__18103\,
            lcout => \b2v_inst1.r_Bit_IndexZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22455\,
            ce => 'H',
            sr => \N__24081\
        );

    \b2v_inst1.r_Bit_Index_1_LC_11_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__18102\,
            in1 => \N__18187\,
            in2 => \_gnd_net_\,
            in3 => \N__21310\,
            lcout => \b2v_inst1.r_Bit_IndexZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22455\,
            ce => 'H',
            sr => \N__24081\
        );

    \b2v_inst1.r_Clk_Count_RNO_0_5_LC_11_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111101001111"
        )
    port map (
            in0 => \N__21661\,
            in1 => \N__18455\,
            in2 => \N__23351\,
            in3 => \N__18448\,
            lcout => \b2v_inst1.N_14_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_SM_Main_ns_2_0__m22_ns_1_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100001100"
        )
    port map (
            in0 => \N__23992\,
            in1 => \N__23727\,
            in2 => \N__22709\,
            in3 => \N__23589\,
            lcout => \b2v_inst1.m22_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_Clk_Count_RNO_9_4_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001011111010"
        )
    port map (
            in0 => \N__23588\,
            in1 => \N__23903\,
            in2 => \N__23748\,
            in3 => \N__23991\,
            lcout => \b2v_inst1.N_9_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_SM_Main_ns_2_0__m2_0_LC_11_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21439\,
            in2 => \_gnd_net_\,
            in3 => \N__21527\,
            lcout => \b2v_inst1.un1_r_Clk_Count_ac0_1_out\,
            ltout => \b2v_inst1.un1_r_Clk_Count_ac0_1_out_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_SM_Main_ns_2_0__m6_LC_11_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__21660\,
            in1 => \N__19415\,
            in2 => \N__18437\,
            in3 => \N__23315\,
            lcout => \b2v_inst1.N_29_mux\,
            ltout => \b2v_inst1.N_29_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_SM_Main_1_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111010100000"
        )
    port map (
            in0 => \N__18434\,
            in1 => \N__21352\,
            in2 => \N__18428\,
            in3 => \N__23590\,
            lcout => \b2v_inst1.r_SM_MainZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22561\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_SM_Main_ns_2_0__m10_LC_11_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21528\,
            in1 => \N__23902\,
            in2 => \N__21462\,
            in3 => \N__23820\,
            lcout => OPEN,
            ltout => \b2v_inst1.N_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_SM_Main_ns_2_0__m12_LC_11_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101000111"
        )
    port map (
            in0 => \N__23904\,
            in1 => \N__23347\,
            in2 => \N__18425\,
            in3 => \N__21659\,
            lcout => \b2v_inst1.N_28_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_Clk_Count_5_LC_11_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100000001"
        )
    port map (
            in0 => \N__18422\,
            in1 => \N__18413\,
            in2 => \N__18407\,
            in3 => \N__23901\,
            lcout => \b2v_inst1.r_Clk_CountZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22550\,
            ce => 'H',
            sr => \N__24093\
        );

    \b2v_inst1.r_SM_Main_ns_2_0__m6_2_LC_11_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__23984\,
            in1 => \N__23900\,
            in2 => \_gnd_net_\,
            in3 => \N__23809\,
            lcout => \b2v_inst1.m6_2\,
            ltout => \b2v_inst1.m6_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_SM_Main_ns_2_0__g0_6_LC_11_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__21656\,
            in1 => \N__23285\,
            in2 => \N__18512\,
            in3 => \N__21723\,
            lcout => \b2v_inst1.N_29_mux_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_Clk_Count_RNO_2_6_LC_11_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100100000"
        )
    port map (
            in0 => \N__23985\,
            in1 => \N__23612\,
            in2 => \N__23742\,
            in3 => \N__18509\,
            lcout => OPEN,
            ltout => \b2v_inst1.g0_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_Clk_Count_6_LC_11_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001100001011"
        )
    port map (
            in0 => \N__23613\,
            in1 => \N__18500\,
            in2 => \N__18488\,
            in3 => \N__18485\,
            lcout => \b2v_inst1.r_Clk_CountZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22550\,
            ce => 'H',
            sr => \N__24093\
        );

    \b2v_inst1.r_SM_Main_ns_2_0__m9_LC_11_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__23708\,
            in1 => \_gnd_net_\,
            in2 => \N__22699\,
            in3 => \N__21767\,
            lcout => OPEN,
            ltout => \b2v_inst1.N_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_SM_Main_0_LC_11_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000000101"
        )
    port map (
            in0 => \N__23482\,
            in1 => \N__18476\,
            in2 => \N__18467\,
            in3 => \N__23622\,
            lcout => \b2v_inst1.r_SM_MainZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22510\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_Clk_Count_RNIAI9K1_1_LC_11_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__21443\,
            in1 => \N__21532\,
            in2 => \N__21695\,
            in3 => \N__23821\,
            lcout => \b2v_inst1.N_11_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_Clk_Count_RNO_3_1_LC_11_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__21533\,
            in1 => \N__23762\,
            in2 => \N__21692\,
            in3 => \N__21444\,
            lcout => OPEN,
            ltout => \b2v_inst1.g2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_Clk_Count_RNO_0_1_LC_11_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110011"
        )
    port map (
            in0 => \N__21578\,
            in1 => \N__23707\,
            in2 => \N__18464\,
            in3 => \N__23621\,
            lcout => \b2v_inst1.g2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_Clk_Count_RNO_0_4_LC_11_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__22679\,
            in1 => \N__19417\,
            in2 => \_gnd_net_\,
            in3 => \N__21733\,
            lcout => \b2v_inst1.N_7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_RNO_4_5_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__19301\,
            in1 => \N__19200\,
            in2 => \N__19331\,
            in3 => \N__19757\,
            lcout => \b2v_inst.un2_indice_0_d1_c5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_RNIJMO11_4_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__19361\,
            in1 => \N__19806\,
            in2 => \_gnd_net_\,
            in3 => \N__19874\,
            lcout => \b2v_inst.un2_indice_0_d1_ac0_7_s_0_0\,
            ltout => \b2v_inst.un2_indice_0_d1_ac0_7_s_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_RNO_4_7_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__19302\,
            in1 => \N__19265\,
            in2 => \N__19220\,
            in3 => \N__19201\,
            lcout => OPEN,
            ltout => \b2v_inst.un2_indice_0_d1_ac0_9_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_RNO_1_7_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001110011001100"
        )
    port map (
            in0 => \N__19759\,
            in1 => \N__19149\,
            in2 => \N__19130\,
            in3 => \N__19126\,
            lcout => \b2v_inst.un2_indice_21_s1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNIVTJP1_15_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__19081\,
            in1 => \N__18997\,
            in2 => \N__18940\,
            in3 => \N__18765\,
            lcout => OPEN,
            ltout => \b2v_inst.N_384_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.state_RNIM5P55_15_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18552\,
            in2 => \N__18539\,
            in3 => \N__18536\,
            lcout => \b2v_inst.un2_indice_3_0_iv_0_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_RNO_1_1_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001100110"
        )
    port map (
            in0 => \N__19875\,
            in1 => \N__19807\,
            in2 => \_gnd_net_\,
            in3 => \N__19758\,
            lcout => \b2v_inst.un2_indice_21_s1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_fast_0_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1011001100110011"
        )
    port map (
            in0 => \N__19587\,
            in1 => \N__19550\,
            in2 => \N__21002\,
            in3 => \N__19666\,
            lcout => \b2v_inst.indice_fastZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22102\,
            ce => \N__22948\,
            sr => \N__22917\
        );

    \b2v_inst.indice_RNITPHB_6_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20617\,
            in2 => \_gnd_net_\,
            in3 => \N__20476\,
            lcout => \b2v_inst.CO1\,
            ltout => \b2v_inst.CO1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_2_rep1_RNI6ULR_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__19467\,
            in1 => \N__20685\,
            in2 => \N__19556\,
            in3 => \N__20019\,
            lcout => \b2v_inst.un8_dir_mem_1_c7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_fast_RNIDE54_0_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__19549\,
            in1 => \_gnd_net_\,
            in2 => \N__19538\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst.un2_dir_mem_2_c2\,
            ltout => \b2v_inst.un2_dir_mem_2_c2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_1_RNO_0_5_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__20477\,
            in1 => \N__19472\,
            in2 => \N__19553\,
            in3 => \N__20686\,
            lcout => \b2v_inst.dir_mem_1_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_fast_RNIF91E_0_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011111111111"
        )
    port map (
            in0 => \N__19548\,
            in1 => \N__19466\,
            in2 => \N__19537\,
            in3 => \N__20723\,
            lcout => \b2v_inst.indice_fast_RNIF91EZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_fast_1_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23206\,
            in2 => \_gnd_net_\,
            in3 => \N__19536\,
            lcout => \b2v_inst.indice_fastZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22102\,
            ce => \N__22948\,
            sr => \N__22917\
        );

    \b2v_inst.indice_2_rep1_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001001100100000"
        )
    port map (
            in0 => \N__23021\,
            in1 => \N__21266\,
            in2 => \N__23217\,
            in3 => \N__19468\,
            lcout => \b2v_inst.indice_2_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22102\,
            ce => \N__22948\,
            sr => \N__22917\
        );

    \b2v_inst.dir_mem_1_RNO_0_3_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011011001100"
        )
    port map (
            in0 => \N__23022\,
            in1 => \N__20327\,
            in2 => \N__23216\,
            in3 => \N__20141\,
            lcout => OPEN,
            ltout => \b2v_inst.dir_mem_1_RNO_0Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_1_3_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__20328\,
            in1 => \_gnd_net_\,
            in2 => \N__20213\,
            in3 => \N__19963\,
            lcout => \b2v_inst.dir_mem_1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22388\,
            ce => \N__19934\,
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_fast_RNI6ULR_4_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001110111111"
        )
    port map (
            in0 => \N__20198\,
            in1 => \N__20579\,
            in2 => \N__20764\,
            in3 => \N__20484\,
            lcout => \b2v_inst.dir_mem_115lto8_1\,
            ltout => \b2v_inst.dir_mem_115lto8_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_RNI36K43_7_LC_12_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110001"
        )
    port map (
            in0 => \N__20186\,
            in1 => \N__20179\,
            in2 => \N__20168\,
            in3 => \N__20927\,
            lcout => \b2v_inst.dir_mem_115_0\,
            ltout => \b2v_inst.dir_mem_115_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_1_0_LC_12_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__23199\,
            in1 => \_gnd_net_\,
            in2 => \N__20165\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst.dir_mem_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22388\,
            ce => \N__19934\,
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_1_2_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__20142\,
            in1 => \N__20020\,
            in2 => \_gnd_net_\,
            in3 => \N__19962\,
            lcout => \b2v_inst.dir_mem_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22388\,
            ce => \N__19934\,
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_1_5_LC_12_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__19964\,
            in1 => \N__19985\,
            in2 => \_gnd_net_\,
            in3 => \N__20485\,
            lcout => \b2v_inst.dir_mem_1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22388\,
            ce => \N__19934\,
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_1_1_LC_12_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100111001100"
        )
    port map (
            in0 => \N__23200\,
            in1 => \N__23023\,
            in2 => \_gnd_net_\,
            in3 => \N__19961\,
            lcout => \b2v_inst.dir_mem_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22388\,
            ce => \N__19934\,
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_4_rep1_RNIP76I_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21232\,
            in2 => \_gnd_net_\,
            in3 => \N__20482\,
            lcout => \b2v_inst.un8_dir_mem_3_ac0_9_0\,
            ltout => \b2v_inst.un8_dir_mem_3_ac0_9_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_6_LC_12_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101010"
        )
    port map (
            in0 => \N__20577\,
            in1 => \N__20826\,
            in2 => \N__21269\,
            in3 => \N__21261\,
            lcout => \b2v_inst.indiceZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21884\,
            ce => \N__22946\,
            sr => \N__22920\
        );

    \b2v_inst.indice_4_rep1_RNICTP21_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__21233\,
            in1 => \N__21173\,
            in2 => \N__20899\,
            in3 => \N__21086\,
            lcout => \b2v_inst.un10_indice_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_7_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__20578\,
            in1 => \N__20872\,
            in2 => \N__20953\,
            in3 => \N__20827\,
            lcout => \b2v_inst.indiceZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21884\,
            ce => \N__22946\,
            sr => \N__22920\
        );

    \b2v_inst.indice_fast_4_LC_12_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__20755\,
            in1 => \_gnd_net_\,
            in2 => \N__20831\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst.indice_fastZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21884\,
            ce => \N__22946\,
            sr => \N__22920\
        );

    \b2v_inst.indice_fast_RNIJK54_3_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20754\,
            in2 => \_gnd_net_\,
            in3 => \N__20722\,
            lcout => \b2v_inst.un8_dir_mem_1_ac0_7_out\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.dir_mem_2_RNO_1_6_LC_12_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20665\,
            in1 => \N__20576\,
            in2 => \_gnd_net_\,
            in3 => \N__20483\,
            lcout => \b2v_inst.dir_mem_2_RNO_1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_Clk_Count_RNO_5_6_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__21658\,
            in1 => \N__23921\,
            in2 => \N__23346\,
            in3 => \N__23835\,
            lcout => \b2v_inst1.g0_i_o5_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_SM_Main_ns_2_0__g0_1_4_LC_12_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__24014\,
            in1 => \N__23920\,
            in2 => \N__23345\,
            in3 => \N__23834\,
            lcout => OPEN,
            ltout => \b2v_inst1.g0_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_SM_Main_ns_2_0__g0_0_LC_12_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__21662\,
            in1 => \N__21479\,
            in2 => \N__21362\,
            in3 => \N__21561\,
            lcout => \b2v_inst1.N_29_mux_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_SM_Main_RNIAP3K3_2_LC_12_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__23497\,
            in1 => \N__23739\,
            in2 => \N__21355\,
            in3 => \N__24015\,
            lcout => \b2v_inst1.un1_r_SM_Main_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_SM_Main_ns_2_0__g0_1_0_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__21477\,
            in1 => \N__21542\,
            in2 => \N__21666\,
            in3 => \N__23831\,
            lcout => OPEN,
            ltout => \b2v_inst1.g0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_SM_Main_ns_2_0__g0_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110000000000"
        )
    port map (
            in0 => \N__23314\,
            in1 => \N__24005\,
            in2 => \N__21299\,
            in3 => \N__23913\,
            lcout => OPEN,
            ltout => \b2v_inst1.N_14_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_SM_Main_RNIVAI26_0_LC_12_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011110101"
        )
    port map (
            in0 => \N__23599\,
            in1 => \N__21296\,
            in2 => \N__21290\,
            in3 => \N__23740\,
            lcout => \b2v_inst1.un1_r_SM_Main_1_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_Clk_Count_RNO_8_4_LC_12_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__21543\,
            in1 => \N__23598\,
            in2 => \N__23484\,
            in3 => \N__21478\,
            lcout => OPEN,
            ltout => \b2v_inst1.g0_0_i_a6_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_Clk_Count_RNO_3_4_LC_12_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__23912\,
            in1 => \N__21284\,
            in2 => \N__21287\,
            in3 => \N__23830\,
            lcout => \b2v_inst1.g0_0_i_a6_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_Clk_Count_RNO_7_4_LC_12_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21639\,
            in2 => \_gnd_net_\,
            in3 => \N__24004\,
            lcout => \b2v_inst1.g0_0_i_a6_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_Clk_Count_3_LC_12_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001101000010010"
        )
    port map (
            in0 => \N__21643\,
            in1 => \N__21747\,
            in2 => \N__21278\,
            in3 => \N__23455\,
            lcout => \b2v_inst1.r_Clk_CountZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22251\,
            ce => 'H',
            sr => \N__24094\
        );

    \b2v_inst1.r_Clk_Count_RNO_0_0_LC_12_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__23704\,
            in1 => \N__21766\,
            in2 => \N__22689\,
            in3 => \N__23608\,
            lcout => OPEN,
            ltout => \b2v_inst1.r_SM_Main_1_sqmuxa_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_Clk_Count_0_LC_12_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100111110001"
        )
    port map (
            in0 => \N__21531\,
            in1 => \N__21748\,
            in2 => \N__21752\,
            in3 => \N__23490\,
            lcout => \b2v_inst1.r_Clk_CountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22461\,
            ce => 'H',
            sr => \N__24092\
        );

    \b2v_inst1.r_Clk_Count_2_LC_12_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001000110100010"
        )
    port map (
            in0 => \N__23823\,
            in1 => \N__21749\,
            in2 => \N__23498\,
            in3 => \N__21732\,
            lcout => \b2v_inst1.r_Clk_CountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22461\,
            ce => 'H',
            sr => \N__24092\
        );

    \b2v_inst1.r_SM_Main_ns_2_0__g0_3_1_LC_12_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__21453\,
            in1 => \N__21529\,
            in2 => \N__21691\,
            in3 => \N__23822\,
            lcout => OPEN,
            ltout => \b2v_inst1.g0_3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_SM_Main_ns_2_0__g0_3_LC_12_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110000000000"
        )
    port map (
            in0 => \N__23313\,
            in1 => \N__23990\,
            in2 => \N__21581\,
            in3 => \N__23917\,
            lcout => \b2v_inst1.N_14_0_0\,
            ltout => \b2v_inst1.N_14_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_Clk_Count_RNO_4_1_LC_12_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000101110"
        )
    port map (
            in0 => \N__23703\,
            in1 => \N__23607\,
            in2 => \N__21572\,
            in3 => \N__21569\,
            lcout => OPEN,
            ltout => \b2v_inst1.g3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_Clk_Count_RNO_1_1_LC_12_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__21530\,
            in1 => \_gnd_net_\,
            in2 => \N__21482\,
            in3 => \N__21454\,
            lcout => \b2v_inst1.g3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_Clk_Count_RNO_5_4_LC_12_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__23365\,
            in1 => \N__21386\,
            in2 => \_gnd_net_\,
            in3 => \N__23294\,
            lcout => OPEN,
            ltout => \b2v_inst1.N_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_Clk_Count_RNO_2_4_LC_12_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111110000"
        )
    port map (
            in0 => \N__23295\,
            in1 => \N__23489\,
            in2 => \N__21377\,
            in3 => \N__21374\,
            lcout => OPEN,
            ltout => \b2v_inst1.g0_0_i_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_Clk_Count_4_LC_12_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100000011"
        )
    port map (
            in0 => \N__24113\,
            in1 => \N__23225\,
            in2 => \N__24104\,
            in3 => \N__24101\,
            lcout => \b2v_inst1.r_Clk_CountZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21890\,
            ce => 'H',
            sr => \N__24095\
        );

    \b2v_inst1.r_Clk_Count_RNO_6_1_LC_12_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__23986\,
            in1 => \N__23914\,
            in2 => \N__23320\,
            in3 => \N__23829\,
            lcout => \b2v_inst1.g2_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_Clk_Count_RNO_4_4_LC_12_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23706\,
            in2 => \_gnd_net_\,
            in3 => \N__23624\,
            lcout => OPEN,
            ltout => \b2v_inst1.g0_0_i_a6_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_Clk_Count_RNO_1_4_LC_12_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011111100"
        )
    port map (
            in0 => \N__23488\,
            in1 => \N__23366\,
            in2 => \N__23354\,
            in3 => \N__23301\,
            lcout => \b2v_inst1.g0_0_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst.indice_1_LC_13_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23218\,
            in2 => \_gnd_net_\,
            in3 => \N__22996\,
            lcout => \b2v_inst.indiceZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22500\,
            ce => \N__22945\,
            sr => \N__22922\
        );

    \b2v_inst1.r_RX_Data_R_LC_13_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22772\,
            lcout => \b2v_inst1.r_RX_Data_RZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22252\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst1.r_RX_Data_LC_13_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22757\,
            lcout => \b2v_inst1.r_RX_DataZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22252\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
