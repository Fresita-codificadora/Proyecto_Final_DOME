// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Oct 31 2024 19:51:40

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "anda_plis_2" view "INTERFACE"

module anda_plis_2 (
    leds,
    swit,
    uart_tx_o,
    uart_rx_i,
    clk,
    reset);

    output [13:0] leds;
    input [10:0] swit;
    output uart_tx_o;
    input uart_rx_i;
    input clk;
    input reset;

    wire N__39656;
    wire N__39655;
    wire N__39654;
    wire N__39645;
    wire N__39644;
    wire N__39643;
    wire N__39636;
    wire N__39635;
    wire N__39634;
    wire N__39627;
    wire N__39626;
    wire N__39625;
    wire N__39618;
    wire N__39617;
    wire N__39616;
    wire N__39609;
    wire N__39608;
    wire N__39607;
    wire N__39600;
    wire N__39599;
    wire N__39598;
    wire N__39591;
    wire N__39590;
    wire N__39589;
    wire N__39582;
    wire N__39581;
    wire N__39580;
    wire N__39573;
    wire N__39572;
    wire N__39571;
    wire N__39564;
    wire N__39563;
    wire N__39562;
    wire N__39555;
    wire N__39554;
    wire N__39553;
    wire N__39546;
    wire N__39545;
    wire N__39544;
    wire N__39537;
    wire N__39536;
    wire N__39535;
    wire N__39528;
    wire N__39527;
    wire N__39526;
    wire N__39519;
    wire N__39518;
    wire N__39517;
    wire N__39510;
    wire N__39509;
    wire N__39508;
    wire N__39501;
    wire N__39500;
    wire N__39499;
    wire N__39492;
    wire N__39491;
    wire N__39490;
    wire N__39483;
    wire N__39482;
    wire N__39481;
    wire N__39474;
    wire N__39473;
    wire N__39472;
    wire N__39465;
    wire N__39464;
    wire N__39463;
    wire N__39456;
    wire N__39455;
    wire N__39454;
    wire N__39447;
    wire N__39446;
    wire N__39445;
    wire N__39438;
    wire N__39437;
    wire N__39436;
    wire N__39429;
    wire N__39428;
    wire N__39427;
    wire N__39420;
    wire N__39419;
    wire N__39418;
    wire N__39411;
    wire N__39410;
    wire N__39409;
    wire N__39402;
    wire N__39401;
    wire N__39400;
    wire N__39383;
    wire N__39380;
    wire N__39377;
    wire N__39376;
    wire N__39373;
    wire N__39370;
    wire N__39369;
    wire N__39366;
    wire N__39363;
    wire N__39360;
    wire N__39359;
    wire N__39356;
    wire N__39351;
    wire N__39350;
    wire N__39349;
    wire N__39346;
    wire N__39343;
    wire N__39340;
    wire N__39337;
    wire N__39334;
    wire N__39323;
    wire N__39322;
    wire N__39319;
    wire N__39318;
    wire N__39317;
    wire N__39316;
    wire N__39313;
    wire N__39310;
    wire N__39307;
    wire N__39306;
    wire N__39305;
    wire N__39304;
    wire N__39303;
    wire N__39300;
    wire N__39297;
    wire N__39294;
    wire N__39289;
    wire N__39286;
    wire N__39283;
    wire N__39280;
    wire N__39277;
    wire N__39274;
    wire N__39273;
    wire N__39270;
    wire N__39267;
    wire N__39264;
    wire N__39261;
    wire N__39258;
    wire N__39255;
    wire N__39252;
    wire N__39249;
    wire N__39246;
    wire N__39243;
    wire N__39242;
    wire N__39237;
    wire N__39228;
    wire N__39227;
    wire N__39226;
    wire N__39223;
    wire N__39220;
    wire N__39217;
    wire N__39214;
    wire N__39209;
    wire N__39204;
    wire N__39199;
    wire N__39188;
    wire N__39187;
    wire N__39184;
    wire N__39181;
    wire N__39178;
    wire N__39175;
    wire N__39172;
    wire N__39169;
    wire N__39166;
    wire N__39163;
    wire N__39160;
    wire N__39157;
    wire N__39154;
    wire N__39151;
    wire N__39146;
    wire N__39143;
    wire N__39140;
    wire N__39139;
    wire N__39138;
    wire N__39135;
    wire N__39132;
    wire N__39129;
    wire N__39124;
    wire N__39123;
    wire N__39122;
    wire N__39119;
    wire N__39116;
    wire N__39113;
    wire N__39110;
    wire N__39101;
    wire N__39100;
    wire N__39097;
    wire N__39094;
    wire N__39091;
    wire N__39088;
    wire N__39085;
    wire N__39082;
    wire N__39081;
    wire N__39080;
    wire N__39079;
    wire N__39076;
    wire N__39073;
    wire N__39070;
    wire N__39069;
    wire N__39068;
    wire N__39065;
    wire N__39062;
    wire N__39059;
    wire N__39058;
    wire N__39053;
    wire N__39050;
    wire N__39049;
    wire N__39046;
    wire N__39041;
    wire N__39038;
    wire N__39035;
    wire N__39034;
    wire N__39031;
    wire N__39028;
    wire N__39027;
    wire N__39026;
    wire N__39023;
    wire N__39018;
    wire N__39013;
    wire N__39010;
    wire N__39007;
    wire N__39004;
    wire N__39001;
    wire N__38998;
    wire N__38995;
    wire N__38992;
    wire N__38987;
    wire N__38980;
    wire N__38969;
    wire N__38968;
    wire N__38965;
    wire N__38962;
    wire N__38959;
    wire N__38956;
    wire N__38953;
    wire N__38950;
    wire N__38947;
    wire N__38944;
    wire N__38941;
    wire N__38938;
    wire N__38935;
    wire N__38932;
    wire N__38927;
    wire N__38924;
    wire N__38921;
    wire N__38918;
    wire N__38917;
    wire N__38914;
    wire N__38911;
    wire N__38910;
    wire N__38909;
    wire N__38906;
    wire N__38905;
    wire N__38902;
    wire N__38899;
    wire N__38896;
    wire N__38893;
    wire N__38890;
    wire N__38887;
    wire N__38884;
    wire N__38881;
    wire N__38870;
    wire N__38867;
    wire N__38866;
    wire N__38863;
    wire N__38862;
    wire N__38861;
    wire N__38860;
    wire N__38857;
    wire N__38854;
    wire N__38851;
    wire N__38848;
    wire N__38847;
    wire N__38844;
    wire N__38843;
    wire N__38840;
    wire N__38837;
    wire N__38836;
    wire N__38833;
    wire N__38830;
    wire N__38829;
    wire N__38828;
    wire N__38825;
    wire N__38822;
    wire N__38819;
    wire N__38814;
    wire N__38811;
    wire N__38808;
    wire N__38805;
    wire N__38802;
    wire N__38799;
    wire N__38794;
    wire N__38793;
    wire N__38790;
    wire N__38785;
    wire N__38782;
    wire N__38779;
    wire N__38772;
    wire N__38769;
    wire N__38756;
    wire N__38755;
    wire N__38752;
    wire N__38749;
    wire N__38746;
    wire N__38743;
    wire N__38740;
    wire N__38737;
    wire N__38734;
    wire N__38731;
    wire N__38728;
    wire N__38725;
    wire N__38722;
    wire N__38719;
    wire N__38714;
    wire N__38711;
    wire N__38708;
    wire N__38707;
    wire N__38704;
    wire N__38701;
    wire N__38698;
    wire N__38697;
    wire N__38694;
    wire N__38693;
    wire N__38692;
    wire N__38689;
    wire N__38686;
    wire N__38683;
    wire N__38680;
    wire N__38677;
    wire N__38666;
    wire N__38665;
    wire N__38664;
    wire N__38661;
    wire N__38660;
    wire N__38657;
    wire N__38656;
    wire N__38653;
    wire N__38650;
    wire N__38647;
    wire N__38646;
    wire N__38643;
    wire N__38642;
    wire N__38641;
    wire N__38640;
    wire N__38637;
    wire N__38634;
    wire N__38629;
    wire N__38626;
    wire N__38625;
    wire N__38622;
    wire N__38619;
    wire N__38616;
    wire N__38613;
    wire N__38610;
    wire N__38607;
    wire N__38604;
    wire N__38603;
    wire N__38600;
    wire N__38597;
    wire N__38594;
    wire N__38591;
    wire N__38588;
    wire N__38587;
    wire N__38584;
    wire N__38579;
    wire N__38576;
    wire N__38575;
    wire N__38574;
    wire N__38573;
    wire N__38570;
    wire N__38567;
    wire N__38564;
    wire N__38559;
    wire N__38556;
    wire N__38553;
    wire N__38548;
    wire N__38545;
    wire N__38540;
    wire N__38537;
    wire N__38534;
    wire N__38523;
    wire N__38510;
    wire N__38509;
    wire N__38506;
    wire N__38503;
    wire N__38500;
    wire N__38497;
    wire N__38494;
    wire N__38491;
    wire N__38488;
    wire N__38485;
    wire N__38482;
    wire N__38479;
    wire N__38476;
    wire N__38473;
    wire N__38468;
    wire N__38467;
    wire N__38466;
    wire N__38465;
    wire N__38464;
    wire N__38463;
    wire N__38462;
    wire N__38461;
    wire N__38460;
    wire N__38459;
    wire N__38458;
    wire N__38447;
    wire N__38434;
    wire N__38429;
    wire N__38426;
    wire N__38423;
    wire N__38422;
    wire N__38419;
    wire N__38416;
    wire N__38413;
    wire N__38412;
    wire N__38409;
    wire N__38408;
    wire N__38407;
    wire N__38404;
    wire N__38401;
    wire N__38398;
    wire N__38395;
    wire N__38392;
    wire N__38381;
    wire N__38378;
    wire N__38377;
    wire N__38374;
    wire N__38371;
    wire N__38370;
    wire N__38369;
    wire N__38366;
    wire N__38363;
    wire N__38360;
    wire N__38359;
    wire N__38356;
    wire N__38355;
    wire N__38352;
    wire N__38349;
    wire N__38346;
    wire N__38343;
    wire N__38342;
    wire N__38339;
    wire N__38338;
    wire N__38337;
    wire N__38334;
    wire N__38331;
    wire N__38328;
    wire N__38327;
    wire N__38326;
    wire N__38323;
    wire N__38320;
    wire N__38317;
    wire N__38314;
    wire N__38313;
    wire N__38310;
    wire N__38307;
    wire N__38300;
    wire N__38297;
    wire N__38294;
    wire N__38289;
    wire N__38284;
    wire N__38281;
    wire N__38264;
    wire N__38263;
    wire N__38262;
    wire N__38261;
    wire N__38260;
    wire N__38259;
    wire N__38248;
    wire N__38247;
    wire N__38246;
    wire N__38245;
    wire N__38244;
    wire N__38243;
    wire N__38242;
    wire N__38239;
    wire N__38236;
    wire N__38231;
    wire N__38222;
    wire N__38219;
    wire N__38212;
    wire N__38209;
    wire N__38206;
    wire N__38203;
    wire N__38198;
    wire N__38197;
    wire N__38194;
    wire N__38191;
    wire N__38188;
    wire N__38185;
    wire N__38182;
    wire N__38179;
    wire N__38176;
    wire N__38173;
    wire N__38170;
    wire N__38167;
    wire N__38164;
    wire N__38161;
    wire N__38156;
    wire N__38155;
    wire N__38152;
    wire N__38151;
    wire N__38150;
    wire N__38145;
    wire N__38140;
    wire N__38139;
    wire N__38138;
    wire N__38137;
    wire N__38136;
    wire N__38135;
    wire N__38134;
    wire N__38133;
    wire N__38132;
    wire N__38131;
    wire N__38130;
    wire N__38129;
    wire N__38128;
    wire N__38125;
    wire N__38124;
    wire N__38123;
    wire N__38120;
    wire N__38119;
    wire N__38118;
    wire N__38117;
    wire N__38116;
    wire N__38115;
    wire N__38114;
    wire N__38113;
    wire N__38112;
    wire N__38111;
    wire N__38110;
    wire N__38109;
    wire N__38108;
    wire N__38107;
    wire N__38106;
    wire N__38105;
    wire N__38104;
    wire N__38103;
    wire N__38102;
    wire N__38101;
    wire N__38100;
    wire N__38099;
    wire N__38098;
    wire N__38097;
    wire N__38096;
    wire N__38095;
    wire N__38094;
    wire N__38093;
    wire N__38092;
    wire N__38091;
    wire N__38090;
    wire N__38089;
    wire N__38088;
    wire N__38087;
    wire N__38086;
    wire N__38085;
    wire N__38084;
    wire N__38083;
    wire N__38082;
    wire N__38081;
    wire N__38080;
    wire N__38079;
    wire N__38078;
    wire N__38077;
    wire N__38076;
    wire N__38075;
    wire N__38074;
    wire N__38073;
    wire N__38072;
    wire N__38071;
    wire N__38070;
    wire N__38069;
    wire N__38068;
    wire N__38067;
    wire N__38066;
    wire N__38065;
    wire N__38064;
    wire N__38063;
    wire N__38062;
    wire N__38061;
    wire N__38060;
    wire N__38059;
    wire N__38058;
    wire N__38057;
    wire N__38056;
    wire N__38055;
    wire N__38054;
    wire N__38053;
    wire N__38052;
    wire N__38051;
    wire N__38050;
    wire N__38049;
    wire N__38048;
    wire N__38047;
    wire N__38046;
    wire N__38045;
    wire N__38044;
    wire N__38043;
    wire N__38042;
    wire N__38041;
    wire N__38040;
    wire N__37847;
    wire N__37844;
    wire N__37841;
    wire N__37840;
    wire N__37837;
    wire N__37836;
    wire N__37835;
    wire N__37832;
    wire N__37831;
    wire N__37830;
    wire N__37827;
    wire N__37824;
    wire N__37823;
    wire N__37820;
    wire N__37819;
    wire N__37814;
    wire N__37813;
    wire N__37810;
    wire N__37809;
    wire N__37808;
    wire N__37807;
    wire N__37802;
    wire N__37799;
    wire N__37794;
    wire N__37793;
    wire N__37792;
    wire N__37791;
    wire N__37790;
    wire N__37789;
    wire N__37786;
    wire N__37783;
    wire N__37778;
    wire N__37773;
    wire N__37766;
    wire N__37763;
    wire N__37760;
    wire N__37759;
    wire N__37754;
    wire N__37753;
    wire N__37750;
    wire N__37741;
    wire N__37734;
    wire N__37733;
    wire N__37732;
    wire N__37729;
    wire N__37728;
    wire N__37725;
    wire N__37722;
    wire N__37719;
    wire N__37716;
    wire N__37713;
    wire N__37710;
    wire N__37709;
    wire N__37706;
    wire N__37701;
    wire N__37698;
    wire N__37695;
    wire N__37692;
    wire N__37685;
    wire N__37682;
    wire N__37681;
    wire N__37680;
    wire N__37679;
    wire N__37678;
    wire N__37673;
    wire N__37664;
    wire N__37661;
    wire N__37658;
    wire N__37653;
    wire N__37650;
    wire N__37637;
    wire N__37634;
    wire N__37631;
    wire N__37628;
    wire N__37627;
    wire N__37626;
    wire N__37623;
    wire N__37620;
    wire N__37617;
    wire N__37614;
    wire N__37611;
    wire N__37608;
    wire N__37605;
    wire N__37602;
    wire N__37599;
    wire N__37598;
    wire N__37597;
    wire N__37594;
    wire N__37591;
    wire N__37588;
    wire N__37585;
    wire N__37582;
    wire N__37573;
    wire N__37570;
    wire N__37567;
    wire N__37562;
    wire N__37561;
    wire N__37560;
    wire N__37557;
    wire N__37554;
    wire N__37551;
    wire N__37550;
    wire N__37549;
    wire N__37548;
    wire N__37547;
    wire N__37546;
    wire N__37545;
    wire N__37544;
    wire N__37543;
    wire N__37540;
    wire N__37537;
    wire N__37532;
    wire N__37531;
    wire N__37530;
    wire N__37527;
    wire N__37524;
    wire N__37521;
    wire N__37516;
    wire N__37511;
    wire N__37510;
    wire N__37509;
    wire N__37504;
    wire N__37503;
    wire N__37502;
    wire N__37499;
    wire N__37498;
    wire N__37497;
    wire N__37496;
    wire N__37491;
    wire N__37480;
    wire N__37479;
    wire N__37474;
    wire N__37471;
    wire N__37468;
    wire N__37467;
    wire N__37466;
    wire N__37465;
    wire N__37462;
    wire N__37461;
    wire N__37460;
    wire N__37459;
    wire N__37456;
    wire N__37453;
    wire N__37450;
    wire N__37449;
    wire N__37446;
    wire N__37441;
    wire N__37438;
    wire N__37431;
    wire N__37426;
    wire N__37423;
    wire N__37420;
    wire N__37415;
    wire N__37412;
    wire N__37407;
    wire N__37406;
    wire N__37405;
    wire N__37404;
    wire N__37401;
    wire N__37398;
    wire N__37397;
    wire N__37396;
    wire N__37393;
    wire N__37390;
    wire N__37385;
    wire N__37384;
    wire N__37381;
    wire N__37370;
    wire N__37365;
    wire N__37362;
    wire N__37359;
    wire N__37356;
    wire N__37351;
    wire N__37348;
    wire N__37343;
    wire N__37340;
    wire N__37335;
    wire N__37316;
    wire N__37313;
    wire N__37310;
    wire N__37307;
    wire N__37304;
    wire N__37303;
    wire N__37302;
    wire N__37301;
    wire N__37300;
    wire N__37299;
    wire N__37298;
    wire N__37297;
    wire N__37296;
    wire N__37293;
    wire N__37292;
    wire N__37289;
    wire N__37288;
    wire N__37287;
    wire N__37286;
    wire N__37285;
    wire N__37284;
    wire N__37283;
    wire N__37282;
    wire N__37273;
    wire N__37266;
    wire N__37265;
    wire N__37264;
    wire N__37263;
    wire N__37260;
    wire N__37257;
    wire N__37256;
    wire N__37253;
    wire N__37250;
    wire N__37249;
    wire N__37246;
    wire N__37243;
    wire N__37242;
    wire N__37239;
    wire N__37236;
    wire N__37235;
    wire N__37232;
    wire N__37231;
    wire N__37228;
    wire N__37227;
    wire N__37226;
    wire N__37221;
    wire N__37218;
    wire N__37217;
    wire N__37214;
    wire N__37213;
    wire N__37212;
    wire N__37209;
    wire N__37206;
    wire N__37203;
    wire N__37200;
    wire N__37199;
    wire N__37198;
    wire N__37195;
    wire N__37192;
    wire N__37189;
    wire N__37184;
    wire N__37181;
    wire N__37176;
    wire N__37173;
    wire N__37170;
    wire N__37167;
    wire N__37164;
    wire N__37161;
    wire N__37160;
    wire N__37159;
    wire N__37158;
    wire N__37157;
    wire N__37156;
    wire N__37155;
    wire N__37154;
    wire N__37153;
    wire N__37152;
    wire N__37151;
    wire N__37148;
    wire N__37143;
    wire N__37140;
    wire N__37137;
    wire N__37134;
    wire N__37133;
    wire N__37130;
    wire N__37129;
    wire N__37126;
    wire N__37119;
    wire N__37116;
    wire N__37113;
    wire N__37112;
    wire N__37107;
    wire N__37100;
    wire N__37095;
    wire N__37090;
    wire N__37085;
    wire N__37082;
    wire N__37079;
    wire N__37076;
    wire N__37073;
    wire N__37070;
    wire N__37067;
    wire N__37064;
    wire N__37063;
    wire N__37060;
    wire N__37057;
    wire N__37056;
    wire N__37053;
    wire N__37050;
    wire N__37047;
    wire N__37044;
    wire N__37039;
    wire N__37036;
    wire N__37033;
    wire N__37030;
    wire N__37029;
    wire N__37026;
    wire N__37019;
    wire N__37016;
    wire N__37015;
    wire N__37014;
    wire N__37013;
    wire N__37012;
    wire N__37009;
    wire N__37004;
    wire N__36997;
    wire N__36996;
    wire N__36991;
    wire N__36984;
    wire N__36975;
    wire N__36970;
    wire N__36967;
    wire N__36960;
    wire N__36957;
    wire N__36952;
    wire N__36949;
    wire N__36942;
    wire N__36939;
    wire N__36938;
    wire N__36935;
    wire N__36932;
    wire N__36929;
    wire N__36922;
    wire N__36921;
    wire N__36918;
    wire N__36915;
    wire N__36908;
    wire N__36905;
    wire N__36900;
    wire N__36891;
    wire N__36888;
    wire N__36883;
    wire N__36880;
    wire N__36877;
    wire N__36874;
    wire N__36871;
    wire N__36868;
    wire N__36865;
    wire N__36862;
    wire N__36859;
    wire N__36854;
    wire N__36851;
    wire N__36848;
    wire N__36847;
    wire N__36844;
    wire N__36841;
    wire N__36838;
    wire N__36837;
    wire N__36836;
    wire N__36831;
    wire N__36826;
    wire N__36819;
    wire N__36816;
    wire N__36809;
    wire N__36806;
    wire N__36803;
    wire N__36788;
    wire N__36787;
    wire N__36784;
    wire N__36781;
    wire N__36780;
    wire N__36777;
    wire N__36776;
    wire N__36773;
    wire N__36770;
    wire N__36767;
    wire N__36764;
    wire N__36759;
    wire N__36752;
    wire N__36751;
    wire N__36748;
    wire N__36747;
    wire N__36746;
    wire N__36745;
    wire N__36742;
    wire N__36739;
    wire N__36738;
    wire N__36735;
    wire N__36732;
    wire N__36729;
    wire N__36728;
    wire N__36727;
    wire N__36726;
    wire N__36723;
    wire N__36720;
    wire N__36717;
    wire N__36714;
    wire N__36711;
    wire N__36710;
    wire N__36707;
    wire N__36704;
    wire N__36701;
    wire N__36698;
    wire N__36697;
    wire N__36692;
    wire N__36689;
    wire N__36684;
    wire N__36681;
    wire N__36674;
    wire N__36671;
    wire N__36668;
    wire N__36665;
    wire N__36662;
    wire N__36657;
    wire N__36652;
    wire N__36649;
    wire N__36644;
    wire N__36641;
    wire N__36638;
    wire N__36629;
    wire N__36626;
    wire N__36625;
    wire N__36622;
    wire N__36619;
    wire N__36616;
    wire N__36613;
    wire N__36610;
    wire N__36607;
    wire N__36604;
    wire N__36601;
    wire N__36598;
    wire N__36595;
    wire N__36592;
    wire N__36589;
    wire N__36586;
    wire N__36581;
    wire N__36580;
    wire N__36577;
    wire N__36574;
    wire N__36573;
    wire N__36572;
    wire N__36571;
    wire N__36570;
    wire N__36569;
    wire N__36566;
    wire N__36565;
    wire N__36562;
    wire N__36559;
    wire N__36556;
    wire N__36553;
    wire N__36550;
    wire N__36547;
    wire N__36544;
    wire N__36541;
    wire N__36536;
    wire N__36531;
    wire N__36528;
    wire N__36527;
    wire N__36524;
    wire N__36523;
    wire N__36520;
    wire N__36513;
    wire N__36512;
    wire N__36509;
    wire N__36506;
    wire N__36503;
    wire N__36500;
    wire N__36499;
    wire N__36496;
    wire N__36493;
    wire N__36490;
    wire N__36481;
    wire N__36478;
    wire N__36467;
    wire N__36464;
    wire N__36463;
    wire N__36460;
    wire N__36457;
    wire N__36454;
    wire N__36453;
    wire N__36450;
    wire N__36449;
    wire N__36448;
    wire N__36445;
    wire N__36442;
    wire N__36439;
    wire N__36436;
    wire N__36433;
    wire N__36422;
    wire N__36421;
    wire N__36418;
    wire N__36415;
    wire N__36412;
    wire N__36409;
    wire N__36406;
    wire N__36403;
    wire N__36400;
    wire N__36397;
    wire N__36394;
    wire N__36391;
    wire N__36388;
    wire N__36385;
    wire N__36382;
    wire N__36377;
    wire N__36376;
    wire N__36375;
    wire N__36372;
    wire N__36369;
    wire N__36368;
    wire N__36367;
    wire N__36364;
    wire N__36363;
    wire N__36360;
    wire N__36359;
    wire N__36358;
    wire N__36357;
    wire N__36354;
    wire N__36351;
    wire N__36348;
    wire N__36347;
    wire N__36344;
    wire N__36341;
    wire N__36338;
    wire N__36337;
    wire N__36334;
    wire N__36331;
    wire N__36328;
    wire N__36325;
    wire N__36322;
    wire N__36319;
    wire N__36316;
    wire N__36313;
    wire N__36310;
    wire N__36309;
    wire N__36306;
    wire N__36303;
    wire N__36296;
    wire N__36293;
    wire N__36286;
    wire N__36283;
    wire N__36280;
    wire N__36277;
    wire N__36270;
    wire N__36257;
    wire N__36254;
    wire N__36251;
    wire N__36248;
    wire N__36247;
    wire N__36246;
    wire N__36243;
    wire N__36240;
    wire N__36237;
    wire N__36236;
    wire N__36233;
    wire N__36230;
    wire N__36227;
    wire N__36224;
    wire N__36219;
    wire N__36214;
    wire N__36209;
    wire N__36208;
    wire N__36205;
    wire N__36202;
    wire N__36199;
    wire N__36196;
    wire N__36193;
    wire N__36190;
    wire N__36187;
    wire N__36184;
    wire N__36181;
    wire N__36178;
    wire N__36175;
    wire N__36172;
    wire N__36169;
    wire N__36164;
    wire N__36161;
    wire N__36158;
    wire N__36155;
    wire N__36154;
    wire N__36151;
    wire N__36148;
    wire N__36147;
    wire N__36146;
    wire N__36143;
    wire N__36140;
    wire N__36137;
    wire N__36134;
    wire N__36127;
    wire N__36122;
    wire N__36121;
    wire N__36118;
    wire N__36115;
    wire N__36114;
    wire N__36113;
    wire N__36110;
    wire N__36107;
    wire N__36104;
    wire N__36103;
    wire N__36100;
    wire N__36097;
    wire N__36096;
    wire N__36093;
    wire N__36092;
    wire N__36089;
    wire N__36086;
    wire N__36083;
    wire N__36080;
    wire N__36077;
    wire N__36076;
    wire N__36073;
    wire N__36070;
    wire N__36067;
    wire N__36064;
    wire N__36057;
    wire N__36054;
    wire N__36051;
    wire N__36050;
    wire N__36045;
    wire N__36044;
    wire N__36043;
    wire N__36040;
    wire N__36037;
    wire N__36034;
    wire N__36031;
    wire N__36028;
    wire N__36025;
    wire N__36022;
    wire N__36019;
    wire N__36012;
    wire N__35999;
    wire N__35998;
    wire N__35995;
    wire N__35992;
    wire N__35989;
    wire N__35986;
    wire N__35983;
    wire N__35980;
    wire N__35977;
    wire N__35974;
    wire N__35971;
    wire N__35968;
    wire N__35965;
    wire N__35962;
    wire N__35959;
    wire N__35954;
    wire N__35953;
    wire N__35952;
    wire N__35949;
    wire N__35946;
    wire N__35943;
    wire N__35940;
    wire N__35939;
    wire N__35938;
    wire N__35937;
    wire N__35934;
    wire N__35933;
    wire N__35930;
    wire N__35927;
    wire N__35924;
    wire N__35921;
    wire N__35920;
    wire N__35919;
    wire N__35916;
    wire N__35915;
    wire N__35912;
    wire N__35911;
    wire N__35910;
    wire N__35907;
    wire N__35904;
    wire N__35897;
    wire N__35892;
    wire N__35889;
    wire N__35886;
    wire N__35883;
    wire N__35880;
    wire N__35877;
    wire N__35874;
    wire N__35871;
    wire N__35866;
    wire N__35863;
    wire N__35860;
    wire N__35857;
    wire N__35854;
    wire N__35847;
    wire N__35844;
    wire N__35831;
    wire N__35828;
    wire N__35827;
    wire N__35824;
    wire N__35823;
    wire N__35820;
    wire N__35819;
    wire N__35816;
    wire N__35813;
    wire N__35812;
    wire N__35809;
    wire N__35806;
    wire N__35803;
    wire N__35800;
    wire N__35797;
    wire N__35792;
    wire N__35789;
    wire N__35786;
    wire N__35783;
    wire N__35780;
    wire N__35771;
    wire N__35770;
    wire N__35767;
    wire N__35764;
    wire N__35761;
    wire N__35758;
    wire N__35755;
    wire N__35752;
    wire N__35749;
    wire N__35746;
    wire N__35743;
    wire N__35740;
    wire N__35737;
    wire N__35734;
    wire N__35731;
    wire N__35726;
    wire N__35723;
    wire N__35722;
    wire N__35719;
    wire N__35716;
    wire N__35715;
    wire N__35712;
    wire N__35711;
    wire N__35710;
    wire N__35707;
    wire N__35706;
    wire N__35705;
    wire N__35702;
    wire N__35701;
    wire N__35700;
    wire N__35697;
    wire N__35694;
    wire N__35691;
    wire N__35690;
    wire N__35687;
    wire N__35684;
    wire N__35683;
    wire N__35682;
    wire N__35679;
    wire N__35676;
    wire N__35673;
    wire N__35670;
    wire N__35669;
    wire N__35664;
    wire N__35661;
    wire N__35658;
    wire N__35655;
    wire N__35652;
    wire N__35649;
    wire N__35646;
    wire N__35641;
    wire N__35636;
    wire N__35633;
    wire N__35626;
    wire N__35621;
    wire N__35618;
    wire N__35615;
    wire N__35608;
    wire N__35605;
    wire N__35594;
    wire N__35591;
    wire N__35588;
    wire N__35585;
    wire N__35584;
    wire N__35581;
    wire N__35578;
    wire N__35577;
    wire N__35572;
    wire N__35571;
    wire N__35570;
    wire N__35567;
    wire N__35564;
    wire N__35561;
    wire N__35558;
    wire N__35549;
    wire N__35548;
    wire N__35545;
    wire N__35542;
    wire N__35539;
    wire N__35536;
    wire N__35533;
    wire N__35530;
    wire N__35527;
    wire N__35524;
    wire N__35521;
    wire N__35518;
    wire N__35515;
    wire N__35512;
    wire N__35509;
    wire N__35504;
    wire N__35501;
    wire N__35500;
    wire N__35497;
    wire N__35494;
    wire N__35493;
    wire N__35488;
    wire N__35485;
    wire N__35484;
    wire N__35479;
    wire N__35476;
    wire N__35473;
    wire N__35470;
    wire N__35467;
    wire N__35462;
    wire N__35459;
    wire N__35456;
    wire N__35453;
    wire N__35450;
    wire N__35447;
    wire N__35444;
    wire N__35441;
    wire N__35438;
    wire N__35435;
    wire N__35432;
    wire N__35429;
    wire N__35426;
    wire N__35423;
    wire N__35420;
    wire N__35417;
    wire N__35414;
    wire N__35411;
    wire N__35410;
    wire N__35407;
    wire N__35404;
    wire N__35401;
    wire N__35398;
    wire N__35395;
    wire N__35392;
    wire N__35389;
    wire N__35386;
    wire N__35383;
    wire N__35380;
    wire N__35377;
    wire N__35374;
    wire N__35371;
    wire N__35368;
    wire N__35365;
    wire N__35362;
    wire N__35359;
    wire N__35356;
    wire N__35353;
    wire N__35350;
    wire N__35347;
    wire N__35344;
    wire N__35341;
    wire N__35338;
    wire N__35335;
    wire N__35330;
    wire N__35327;
    wire N__35326;
    wire N__35323;
    wire N__35322;
    wire N__35319;
    wire N__35316;
    wire N__35315;
    wire N__35312;
    wire N__35309;
    wire N__35306;
    wire N__35303;
    wire N__35300;
    wire N__35297;
    wire N__35294;
    wire N__35291;
    wire N__35288;
    wire N__35285;
    wire N__35280;
    wire N__35277;
    wire N__35270;
    wire N__35267;
    wire N__35264;
    wire N__35261;
    wire N__35258;
    wire N__35255;
    wire N__35252;
    wire N__35249;
    wire N__35246;
    wire N__35243;
    wire N__35242;
    wire N__35241;
    wire N__35240;
    wire N__35239;
    wire N__35238;
    wire N__35237;
    wire N__35228;
    wire N__35223;
    wire N__35220;
    wire N__35219;
    wire N__35218;
    wire N__35217;
    wire N__35216;
    wire N__35215;
    wire N__35210;
    wire N__35209;
    wire N__35208;
    wire N__35207;
    wire N__35204;
    wire N__35197;
    wire N__35196;
    wire N__35193;
    wire N__35190;
    wire N__35189;
    wire N__35188;
    wire N__35187;
    wire N__35186;
    wire N__35185;
    wire N__35182;
    wire N__35179;
    wire N__35176;
    wire N__35173;
    wire N__35172;
    wire N__35167;
    wire N__35166;
    wire N__35163;
    wire N__35160;
    wire N__35157;
    wire N__35148;
    wire N__35145;
    wire N__35140;
    wire N__35137;
    wire N__35134;
    wire N__35131;
    wire N__35128;
    wire N__35125;
    wire N__35122;
    wire N__35119;
    wire N__35116;
    wire N__35113;
    wire N__35108;
    wire N__35105;
    wire N__35100;
    wire N__35095;
    wire N__35092;
    wire N__35075;
    wire N__35072;
    wire N__35069;
    wire N__35066;
    wire N__35063;
    wire N__35060;
    wire N__35057;
    wire N__35056;
    wire N__35053;
    wire N__35050;
    wire N__35047;
    wire N__35044;
    wire N__35041;
    wire N__35038;
    wire N__35035;
    wire N__35032;
    wire N__35029;
    wire N__35026;
    wire N__35023;
    wire N__35020;
    wire N__35017;
    wire N__35014;
    wire N__35011;
    wire N__35008;
    wire N__35005;
    wire N__35002;
    wire N__34999;
    wire N__34996;
    wire N__34993;
    wire N__34990;
    wire N__34987;
    wire N__34984;
    wire N__34979;
    wire N__34976;
    wire N__34975;
    wire N__34974;
    wire N__34973;
    wire N__34970;
    wire N__34967;
    wire N__34966;
    wire N__34963;
    wire N__34960;
    wire N__34957;
    wire N__34954;
    wire N__34951;
    wire N__34948;
    wire N__34945;
    wire N__34942;
    wire N__34939;
    wire N__34936;
    wire N__34931;
    wire N__34928;
    wire N__34921;
    wire N__34916;
    wire N__34913;
    wire N__34910;
    wire N__34909;
    wire N__34908;
    wire N__34907;
    wire N__34904;
    wire N__34903;
    wire N__34900;
    wire N__34897;
    wire N__34894;
    wire N__34891;
    wire N__34888;
    wire N__34885;
    wire N__34874;
    wire N__34871;
    wire N__34870;
    wire N__34867;
    wire N__34866;
    wire N__34865;
    wire N__34862;
    wire N__34859;
    wire N__34856;
    wire N__34853;
    wire N__34844;
    wire N__34841;
    wire N__34840;
    wire N__34839;
    wire N__34838;
    wire N__34835;
    wire N__34832;
    wire N__34829;
    wire N__34826;
    wire N__34825;
    wire N__34822;
    wire N__34819;
    wire N__34816;
    wire N__34813;
    wire N__34810;
    wire N__34807;
    wire N__34804;
    wire N__34801;
    wire N__34798;
    wire N__34795;
    wire N__34792;
    wire N__34787;
    wire N__34782;
    wire N__34775;
    wire N__34772;
    wire N__34769;
    wire N__34766;
    wire N__34765;
    wire N__34764;
    wire N__34763;
    wire N__34762;
    wire N__34761;
    wire N__34758;
    wire N__34755;
    wire N__34752;
    wire N__34747;
    wire N__34746;
    wire N__34745;
    wire N__34742;
    wire N__34741;
    wire N__34738;
    wire N__34731;
    wire N__34728;
    wire N__34727;
    wire N__34726;
    wire N__34725;
    wire N__34722;
    wire N__34719;
    wire N__34716;
    wire N__34713;
    wire N__34710;
    wire N__34707;
    wire N__34706;
    wire N__34703;
    wire N__34698;
    wire N__34695;
    wire N__34694;
    wire N__34691;
    wire N__34688;
    wire N__34681;
    wire N__34676;
    wire N__34673;
    wire N__34670;
    wire N__34667;
    wire N__34652;
    wire N__34649;
    wire N__34646;
    wire N__34643;
    wire N__34642;
    wire N__34639;
    wire N__34636;
    wire N__34633;
    wire N__34630;
    wire N__34629;
    wire N__34628;
    wire N__34627;
    wire N__34626;
    wire N__34625;
    wire N__34624;
    wire N__34623;
    wire N__34620;
    wire N__34617;
    wire N__34610;
    wire N__34607;
    wire N__34604;
    wire N__34599;
    wire N__34592;
    wire N__34589;
    wire N__34588;
    wire N__34583;
    wire N__34582;
    wire N__34579;
    wire N__34576;
    wire N__34573;
    wire N__34570;
    wire N__34567;
    wire N__34556;
    wire N__34553;
    wire N__34550;
    wire N__34549;
    wire N__34546;
    wire N__34545;
    wire N__34542;
    wire N__34539;
    wire N__34536;
    wire N__34529;
    wire N__34528;
    wire N__34527;
    wire N__34526;
    wire N__34525;
    wire N__34524;
    wire N__34523;
    wire N__34522;
    wire N__34521;
    wire N__34520;
    wire N__34519;
    wire N__34518;
    wire N__34517;
    wire N__34516;
    wire N__34515;
    wire N__34514;
    wire N__34513;
    wire N__34512;
    wire N__34511;
    wire N__34510;
    wire N__34509;
    wire N__34508;
    wire N__34507;
    wire N__34506;
    wire N__34505;
    wire N__34504;
    wire N__34503;
    wire N__34502;
    wire N__34501;
    wire N__34500;
    wire N__34499;
    wire N__34498;
    wire N__34497;
    wire N__34496;
    wire N__34495;
    wire N__34494;
    wire N__34493;
    wire N__34492;
    wire N__34491;
    wire N__34490;
    wire N__34489;
    wire N__34488;
    wire N__34487;
    wire N__34486;
    wire N__34485;
    wire N__34484;
    wire N__34483;
    wire N__34482;
    wire N__34481;
    wire N__34480;
    wire N__34479;
    wire N__34478;
    wire N__34477;
    wire N__34476;
    wire N__34475;
    wire N__34474;
    wire N__34473;
    wire N__34472;
    wire N__34471;
    wire N__34470;
    wire N__34469;
    wire N__34468;
    wire N__34467;
    wire N__34466;
    wire N__34465;
    wire N__34464;
    wire N__34463;
    wire N__34462;
    wire N__34461;
    wire N__34460;
    wire N__34459;
    wire N__34458;
    wire N__34457;
    wire N__34456;
    wire N__34455;
    wire N__34454;
    wire N__34453;
    wire N__34452;
    wire N__34451;
    wire N__34450;
    wire N__34449;
    wire N__34448;
    wire N__34447;
    wire N__34446;
    wire N__34445;
    wire N__34444;
    wire N__34443;
    wire N__34442;
    wire N__34441;
    wire N__34440;
    wire N__34439;
    wire N__34438;
    wire N__34437;
    wire N__34436;
    wire N__34435;
    wire N__34434;
    wire N__34433;
    wire N__34432;
    wire N__34431;
    wire N__34430;
    wire N__34429;
    wire N__34428;
    wire N__34427;
    wire N__34426;
    wire N__34425;
    wire N__34424;
    wire N__34423;
    wire N__34422;
    wire N__34421;
    wire N__34420;
    wire N__34419;
    wire N__34418;
    wire N__34417;
    wire N__34416;
    wire N__34415;
    wire N__34414;
    wire N__34413;
    wire N__34412;
    wire N__34411;
    wire N__34410;
    wire N__34409;
    wire N__34408;
    wire N__34407;
    wire N__34406;
    wire N__34405;
    wire N__34404;
    wire N__34403;
    wire N__34402;
    wire N__34401;
    wire N__34400;
    wire N__34399;
    wire N__34398;
    wire N__34397;
    wire N__34396;
    wire N__34395;
    wire N__34394;
    wire N__34393;
    wire N__34392;
    wire N__34391;
    wire N__34390;
    wire N__34389;
    wire N__34388;
    wire N__34387;
    wire N__34386;
    wire N__34385;
    wire N__34384;
    wire N__34383;
    wire N__34382;
    wire N__34381;
    wire N__34380;
    wire N__34379;
    wire N__34378;
    wire N__34377;
    wire N__34376;
    wire N__34375;
    wire N__34374;
    wire N__34373;
    wire N__34372;
    wire N__34371;
    wire N__34052;
    wire N__34049;
    wire N__34046;
    wire N__34043;
    wire N__34040;
    wire N__34037;
    wire N__34034;
    wire N__34031;
    wire N__34028;
    wire N__34025;
    wire N__34022;
    wire N__34019;
    wire N__34016;
    wire N__34013;
    wire N__34010;
    wire N__34009;
    wire N__34006;
    wire N__34003;
    wire N__34000;
    wire N__33997;
    wire N__33994;
    wire N__33991;
    wire N__33988;
    wire N__33985;
    wire N__33982;
    wire N__33979;
    wire N__33976;
    wire N__33973;
    wire N__33970;
    wire N__33967;
    wire N__33964;
    wire N__33961;
    wire N__33958;
    wire N__33955;
    wire N__33952;
    wire N__33949;
    wire N__33946;
    wire N__33943;
    wire N__33940;
    wire N__33937;
    wire N__33934;
    wire N__33929;
    wire N__33926;
    wire N__33923;
    wire N__33920;
    wire N__33917;
    wire N__33914;
    wire N__33911;
    wire N__33908;
    wire N__33905;
    wire N__33902;
    wire N__33899;
    wire N__33896;
    wire N__33893;
    wire N__33892;
    wire N__33889;
    wire N__33886;
    wire N__33883;
    wire N__33880;
    wire N__33877;
    wire N__33874;
    wire N__33871;
    wire N__33868;
    wire N__33865;
    wire N__33862;
    wire N__33859;
    wire N__33856;
    wire N__33853;
    wire N__33850;
    wire N__33847;
    wire N__33844;
    wire N__33841;
    wire N__33838;
    wire N__33835;
    wire N__33832;
    wire N__33829;
    wire N__33826;
    wire N__33823;
    wire N__33820;
    wire N__33817;
    wire N__33812;
    wire N__33809;
    wire N__33806;
    wire N__33803;
    wire N__33800;
    wire N__33797;
    wire N__33794;
    wire N__33791;
    wire N__33788;
    wire N__33785;
    wire N__33782;
    wire N__33779;
    wire N__33778;
    wire N__33775;
    wire N__33772;
    wire N__33769;
    wire N__33766;
    wire N__33763;
    wire N__33760;
    wire N__33757;
    wire N__33754;
    wire N__33751;
    wire N__33748;
    wire N__33745;
    wire N__33742;
    wire N__33739;
    wire N__33736;
    wire N__33733;
    wire N__33730;
    wire N__33727;
    wire N__33724;
    wire N__33721;
    wire N__33718;
    wire N__33715;
    wire N__33712;
    wire N__33709;
    wire N__33706;
    wire N__33703;
    wire N__33698;
    wire N__33695;
    wire N__33692;
    wire N__33689;
    wire N__33686;
    wire N__33683;
    wire N__33682;
    wire N__33679;
    wire N__33676;
    wire N__33673;
    wire N__33670;
    wire N__33669;
    wire N__33664;
    wire N__33661;
    wire N__33658;
    wire N__33655;
    wire N__33652;
    wire N__33649;
    wire N__33648;
    wire N__33645;
    wire N__33642;
    wire N__33639;
    wire N__33632;
    wire N__33629;
    wire N__33626;
    wire N__33623;
    wire N__33620;
    wire N__33617;
    wire N__33614;
    wire N__33611;
    wire N__33608;
    wire N__33605;
    wire N__33602;
    wire N__33599;
    wire N__33596;
    wire N__33593;
    wire N__33590;
    wire N__33589;
    wire N__33586;
    wire N__33583;
    wire N__33580;
    wire N__33577;
    wire N__33574;
    wire N__33571;
    wire N__33568;
    wire N__33565;
    wire N__33562;
    wire N__33559;
    wire N__33556;
    wire N__33553;
    wire N__33550;
    wire N__33547;
    wire N__33544;
    wire N__33541;
    wire N__33538;
    wire N__33535;
    wire N__33532;
    wire N__33529;
    wire N__33526;
    wire N__33523;
    wire N__33520;
    wire N__33517;
    wire N__33512;
    wire N__33509;
    wire N__33506;
    wire N__33503;
    wire N__33500;
    wire N__33497;
    wire N__33494;
    wire N__33491;
    wire N__33488;
    wire N__33485;
    wire N__33482;
    wire N__33479;
    wire N__33476;
    wire N__33475;
    wire N__33472;
    wire N__33469;
    wire N__33466;
    wire N__33463;
    wire N__33460;
    wire N__33457;
    wire N__33454;
    wire N__33451;
    wire N__33448;
    wire N__33445;
    wire N__33442;
    wire N__33439;
    wire N__33436;
    wire N__33433;
    wire N__33430;
    wire N__33427;
    wire N__33424;
    wire N__33421;
    wire N__33418;
    wire N__33415;
    wire N__33412;
    wire N__33409;
    wire N__33406;
    wire N__33403;
    wire N__33398;
    wire N__33397;
    wire N__33394;
    wire N__33391;
    wire N__33388;
    wire N__33385;
    wire N__33382;
    wire N__33381;
    wire N__33380;
    wire N__33375;
    wire N__33372;
    wire N__33369;
    wire N__33366;
    wire N__33361;
    wire N__33356;
    wire N__33353;
    wire N__33350;
    wire N__33347;
    wire N__33344;
    wire N__33341;
    wire N__33338;
    wire N__33337;
    wire N__33336;
    wire N__33333;
    wire N__33330;
    wire N__33329;
    wire N__33326;
    wire N__33325;
    wire N__33322;
    wire N__33319;
    wire N__33316;
    wire N__33313;
    wire N__33310;
    wire N__33305;
    wire N__33302;
    wire N__33297;
    wire N__33294;
    wire N__33291;
    wire N__33288;
    wire N__33285;
    wire N__33280;
    wire N__33275;
    wire N__33272;
    wire N__33269;
    wire N__33266;
    wire N__33263;
    wire N__33260;
    wire N__33257;
    wire N__33256;
    wire N__33255;
    wire N__33254;
    wire N__33251;
    wire N__33248;
    wire N__33245;
    wire N__33244;
    wire N__33241;
    wire N__33238;
    wire N__33235;
    wire N__33232;
    wire N__33229;
    wire N__33226;
    wire N__33223;
    wire N__33218;
    wire N__33215;
    wire N__33212;
    wire N__33207;
    wire N__33200;
    wire N__33197;
    wire N__33194;
    wire N__33191;
    wire N__33188;
    wire N__33187;
    wire N__33184;
    wire N__33181;
    wire N__33180;
    wire N__33177;
    wire N__33174;
    wire N__33171;
    wire N__33168;
    wire N__33167;
    wire N__33164;
    wire N__33159;
    wire N__33156;
    wire N__33153;
    wire N__33146;
    wire N__33143;
    wire N__33140;
    wire N__33139;
    wire N__33136;
    wire N__33135;
    wire N__33132;
    wire N__33131;
    wire N__33128;
    wire N__33125;
    wire N__33124;
    wire N__33121;
    wire N__33118;
    wire N__33115;
    wire N__33112;
    wire N__33109;
    wire N__33106;
    wire N__33103;
    wire N__33100;
    wire N__33097;
    wire N__33094;
    wire N__33089;
    wire N__33084;
    wire N__33081;
    wire N__33078;
    wire N__33071;
    wire N__33068;
    wire N__33065;
    wire N__33062;
    wire N__33061;
    wire N__33058;
    wire N__33055;
    wire N__33054;
    wire N__33051;
    wire N__33050;
    wire N__33047;
    wire N__33044;
    wire N__33041;
    wire N__33038;
    wire N__33035;
    wire N__33030;
    wire N__33027;
    wire N__33020;
    wire N__33019;
    wire N__33016;
    wire N__33015;
    wire N__33014;
    wire N__33011;
    wire N__33010;
    wire N__33007;
    wire N__33004;
    wire N__33001;
    wire N__32998;
    wire N__32995;
    wire N__32992;
    wire N__32989;
    wire N__32986;
    wire N__32983;
    wire N__32980;
    wire N__32975;
    wire N__32966;
    wire N__32965;
    wire N__32964;
    wire N__32963;
    wire N__32960;
    wire N__32959;
    wire N__32958;
    wire N__32955;
    wire N__32952;
    wire N__32949;
    wire N__32946;
    wire N__32943;
    wire N__32940;
    wire N__32937;
    wire N__32934;
    wire N__32931;
    wire N__32930;
    wire N__32925;
    wire N__32922;
    wire N__32919;
    wire N__32914;
    wire N__32911;
    wire N__32900;
    wire N__32899;
    wire N__32898;
    wire N__32897;
    wire N__32896;
    wire N__32893;
    wire N__32890;
    wire N__32885;
    wire N__32882;
    wire N__32873;
    wire N__32872;
    wire N__32869;
    wire N__32866;
    wire N__32863;
    wire N__32860;
    wire N__32859;
    wire N__32854;
    wire N__32853;
    wire N__32850;
    wire N__32847;
    wire N__32844;
    wire N__32841;
    wire N__32836;
    wire N__32833;
    wire N__32830;
    wire N__32825;
    wire N__32822;
    wire N__32819;
    wire N__32816;
    wire N__32813;
    wire N__32810;
    wire N__32807;
    wire N__32804;
    wire N__32801;
    wire N__32798;
    wire N__32795;
    wire N__32792;
    wire N__32789;
    wire N__32786;
    wire N__32785;
    wire N__32782;
    wire N__32779;
    wire N__32776;
    wire N__32773;
    wire N__32770;
    wire N__32767;
    wire N__32764;
    wire N__32761;
    wire N__32758;
    wire N__32755;
    wire N__32752;
    wire N__32749;
    wire N__32746;
    wire N__32743;
    wire N__32740;
    wire N__32737;
    wire N__32734;
    wire N__32731;
    wire N__32728;
    wire N__32725;
    wire N__32722;
    wire N__32719;
    wire N__32716;
    wire N__32713;
    wire N__32710;
    wire N__32705;
    wire N__32702;
    wire N__32699;
    wire N__32696;
    wire N__32693;
    wire N__32690;
    wire N__32687;
    wire N__32684;
    wire N__32681;
    wire N__32678;
    wire N__32675;
    wire N__32672;
    wire N__32669;
    wire N__32666;
    wire N__32663;
    wire N__32660;
    wire N__32657;
    wire N__32656;
    wire N__32653;
    wire N__32652;
    wire N__32649;
    wire N__32646;
    wire N__32643;
    wire N__32636;
    wire N__32633;
    wire N__32630;
    wire N__32627;
    wire N__32624;
    wire N__32623;
    wire N__32620;
    wire N__32619;
    wire N__32616;
    wire N__32613;
    wire N__32610;
    wire N__32603;
    wire N__32600;
    wire N__32599;
    wire N__32596;
    wire N__32593;
    wire N__32590;
    wire N__32587;
    wire N__32586;
    wire N__32583;
    wire N__32580;
    wire N__32577;
    wire N__32572;
    wire N__32567;
    wire N__32564;
    wire N__32561;
    wire N__32558;
    wire N__32555;
    wire N__32552;
    wire N__32549;
    wire N__32546;
    wire N__32545;
    wire N__32544;
    wire N__32543;
    wire N__32542;
    wire N__32541;
    wire N__32540;
    wire N__32539;
    wire N__32538;
    wire N__32537;
    wire N__32536;
    wire N__32535;
    wire N__32530;
    wire N__32525;
    wire N__32522;
    wire N__32517;
    wire N__32514;
    wire N__32511;
    wire N__32506;
    wire N__32503;
    wire N__32500;
    wire N__32497;
    wire N__32494;
    wire N__32485;
    wire N__32482;
    wire N__32477;
    wire N__32474;
    wire N__32465;
    wire N__32462;
    wire N__32459;
    wire N__32458;
    wire N__32455;
    wire N__32452;
    wire N__32449;
    wire N__32448;
    wire N__32445;
    wire N__32442;
    wire N__32439;
    wire N__32438;
    wire N__32435;
    wire N__32434;
    wire N__32429;
    wire N__32426;
    wire N__32423;
    wire N__32420;
    wire N__32417;
    wire N__32408;
    wire N__32407;
    wire N__32406;
    wire N__32405;
    wire N__32402;
    wire N__32399;
    wire N__32398;
    wire N__32397;
    wire N__32396;
    wire N__32395;
    wire N__32394;
    wire N__32393;
    wire N__32392;
    wire N__32391;
    wire N__32386;
    wire N__32383;
    wire N__32380;
    wire N__32377;
    wire N__32374;
    wire N__32369;
    wire N__32366;
    wire N__32359;
    wire N__32350;
    wire N__32349;
    wire N__32344;
    wire N__32341;
    wire N__32336;
    wire N__32333;
    wire N__32324;
    wire N__32321;
    wire N__32318;
    wire N__32315;
    wire N__32312;
    wire N__32309;
    wire N__32306;
    wire N__32305;
    wire N__32302;
    wire N__32301;
    wire N__32298;
    wire N__32295;
    wire N__32292;
    wire N__32285;
    wire N__32284;
    wire N__32283;
    wire N__32282;
    wire N__32279;
    wire N__32276;
    wire N__32273;
    wire N__32270;
    wire N__32267;
    wire N__32264;
    wire N__32261;
    wire N__32258;
    wire N__32255;
    wire N__32252;
    wire N__32249;
    wire N__32246;
    wire N__32241;
    wire N__32236;
    wire N__32231;
    wire N__32230;
    wire N__32229;
    wire N__32226;
    wire N__32223;
    wire N__32220;
    wire N__32215;
    wire N__32210;
    wire N__32209;
    wire N__32206;
    wire N__32205;
    wire N__32204;
    wire N__32201;
    wire N__32198;
    wire N__32195;
    wire N__32192;
    wire N__32189;
    wire N__32186;
    wire N__32183;
    wire N__32180;
    wire N__32177;
    wire N__32172;
    wire N__32169;
    wire N__32166;
    wire N__32163;
    wire N__32160;
    wire N__32153;
    wire N__32152;
    wire N__32151;
    wire N__32148;
    wire N__32145;
    wire N__32142;
    wire N__32139;
    wire N__32132;
    wire N__32131;
    wire N__32128;
    wire N__32125;
    wire N__32124;
    wire N__32121;
    wire N__32118;
    wire N__32117;
    wire N__32114;
    wire N__32111;
    wire N__32108;
    wire N__32105;
    wire N__32102;
    wire N__32099;
    wire N__32096;
    wire N__32093;
    wire N__32084;
    wire N__32083;
    wire N__32082;
    wire N__32079;
    wire N__32076;
    wire N__32073;
    wire N__32070;
    wire N__32065;
    wire N__32060;
    wire N__32059;
    wire N__32056;
    wire N__32053;
    wire N__32052;
    wire N__32051;
    wire N__32048;
    wire N__32045;
    wire N__32042;
    wire N__32039;
    wire N__32036;
    wire N__32033;
    wire N__32030;
    wire N__32027;
    wire N__32026;
    wire N__32025;
    wire N__32024;
    wire N__32021;
    wire N__32016;
    wire N__32013;
    wire N__32008;
    wire N__32005;
    wire N__31994;
    wire N__31993;
    wire N__31990;
    wire N__31989;
    wire N__31986;
    wire N__31985;
    wire N__31982;
    wire N__31979;
    wire N__31976;
    wire N__31973;
    wire N__31966;
    wire N__31963;
    wire N__31958;
    wire N__31955;
    wire N__31954;
    wire N__31951;
    wire N__31950;
    wire N__31947;
    wire N__31946;
    wire N__31943;
    wire N__31940;
    wire N__31937;
    wire N__31934;
    wire N__31931;
    wire N__31928;
    wire N__31919;
    wire N__31918;
    wire N__31917;
    wire N__31914;
    wire N__31909;
    wire N__31908;
    wire N__31907;
    wire N__31906;
    wire N__31905;
    wire N__31904;
    wire N__31903;
    wire N__31902;
    wire N__31901;
    wire N__31900;
    wire N__31899;
    wire N__31898;
    wire N__31897;
    wire N__31896;
    wire N__31895;
    wire N__31894;
    wire N__31889;
    wire N__31876;
    wire N__31873;
    wire N__31864;
    wire N__31859;
    wire N__31858;
    wire N__31853;
    wire N__31848;
    wire N__31843;
    wire N__31840;
    wire N__31837;
    wire N__31834;
    wire N__31833;
    wire N__31832;
    wire N__31831;
    wire N__31828;
    wire N__31825;
    wire N__31820;
    wire N__31817;
    wire N__31814;
    wire N__31809;
    wire N__31802;
    wire N__31795;
    wire N__31792;
    wire N__31789;
    wire N__31786;
    wire N__31781;
    wire N__31780;
    wire N__31777;
    wire N__31776;
    wire N__31773;
    wire N__31772;
    wire N__31769;
    wire N__31766;
    wire N__31763;
    wire N__31760;
    wire N__31757;
    wire N__31754;
    wire N__31751;
    wire N__31748;
    wire N__31745;
    wire N__31742;
    wire N__31737;
    wire N__31730;
    wire N__31727;
    wire N__31726;
    wire N__31723;
    wire N__31720;
    wire N__31719;
    wire N__31718;
    wire N__31715;
    wire N__31712;
    wire N__31709;
    wire N__31706;
    wire N__31703;
    wire N__31700;
    wire N__31697;
    wire N__31688;
    wire N__31687;
    wire N__31686;
    wire N__31683;
    wire N__31680;
    wire N__31677;
    wire N__31674;
    wire N__31673;
    wire N__31672;
    wire N__31671;
    wire N__31668;
    wire N__31667;
    wire N__31666;
    wire N__31663;
    wire N__31660;
    wire N__31657;
    wire N__31654;
    wire N__31651;
    wire N__31648;
    wire N__31645;
    wire N__31642;
    wire N__31639;
    wire N__31634;
    wire N__31631;
    wire N__31626;
    wire N__31623;
    wire N__31622;
    wire N__31619;
    wire N__31614;
    wire N__31613;
    wire N__31610;
    wire N__31605;
    wire N__31604;
    wire N__31601;
    wire N__31598;
    wire N__31595;
    wire N__31592;
    wire N__31587;
    wire N__31584;
    wire N__31571;
    wire N__31570;
    wire N__31567;
    wire N__31564;
    wire N__31563;
    wire N__31562;
    wire N__31559;
    wire N__31556;
    wire N__31553;
    wire N__31550;
    wire N__31543;
    wire N__31540;
    wire N__31537;
    wire N__31534;
    wire N__31529;
    wire N__31526;
    wire N__31525;
    wire N__31522;
    wire N__31519;
    wire N__31518;
    wire N__31515;
    wire N__31514;
    wire N__31511;
    wire N__31508;
    wire N__31505;
    wire N__31502;
    wire N__31499;
    wire N__31490;
    wire N__31489;
    wire N__31488;
    wire N__31487;
    wire N__31484;
    wire N__31483;
    wire N__31480;
    wire N__31477;
    wire N__31474;
    wire N__31471;
    wire N__31468;
    wire N__31465;
    wire N__31462;
    wire N__31459;
    wire N__31450;
    wire N__31445;
    wire N__31442;
    wire N__31439;
    wire N__31438;
    wire N__31435;
    wire N__31432;
    wire N__31427;
    wire N__31426;
    wire N__31423;
    wire N__31420;
    wire N__31415;
    wire N__31412;
    wire N__31409;
    wire N__31406;
    wire N__31403;
    wire N__31400;
    wire N__31397;
    wire N__31396;
    wire N__31395;
    wire N__31394;
    wire N__31391;
    wire N__31388;
    wire N__31385;
    wire N__31382;
    wire N__31377;
    wire N__31374;
    wire N__31371;
    wire N__31368;
    wire N__31363;
    wire N__31360;
    wire N__31357;
    wire N__31352;
    wire N__31351;
    wire N__31350;
    wire N__31347;
    wire N__31346;
    wire N__31343;
    wire N__31340;
    wire N__31337;
    wire N__31334;
    wire N__31331;
    wire N__31330;
    wire N__31327;
    wire N__31322;
    wire N__31319;
    wire N__31316;
    wire N__31311;
    wire N__31304;
    wire N__31301;
    wire N__31300;
    wire N__31299;
    wire N__31296;
    wire N__31293;
    wire N__31290;
    wire N__31287;
    wire N__31284;
    wire N__31283;
    wire N__31282;
    wire N__31279;
    wire N__31276;
    wire N__31273;
    wire N__31268;
    wire N__31265;
    wire N__31256;
    wire N__31255;
    wire N__31252;
    wire N__31249;
    wire N__31246;
    wire N__31245;
    wire N__31242;
    wire N__31241;
    wire N__31238;
    wire N__31235;
    wire N__31232;
    wire N__31229;
    wire N__31224;
    wire N__31223;
    wire N__31220;
    wire N__31217;
    wire N__31214;
    wire N__31211;
    wire N__31202;
    wire N__31199;
    wire N__31196;
    wire N__31195;
    wire N__31192;
    wire N__31189;
    wire N__31184;
    wire N__31181;
    wire N__31180;
    wire N__31179;
    wire N__31178;
    wire N__31177;
    wire N__31176;
    wire N__31175;
    wire N__31174;
    wire N__31173;
    wire N__31172;
    wire N__31171;
    wire N__31170;
    wire N__31169;
    wire N__31168;
    wire N__31167;
    wire N__31166;
    wire N__31165;
    wire N__31164;
    wire N__31161;
    wire N__31158;
    wire N__31151;
    wire N__31148;
    wire N__31139;
    wire N__31130;
    wire N__31129;
    wire N__31120;
    wire N__31119;
    wire N__31118;
    wire N__31117;
    wire N__31116;
    wire N__31115;
    wire N__31114;
    wire N__31113;
    wire N__31112;
    wire N__31111;
    wire N__31110;
    wire N__31105;
    wire N__31096;
    wire N__31093;
    wire N__31090;
    wire N__31077;
    wire N__31068;
    wire N__31061;
    wire N__31056;
    wire N__31049;
    wire N__31046;
    wire N__31043;
    wire N__31042;
    wire N__31041;
    wire N__31038;
    wire N__31037;
    wire N__31034;
    wire N__31031;
    wire N__31028;
    wire N__31025;
    wire N__31022;
    wire N__31019;
    wire N__31014;
    wire N__31011;
    wire N__31010;
    wire N__31007;
    wire N__31002;
    wire N__30999;
    wire N__30992;
    wire N__30991;
    wire N__30990;
    wire N__30989;
    wire N__30988;
    wire N__30987;
    wire N__30984;
    wire N__30983;
    wire N__30982;
    wire N__30981;
    wire N__30980;
    wire N__30979;
    wire N__30978;
    wire N__30977;
    wire N__30972;
    wire N__30971;
    wire N__30968;
    wire N__30965;
    wire N__30962;
    wire N__30961;
    wire N__30958;
    wire N__30957;
    wire N__30956;
    wire N__30953;
    wire N__30950;
    wire N__30947;
    wire N__30946;
    wire N__30945;
    wire N__30942;
    wire N__30941;
    wire N__30938;
    wire N__30935;
    wire N__30932;
    wire N__30931;
    wire N__30928;
    wire N__30925;
    wire N__30922;
    wire N__30915;
    wire N__30912;
    wire N__30911;
    wire N__30910;
    wire N__30907;
    wire N__30904;
    wire N__30901;
    wire N__30894;
    wire N__30889;
    wire N__30882;
    wire N__30879;
    wire N__30876;
    wire N__30875;
    wire N__30874;
    wire N__30869;
    wire N__30862;
    wire N__30861;
    wire N__30860;
    wire N__30857;
    wire N__30854;
    wire N__30849;
    wire N__30846;
    wire N__30843;
    wire N__30840;
    wire N__30837;
    wire N__30834;
    wire N__30831;
    wire N__30828;
    wire N__30825;
    wire N__30820;
    wire N__30811;
    wire N__30806;
    wire N__30799;
    wire N__30792;
    wire N__30787;
    wire N__30780;
    wire N__30777;
    wire N__30770;
    wire N__30769;
    wire N__30768;
    wire N__30765;
    wire N__30762;
    wire N__30761;
    wire N__30758;
    wire N__30755;
    wire N__30752;
    wire N__30749;
    wire N__30746;
    wire N__30743;
    wire N__30738;
    wire N__30733;
    wire N__30728;
    wire N__30725;
    wire N__30724;
    wire N__30723;
    wire N__30720;
    wire N__30717;
    wire N__30714;
    wire N__30709;
    wire N__30704;
    wire N__30701;
    wire N__30698;
    wire N__30695;
    wire N__30692;
    wire N__30691;
    wire N__30690;
    wire N__30687;
    wire N__30684;
    wire N__30681;
    wire N__30674;
    wire N__30671;
    wire N__30670;
    wire N__30669;
    wire N__30664;
    wire N__30661;
    wire N__30658;
    wire N__30657;
    wire N__30654;
    wire N__30651;
    wire N__30648;
    wire N__30645;
    wire N__30638;
    wire N__30635;
    wire N__30632;
    wire N__30629;
    wire N__30628;
    wire N__30627;
    wire N__30626;
    wire N__30625;
    wire N__30624;
    wire N__30623;
    wire N__30622;
    wire N__30615;
    wire N__30614;
    wire N__30613;
    wire N__30612;
    wire N__30611;
    wire N__30610;
    wire N__30609;
    wire N__30608;
    wire N__30607;
    wire N__30606;
    wire N__30601;
    wire N__30594;
    wire N__30591;
    wire N__30584;
    wire N__30577;
    wire N__30570;
    wire N__30557;
    wire N__30556;
    wire N__30555;
    wire N__30554;
    wire N__30553;
    wire N__30552;
    wire N__30549;
    wire N__30546;
    wire N__30543;
    wire N__30540;
    wire N__30537;
    wire N__30534;
    wire N__30531;
    wire N__30528;
    wire N__30525;
    wire N__30522;
    wire N__30517;
    wire N__30512;
    wire N__30503;
    wire N__30500;
    wire N__30497;
    wire N__30494;
    wire N__30493;
    wire N__30492;
    wire N__30491;
    wire N__30488;
    wire N__30485;
    wire N__30480;
    wire N__30473;
    wire N__30472;
    wire N__30471;
    wire N__30468;
    wire N__30467;
    wire N__30466;
    wire N__30463;
    wire N__30460;
    wire N__30457;
    wire N__30452;
    wire N__30449;
    wire N__30446;
    wire N__30443;
    wire N__30434;
    wire N__30433;
    wire N__30430;
    wire N__30427;
    wire N__30426;
    wire N__30423;
    wire N__30422;
    wire N__30421;
    wire N__30420;
    wire N__30419;
    wire N__30418;
    wire N__30417;
    wire N__30416;
    wire N__30413;
    wire N__30412;
    wire N__30411;
    wire N__30408;
    wire N__30405;
    wire N__30402;
    wire N__30397;
    wire N__30390;
    wire N__30387;
    wire N__30384;
    wire N__30383;
    wire N__30380;
    wire N__30379;
    wire N__30378;
    wire N__30377;
    wire N__30376;
    wire N__30375;
    wire N__30372;
    wire N__30371;
    wire N__30368;
    wire N__30361;
    wire N__30358;
    wire N__30355;
    wire N__30352;
    wire N__30343;
    wire N__30338;
    wire N__30335;
    wire N__30330;
    wire N__30321;
    wire N__30308;
    wire N__30305;
    wire N__30304;
    wire N__30303;
    wire N__30302;
    wire N__30299;
    wire N__30294;
    wire N__30291;
    wire N__30286;
    wire N__30281;
    wire N__30278;
    wire N__30277;
    wire N__30274;
    wire N__30271;
    wire N__30268;
    wire N__30265;
    wire N__30260;
    wire N__30257;
    wire N__30254;
    wire N__30251;
    wire N__30248;
    wire N__30245;
    wire N__30244;
    wire N__30243;
    wire N__30240;
    wire N__30237;
    wire N__30234;
    wire N__30233;
    wire N__30232;
    wire N__30227;
    wire N__30224;
    wire N__30221;
    wire N__30218;
    wire N__30217;
    wire N__30214;
    wire N__30211;
    wire N__30208;
    wire N__30205;
    wire N__30202;
    wire N__30191;
    wire N__30188;
    wire N__30185;
    wire N__30182;
    wire N__30179;
    wire N__30176;
    wire N__30175;
    wire N__30172;
    wire N__30171;
    wire N__30168;
    wire N__30165;
    wire N__30162;
    wire N__30159;
    wire N__30158;
    wire N__30153;
    wire N__30150;
    wire N__30147;
    wire N__30144;
    wire N__30137;
    wire N__30136;
    wire N__30133;
    wire N__30132;
    wire N__30129;
    wire N__30126;
    wire N__30123;
    wire N__30120;
    wire N__30115;
    wire N__30110;
    wire N__30109;
    wire N__30106;
    wire N__30103;
    wire N__30100;
    wire N__30095;
    wire N__30092;
    wire N__30089;
    wire N__30086;
    wire N__30083;
    wire N__30080;
    wire N__30077;
    wire N__30074;
    wire N__30071;
    wire N__30068;
    wire N__30065;
    wire N__30062;
    wire N__30059;
    wire N__30056;
    wire N__30053;
    wire N__30050;
    wire N__30047;
    wire N__30044;
    wire N__30041;
    wire N__30038;
    wire N__30035;
    wire N__30034;
    wire N__30031;
    wire N__30028;
    wire N__30025;
    wire N__30020;
    wire N__30017;
    wire N__30014;
    wire N__30011;
    wire N__30008;
    wire N__30005;
    wire N__30004;
    wire N__30003;
    wire N__30000;
    wire N__29997;
    wire N__29994;
    wire N__29989;
    wire N__29988;
    wire N__29987;
    wire N__29984;
    wire N__29981;
    wire N__29978;
    wire N__29975;
    wire N__29966;
    wire N__29965;
    wire N__29964;
    wire N__29961;
    wire N__29956;
    wire N__29953;
    wire N__29950;
    wire N__29949;
    wire N__29948;
    wire N__29945;
    wire N__29942;
    wire N__29939;
    wire N__29936;
    wire N__29927;
    wire N__29926;
    wire N__29925;
    wire N__29922;
    wire N__29919;
    wire N__29916;
    wire N__29913;
    wire N__29910;
    wire N__29909;
    wire N__29906;
    wire N__29903;
    wire N__29900;
    wire N__29899;
    wire N__29896;
    wire N__29891;
    wire N__29888;
    wire N__29885;
    wire N__29882;
    wire N__29873;
    wire N__29870;
    wire N__29867;
    wire N__29864;
    wire N__29863;
    wire N__29860;
    wire N__29857;
    wire N__29852;
    wire N__29849;
    wire N__29846;
    wire N__29843;
    wire N__29840;
    wire N__29839;
    wire N__29838;
    wire N__29837;
    wire N__29834;
    wire N__29831;
    wire N__29828;
    wire N__29825;
    wire N__29822;
    wire N__29819;
    wire N__29814;
    wire N__29811;
    wire N__29806;
    wire N__29801;
    wire N__29798;
    wire N__29795;
    wire N__29792;
    wire N__29789;
    wire N__29786;
    wire N__29783;
    wire N__29780;
    wire N__29777;
    wire N__29774;
    wire N__29771;
    wire N__29768;
    wire N__29765;
    wire N__29762;
    wire N__29759;
    wire N__29756;
    wire N__29753;
    wire N__29750;
    wire N__29747;
    wire N__29744;
    wire N__29741;
    wire N__29738;
    wire N__29737;
    wire N__29736;
    wire N__29733;
    wire N__29730;
    wire N__29727;
    wire N__29726;
    wire N__29725;
    wire N__29718;
    wire N__29715;
    wire N__29712;
    wire N__29709;
    wire N__29702;
    wire N__29701;
    wire N__29698;
    wire N__29695;
    wire N__29692;
    wire N__29691;
    wire N__29688;
    wire N__29685;
    wire N__29682;
    wire N__29675;
    wire N__29674;
    wire N__29671;
    wire N__29668;
    wire N__29665;
    wire N__29664;
    wire N__29661;
    wire N__29658;
    wire N__29655;
    wire N__29648;
    wire N__29645;
    wire N__29642;
    wire N__29639;
    wire N__29636;
    wire N__29635;
    wire N__29634;
    wire N__29633;
    wire N__29630;
    wire N__29627;
    wire N__29622;
    wire N__29619;
    wire N__29616;
    wire N__29615;
    wire N__29612;
    wire N__29609;
    wire N__29606;
    wire N__29603;
    wire N__29600;
    wire N__29591;
    wire N__29590;
    wire N__29589;
    wire N__29586;
    wire N__29583;
    wire N__29580;
    wire N__29577;
    wire N__29574;
    wire N__29571;
    wire N__29566;
    wire N__29561;
    wire N__29560;
    wire N__29559;
    wire N__29556;
    wire N__29553;
    wire N__29552;
    wire N__29551;
    wire N__29548;
    wire N__29545;
    wire N__29542;
    wire N__29539;
    wire N__29536;
    wire N__29533;
    wire N__29530;
    wire N__29525;
    wire N__29522;
    wire N__29513;
    wire N__29512;
    wire N__29509;
    wire N__29506;
    wire N__29505;
    wire N__29502;
    wire N__29499;
    wire N__29496;
    wire N__29493;
    wire N__29486;
    wire N__29485;
    wire N__29484;
    wire N__29481;
    wire N__29478;
    wire N__29475;
    wire N__29474;
    wire N__29469;
    wire N__29466;
    wire N__29465;
    wire N__29462;
    wire N__29457;
    wire N__29454;
    wire N__29451;
    wire N__29444;
    wire N__29443;
    wire N__29442;
    wire N__29439;
    wire N__29436;
    wire N__29433;
    wire N__29426;
    wire N__29425;
    wire N__29424;
    wire N__29421;
    wire N__29418;
    wire N__29415;
    wire N__29412;
    wire N__29409;
    wire N__29406;
    wire N__29401;
    wire N__29396;
    wire N__29395;
    wire N__29392;
    wire N__29391;
    wire N__29390;
    wire N__29387;
    wire N__29386;
    wire N__29383;
    wire N__29380;
    wire N__29375;
    wire N__29372;
    wire N__29369;
    wire N__29366;
    wire N__29363;
    wire N__29360;
    wire N__29351;
    wire N__29350;
    wire N__29349;
    wire N__29346;
    wire N__29343;
    wire N__29340;
    wire N__29337;
    wire N__29334;
    wire N__29331;
    wire N__29326;
    wire N__29321;
    wire N__29320;
    wire N__29319;
    wire N__29316;
    wire N__29313;
    wire N__29310;
    wire N__29307;
    wire N__29304;
    wire N__29301;
    wire N__29298;
    wire N__29291;
    wire N__29290;
    wire N__29287;
    wire N__29286;
    wire N__29283;
    wire N__29280;
    wire N__29277;
    wire N__29274;
    wire N__29271;
    wire N__29268;
    wire N__29265;
    wire N__29258;
    wire N__29257;
    wire N__29256;
    wire N__29253;
    wire N__29250;
    wire N__29247;
    wire N__29246;
    wire N__29245;
    wire N__29240;
    wire N__29237;
    wire N__29234;
    wire N__29231;
    wire N__29228;
    wire N__29225;
    wire N__29220;
    wire N__29213;
    wire N__29212;
    wire N__29209;
    wire N__29208;
    wire N__29205;
    wire N__29202;
    wire N__29199;
    wire N__29196;
    wire N__29193;
    wire N__29190;
    wire N__29187;
    wire N__29180;
    wire N__29177;
    wire N__29174;
    wire N__29171;
    wire N__29168;
    wire N__29165;
    wire N__29162;
    wire N__29159;
    wire N__29158;
    wire N__29157;
    wire N__29154;
    wire N__29153;
    wire N__29150;
    wire N__29147;
    wire N__29144;
    wire N__29141;
    wire N__29138;
    wire N__29135;
    wire N__29130;
    wire N__29127;
    wire N__29120;
    wire N__29117;
    wire N__29114;
    wire N__29111;
    wire N__29108;
    wire N__29105;
    wire N__29102;
    wire N__29101;
    wire N__29098;
    wire N__29097;
    wire N__29094;
    wire N__29091;
    wire N__29090;
    wire N__29087;
    wire N__29084;
    wire N__29081;
    wire N__29078;
    wire N__29073;
    wire N__29066;
    wire N__29065;
    wire N__29062;
    wire N__29061;
    wire N__29060;
    wire N__29057;
    wire N__29054;
    wire N__29049;
    wire N__29046;
    wire N__29045;
    wire N__29042;
    wire N__29039;
    wire N__29036;
    wire N__29033;
    wire N__29024;
    wire N__29023;
    wire N__29022;
    wire N__29019;
    wire N__29016;
    wire N__29013;
    wire N__29010;
    wire N__29007;
    wire N__29004;
    wire N__29001;
    wire N__28994;
    wire N__28991;
    wire N__28990;
    wire N__28987;
    wire N__28984;
    wire N__28983;
    wire N__28982;
    wire N__28977;
    wire N__28972;
    wire N__28971;
    wire N__28968;
    wire N__28965;
    wire N__28962;
    wire N__28959;
    wire N__28952;
    wire N__28951;
    wire N__28948;
    wire N__28945;
    wire N__28944;
    wire N__28941;
    wire N__28938;
    wire N__28935;
    wire N__28932;
    wire N__28929;
    wire N__28926;
    wire N__28923;
    wire N__28916;
    wire N__28915;
    wire N__28912;
    wire N__28911;
    wire N__28908;
    wire N__28905;
    wire N__28902;
    wire N__28899;
    wire N__28896;
    wire N__28893;
    wire N__28890;
    wire N__28883;
    wire N__28882;
    wire N__28881;
    wire N__28878;
    wire N__28875;
    wire N__28872;
    wire N__28869;
    wire N__28866;
    wire N__28863;
    wire N__28860;
    wire N__28853;
    wire N__28852;
    wire N__28849;
    wire N__28846;
    wire N__28841;
    wire N__28840;
    wire N__28839;
    wire N__28836;
    wire N__28833;
    wire N__28830;
    wire N__28823;
    wire N__28820;
    wire N__28817;
    wire N__28814;
    wire N__28813;
    wire N__28810;
    wire N__28807;
    wire N__28802;
    wire N__28799;
    wire N__28796;
    wire N__28795;
    wire N__28792;
    wire N__28789;
    wire N__28784;
    wire N__28783;
    wire N__28780;
    wire N__28779;
    wire N__28776;
    wire N__28773;
    wire N__28770;
    wire N__28767;
    wire N__28764;
    wire N__28761;
    wire N__28760;
    wire N__28757;
    wire N__28752;
    wire N__28751;
    wire N__28748;
    wire N__28745;
    wire N__28742;
    wire N__28739;
    wire N__28736;
    wire N__28727;
    wire N__28726;
    wire N__28723;
    wire N__28720;
    wire N__28717;
    wire N__28712;
    wire N__28709;
    wire N__28708;
    wire N__28707;
    wire N__28704;
    wire N__28699;
    wire N__28694;
    wire N__28693;
    wire N__28692;
    wire N__28689;
    wire N__28684;
    wire N__28679;
    wire N__28676;
    wire N__28675;
    wire N__28672;
    wire N__28671;
    wire N__28668;
    wire N__28663;
    wire N__28658;
    wire N__28655;
    wire N__28654;
    wire N__28653;
    wire N__28652;
    wire N__28647;
    wire N__28642;
    wire N__28637;
    wire N__28634;
    wire N__28633;
    wire N__28632;
    wire N__28629;
    wire N__28624;
    wire N__28619;
    wire N__28616;
    wire N__28615;
    wire N__28614;
    wire N__28611;
    wire N__28610;
    wire N__28607;
    wire N__28604;
    wire N__28601;
    wire N__28598;
    wire N__28589;
    wire N__28588;
    wire N__28585;
    wire N__28584;
    wire N__28581;
    wire N__28578;
    wire N__28575;
    wire N__28574;
    wire N__28571;
    wire N__28566;
    wire N__28563;
    wire N__28558;
    wire N__28553;
    wire N__28550;
    wire N__28547;
    wire N__28546;
    wire N__28543;
    wire N__28540;
    wire N__28537;
    wire N__28534;
    wire N__28529;
    wire N__28526;
    wire N__28525;
    wire N__28522;
    wire N__28521;
    wire N__28518;
    wire N__28515;
    wire N__28514;
    wire N__28511;
    wire N__28508;
    wire N__28505;
    wire N__28502;
    wire N__28497;
    wire N__28490;
    wire N__28487;
    wire N__28484;
    wire N__28481;
    wire N__28480;
    wire N__28477;
    wire N__28474;
    wire N__28469;
    wire N__28466;
    wire N__28463;
    wire N__28460;
    wire N__28457;
    wire N__28454;
    wire N__28453;
    wire N__28452;
    wire N__28449;
    wire N__28446;
    wire N__28441;
    wire N__28436;
    wire N__28433;
    wire N__28430;
    wire N__28427;
    wire N__28426;
    wire N__28425;
    wire N__28422;
    wire N__28419;
    wire N__28418;
    wire N__28409;
    wire N__28406;
    wire N__28405;
    wire N__28402;
    wire N__28399;
    wire N__28396;
    wire N__28393;
    wire N__28390;
    wire N__28385;
    wire N__28384;
    wire N__28381;
    wire N__28378;
    wire N__28375;
    wire N__28372;
    wire N__28369;
    wire N__28364;
    wire N__28361;
    wire N__28358;
    wire N__28355;
    wire N__28352;
    wire N__28349;
    wire N__28346;
    wire N__28343;
    wire N__28340;
    wire N__28339;
    wire N__28338;
    wire N__28337;
    wire N__28334;
    wire N__28333;
    wire N__28332;
    wire N__28331;
    wire N__28328;
    wire N__28325;
    wire N__28322;
    wire N__28319;
    wire N__28314;
    wire N__28313;
    wire N__28310;
    wire N__28307;
    wire N__28304;
    wire N__28301;
    wire N__28298;
    wire N__28297;
    wire N__28294;
    wire N__28293;
    wire N__28290;
    wire N__28287;
    wire N__28282;
    wire N__28277;
    wire N__28274;
    wire N__28271;
    wire N__28268;
    wire N__28253;
    wire N__28252;
    wire N__28249;
    wire N__28246;
    wire N__28243;
    wire N__28240;
    wire N__28239;
    wire N__28238;
    wire N__28235;
    wire N__28234;
    wire N__28233;
    wire N__28230;
    wire N__28225;
    wire N__28222;
    wire N__28217;
    wire N__28208;
    wire N__28207;
    wire N__28206;
    wire N__28205;
    wire N__28204;
    wire N__28203;
    wire N__28202;
    wire N__28201;
    wire N__28198;
    wire N__28197;
    wire N__28192;
    wire N__28189;
    wire N__28186;
    wire N__28185;
    wire N__28184;
    wire N__28183;
    wire N__28178;
    wire N__28175;
    wire N__28174;
    wire N__28173;
    wire N__28170;
    wire N__28167;
    wire N__28164;
    wire N__28161;
    wire N__28158;
    wire N__28151;
    wire N__28148;
    wire N__28145;
    wire N__28142;
    wire N__28139;
    wire N__28138;
    wire N__28137;
    wire N__28136;
    wire N__28133;
    wire N__28130;
    wire N__28127;
    wire N__28116;
    wire N__28113;
    wire N__28110;
    wire N__28107;
    wire N__28102;
    wire N__28099;
    wire N__28096;
    wire N__28091;
    wire N__28076;
    wire N__28073;
    wire N__28070;
    wire N__28067;
    wire N__28066;
    wire N__28065;
    wire N__28064;
    wire N__28061;
    wire N__28058;
    wire N__28053;
    wire N__28050;
    wire N__28047;
    wire N__28046;
    wire N__28045;
    wire N__28040;
    wire N__28037;
    wire N__28032;
    wire N__28025;
    wire N__28022;
    wire N__28019;
    wire N__28016;
    wire N__28013;
    wire N__28010;
    wire N__28007;
    wire N__28004;
    wire N__28003;
    wire N__27998;
    wire N__27997;
    wire N__27994;
    wire N__27993;
    wire N__27990;
    wire N__27987;
    wire N__27984;
    wire N__27983;
    wire N__27980;
    wire N__27975;
    wire N__27972;
    wire N__27967;
    wire N__27962;
    wire N__27961;
    wire N__27960;
    wire N__27959;
    wire N__27954;
    wire N__27951;
    wire N__27950;
    wire N__27947;
    wire N__27944;
    wire N__27941;
    wire N__27938;
    wire N__27935;
    wire N__27932;
    wire N__27925;
    wire N__27920;
    wire N__27919;
    wire N__27918;
    wire N__27917;
    wire N__27914;
    wire N__27911;
    wire N__27910;
    wire N__27909;
    wire N__27902;
    wire N__27899;
    wire N__27896;
    wire N__27893;
    wire N__27890;
    wire N__27887;
    wire N__27886;
    wire N__27883;
    wire N__27880;
    wire N__27877;
    wire N__27874;
    wire N__27871;
    wire N__27866;
    wire N__27859;
    wire N__27856;
    wire N__27853;
    wire N__27850;
    wire N__27845;
    wire N__27844;
    wire N__27841;
    wire N__27840;
    wire N__27839;
    wire N__27838;
    wire N__27837;
    wire N__27834;
    wire N__27833;
    wire N__27830;
    wire N__27827;
    wire N__27822;
    wire N__27819;
    wire N__27816;
    wire N__27813;
    wire N__27808;
    wire N__27805;
    wire N__27802;
    wire N__27799;
    wire N__27796;
    wire N__27793;
    wire N__27788;
    wire N__27787;
    wire N__27782;
    wire N__27779;
    wire N__27776;
    wire N__27773;
    wire N__27768;
    wire N__27763;
    wire N__27760;
    wire N__27757;
    wire N__27754;
    wire N__27751;
    wire N__27746;
    wire N__27745;
    wire N__27742;
    wire N__27739;
    wire N__27736;
    wire N__27733;
    wire N__27728;
    wire N__27727;
    wire N__27724;
    wire N__27721;
    wire N__27718;
    wire N__27715;
    wire N__27710;
    wire N__27709;
    wire N__27706;
    wire N__27703;
    wire N__27700;
    wire N__27697;
    wire N__27692;
    wire N__27691;
    wire N__27688;
    wire N__27685;
    wire N__27682;
    wire N__27679;
    wire N__27676;
    wire N__27671;
    wire N__27670;
    wire N__27667;
    wire N__27664;
    wire N__27661;
    wire N__27658;
    wire N__27655;
    wire N__27650;
    wire N__27649;
    wire N__27646;
    wire N__27643;
    wire N__27640;
    wire N__27637;
    wire N__27632;
    wire N__27631;
    wire N__27628;
    wire N__27625;
    wire N__27622;
    wire N__27619;
    wire N__27616;
    wire N__27611;
    wire N__27610;
    wire N__27607;
    wire N__27604;
    wire N__27601;
    wire N__27598;
    wire N__27595;
    wire N__27590;
    wire N__27587;
    wire N__27586;
    wire N__27585;
    wire N__27582;
    wire N__27579;
    wire N__27576;
    wire N__27575;
    wire N__27572;
    wire N__27569;
    wire N__27566;
    wire N__27563;
    wire N__27562;
    wire N__27559;
    wire N__27552;
    wire N__27549;
    wire N__27542;
    wire N__27539;
    wire N__27536;
    wire N__27533;
    wire N__27530;
    wire N__27527;
    wire N__27524;
    wire N__27521;
    wire N__27520;
    wire N__27517;
    wire N__27514;
    wire N__27511;
    wire N__27506;
    wire N__27505;
    wire N__27502;
    wire N__27499;
    wire N__27496;
    wire N__27493;
    wire N__27488;
    wire N__27487;
    wire N__27486;
    wire N__27483;
    wire N__27480;
    wire N__27479;
    wire N__27476;
    wire N__27471;
    wire N__27468;
    wire N__27465;
    wire N__27460;
    wire N__27455;
    wire N__27452;
    wire N__27449;
    wire N__27448;
    wire N__27445;
    wire N__27442;
    wire N__27441;
    wire N__27438;
    wire N__27435;
    wire N__27434;
    wire N__27431;
    wire N__27430;
    wire N__27425;
    wire N__27422;
    wire N__27419;
    wire N__27416;
    wire N__27413;
    wire N__27410;
    wire N__27405;
    wire N__27398;
    wire N__27395;
    wire N__27394;
    wire N__27393;
    wire N__27390;
    wire N__27387;
    wire N__27384;
    wire N__27383;
    wire N__27380;
    wire N__27377;
    wire N__27374;
    wire N__27371;
    wire N__27370;
    wire N__27365;
    wire N__27360;
    wire N__27357;
    wire N__27350;
    wire N__27349;
    wire N__27348;
    wire N__27345;
    wire N__27342;
    wire N__27339;
    wire N__27336;
    wire N__27333;
    wire N__27330;
    wire N__27327;
    wire N__27324;
    wire N__27321;
    wire N__27320;
    wire N__27319;
    wire N__27312;
    wire N__27309;
    wire N__27306;
    wire N__27299;
    wire N__27296;
    wire N__27293;
    wire N__27290;
    wire N__27287;
    wire N__27284;
    wire N__27283;
    wire N__27280;
    wire N__27277;
    wire N__27276;
    wire N__27271;
    wire N__27270;
    wire N__27267;
    wire N__27264;
    wire N__27261;
    wire N__27254;
    wire N__27251;
    wire N__27250;
    wire N__27249;
    wire N__27248;
    wire N__27245;
    wire N__27242;
    wire N__27239;
    wire N__27236;
    wire N__27233;
    wire N__27228;
    wire N__27225;
    wire N__27222;
    wire N__27217;
    wire N__27214;
    wire N__27211;
    wire N__27206;
    wire N__27205;
    wire N__27204;
    wire N__27203;
    wire N__27200;
    wire N__27197;
    wire N__27196;
    wire N__27193;
    wire N__27192;
    wire N__27191;
    wire N__27190;
    wire N__27189;
    wire N__27188;
    wire N__27183;
    wire N__27182;
    wire N__27179;
    wire N__27174;
    wire N__27171;
    wire N__27168;
    wire N__27163;
    wire N__27162;
    wire N__27159;
    wire N__27156;
    wire N__27153;
    wire N__27150;
    wire N__27147;
    wire N__27146;
    wire N__27143;
    wire N__27138;
    wire N__27133;
    wire N__27130;
    wire N__27127;
    wire N__27122;
    wire N__27119;
    wire N__27104;
    wire N__27101;
    wire N__27098;
    wire N__27097;
    wire N__27094;
    wire N__27091;
    wire N__27086;
    wire N__27083;
    wire N__27080;
    wire N__27077;
    wire N__27074;
    wire N__27073;
    wire N__27070;
    wire N__27067;
    wire N__27062;
    wire N__27059;
    wire N__27058;
    wire N__27055;
    wire N__27052;
    wire N__27049;
    wire N__27046;
    wire N__27043;
    wire N__27040;
    wire N__27035;
    wire N__27032;
    wire N__27029;
    wire N__27026;
    wire N__27023;
    wire N__27022;
    wire N__27019;
    wire N__27018;
    wire N__27015;
    wire N__27012;
    wire N__27009;
    wire N__27006;
    wire N__26999;
    wire N__26998;
    wire N__26995;
    wire N__26992;
    wire N__26987;
    wire N__26986;
    wire N__26983;
    wire N__26982;
    wire N__26979;
    wire N__26976;
    wire N__26971;
    wire N__26966;
    wire N__26965;
    wire N__26962;
    wire N__26959;
    wire N__26954;
    wire N__26951;
    wire N__26950;
    wire N__26947;
    wire N__26944;
    wire N__26941;
    wire N__26938;
    wire N__26935;
    wire N__26934;
    wire N__26929;
    wire N__26926;
    wire N__26921;
    wire N__26918;
    wire N__26915;
    wire N__26912;
    wire N__26909;
    wire N__26906;
    wire N__26903;
    wire N__26902;
    wire N__26901;
    wire N__26900;
    wire N__26899;
    wire N__26898;
    wire N__26897;
    wire N__26894;
    wire N__26891;
    wire N__26886;
    wire N__26885;
    wire N__26884;
    wire N__26883;
    wire N__26882;
    wire N__26881;
    wire N__26878;
    wire N__26875;
    wire N__26874;
    wire N__26871;
    wire N__26866;
    wire N__26863;
    wire N__26856;
    wire N__26851;
    wire N__26848;
    wire N__26845;
    wire N__26842;
    wire N__26837;
    wire N__26828;
    wire N__26819;
    wire N__26816;
    wire N__26813;
    wire N__26810;
    wire N__26807;
    wire N__26804;
    wire N__26801;
    wire N__26800;
    wire N__26797;
    wire N__26796;
    wire N__26793;
    wire N__26790;
    wire N__26785;
    wire N__26780;
    wire N__26777;
    wire N__26774;
    wire N__26773;
    wire N__26770;
    wire N__26767;
    wire N__26762;
    wire N__26761;
    wire N__26758;
    wire N__26755;
    wire N__26752;
    wire N__26749;
    wire N__26744;
    wire N__26741;
    wire N__26738;
    wire N__26737;
    wire N__26734;
    wire N__26731;
    wire N__26728;
    wire N__26725;
    wire N__26720;
    wire N__26717;
    wire N__26716;
    wire N__26713;
    wire N__26712;
    wire N__26709;
    wire N__26706;
    wire N__26703;
    wire N__26700;
    wire N__26697;
    wire N__26690;
    wire N__26689;
    wire N__26686;
    wire N__26683;
    wire N__26678;
    wire N__26675;
    wire N__26674;
    wire N__26671;
    wire N__26668;
    wire N__26665;
    wire N__26660;
    wire N__26657;
    wire N__26654;
    wire N__26651;
    wire N__26648;
    wire N__26647;
    wire N__26644;
    wire N__26641;
    wire N__26638;
    wire N__26635;
    wire N__26630;
    wire N__26627;
    wire N__26624;
    wire N__26621;
    wire N__26618;
    wire N__26617;
    wire N__26614;
    wire N__26611;
    wire N__26608;
    wire N__26603;
    wire N__26600;
    wire N__26597;
    wire N__26594;
    wire N__26591;
    wire N__26590;
    wire N__26587;
    wire N__26584;
    wire N__26579;
    wire N__26576;
    wire N__26573;
    wire N__26570;
    wire N__26569;
    wire N__26566;
    wire N__26563;
    wire N__26558;
    wire N__26555;
    wire N__26552;
    wire N__26551;
    wire N__26548;
    wire N__26545;
    wire N__26540;
    wire N__26537;
    wire N__26534;
    wire N__26531;
    wire N__26528;
    wire N__26527;
    wire N__26526;
    wire N__26525;
    wire N__26524;
    wire N__26523;
    wire N__26522;
    wire N__26521;
    wire N__26520;
    wire N__26519;
    wire N__26518;
    wire N__26503;
    wire N__26500;
    wire N__26493;
    wire N__26490;
    wire N__26485;
    wire N__26482;
    wire N__26479;
    wire N__26476;
    wire N__26473;
    wire N__26470;
    wire N__26467;
    wire N__26462;
    wire N__26459;
    wire N__26458;
    wire N__26455;
    wire N__26452;
    wire N__26451;
    wire N__26450;
    wire N__26449;
    wire N__26446;
    wire N__26443;
    wire N__26442;
    wire N__26441;
    wire N__26436;
    wire N__26433;
    wire N__26430;
    wire N__26427;
    wire N__26422;
    wire N__26417;
    wire N__26408;
    wire N__26405;
    wire N__26402;
    wire N__26399;
    wire N__26396;
    wire N__26393;
    wire N__26390;
    wire N__26387;
    wire N__26384;
    wire N__26381;
    wire N__26378;
    wire N__26375;
    wire N__26372;
    wire N__26369;
    wire N__26366;
    wire N__26363;
    wire N__26360;
    wire N__26357;
    wire N__26354;
    wire N__26351;
    wire N__26348;
    wire N__26345;
    wire N__26342;
    wire N__26339;
    wire N__26336;
    wire N__26333;
    wire N__26330;
    wire N__26327;
    wire N__26324;
    wire N__26321;
    wire N__26318;
    wire N__26315;
    wire N__26312;
    wire N__26309;
    wire N__26306;
    wire N__26303;
    wire N__26300;
    wire N__26297;
    wire N__26294;
    wire N__26291;
    wire N__26288;
    wire N__26285;
    wire N__26282;
    wire N__26279;
    wire N__26276;
    wire N__26273;
    wire N__26270;
    wire N__26267;
    wire N__26264;
    wire N__26261;
    wire N__26260;
    wire N__26257;
    wire N__26254;
    wire N__26251;
    wire N__26248;
    wire N__26245;
    wire N__26242;
    wire N__26239;
    wire N__26236;
    wire N__26233;
    wire N__26230;
    wire N__26225;
    wire N__26222;
    wire N__26221;
    wire N__26218;
    wire N__26215;
    wire N__26210;
    wire N__26207;
    wire N__26206;
    wire N__26205;
    wire N__26202;
    wire N__26199;
    wire N__26198;
    wire N__26197;
    wire N__26194;
    wire N__26191;
    wire N__26190;
    wire N__26187;
    wire N__26184;
    wire N__26181;
    wire N__26180;
    wire N__26177;
    wire N__26174;
    wire N__26171;
    wire N__26168;
    wire N__26163;
    wire N__26160;
    wire N__26153;
    wire N__26150;
    wire N__26145;
    wire N__26144;
    wire N__26141;
    wire N__26136;
    wire N__26133;
    wire N__26130;
    wire N__26127;
    wire N__26124;
    wire N__26121;
    wire N__26116;
    wire N__26111;
    wire N__26108;
    wire N__26105;
    wire N__26102;
    wire N__26099;
    wire N__26096;
    wire N__26093;
    wire N__26090;
    wire N__26087;
    wire N__26084;
    wire N__26081;
    wire N__26078;
    wire N__26075;
    wire N__26074;
    wire N__26071;
    wire N__26068;
    wire N__26067;
    wire N__26062;
    wire N__26061;
    wire N__26060;
    wire N__26057;
    wire N__26054;
    wire N__26051;
    wire N__26048;
    wire N__26045;
    wire N__26042;
    wire N__26033;
    wire N__26032;
    wire N__26031;
    wire N__26028;
    wire N__26025;
    wire N__26022;
    wire N__26021;
    wire N__26018;
    wire N__26015;
    wire N__26014;
    wire N__26011;
    wire N__26008;
    wire N__26005;
    wire N__26004;
    wire N__26001;
    wire N__25998;
    wire N__25995;
    wire N__25992;
    wire N__25989;
    wire N__25986;
    wire N__25981;
    wire N__25978;
    wire N__25975;
    wire N__25970;
    wire N__25963;
    wire N__25958;
    wire N__25957;
    wire N__25956;
    wire N__25955;
    wire N__25954;
    wire N__25953;
    wire N__25952;
    wire N__25951;
    wire N__25942;
    wire N__25939;
    wire N__25936;
    wire N__25935;
    wire N__25934;
    wire N__25933;
    wire N__25930;
    wire N__25927;
    wire N__25922;
    wire N__25919;
    wire N__25916;
    wire N__25913;
    wire N__25912;
    wire N__25911;
    wire N__25910;
    wire N__25909;
    wire N__25906;
    wire N__25903;
    wire N__25900;
    wire N__25899;
    wire N__25896;
    wire N__25893;
    wire N__25890;
    wire N__25887;
    wire N__25876;
    wire N__25873;
    wire N__25870;
    wire N__25867;
    wire N__25864;
    wire N__25861;
    wire N__25858;
    wire N__25853;
    wire N__25850;
    wire N__25847;
    wire N__25844;
    wire N__25829;
    wire N__25828;
    wire N__25827;
    wire N__25824;
    wire N__25821;
    wire N__25818;
    wire N__25817;
    wire N__25816;
    wire N__25815;
    wire N__25814;
    wire N__25807;
    wire N__25804;
    wire N__25799;
    wire N__25796;
    wire N__25793;
    wire N__25784;
    wire N__25781;
    wire N__25778;
    wire N__25775;
    wire N__25774;
    wire N__25771;
    wire N__25768;
    wire N__25763;
    wire N__25760;
    wire N__25757;
    wire N__25754;
    wire N__25751;
    wire N__25748;
    wire N__25745;
    wire N__25742;
    wire N__25739;
    wire N__25738;
    wire N__25735;
    wire N__25732;
    wire N__25731;
    wire N__25728;
    wire N__25725;
    wire N__25724;
    wire N__25723;
    wire N__25722;
    wire N__25721;
    wire N__25718;
    wire N__25713;
    wire N__25708;
    wire N__25701;
    wire N__25698;
    wire N__25691;
    wire N__25688;
    wire N__25687;
    wire N__25686;
    wire N__25685;
    wire N__25682;
    wire N__25679;
    wire N__25676;
    wire N__25673;
    wire N__25672;
    wire N__25667;
    wire N__25664;
    wire N__25661;
    wire N__25658;
    wire N__25655;
    wire N__25650;
    wire N__25647;
    wire N__25640;
    wire N__25639;
    wire N__25636;
    wire N__25635;
    wire N__25634;
    wire N__25633;
    wire N__25632;
    wire N__25629;
    wire N__25628;
    wire N__25625;
    wire N__25624;
    wire N__25617;
    wire N__25614;
    wire N__25609;
    wire N__25606;
    wire N__25603;
    wire N__25598;
    wire N__25595;
    wire N__25590;
    wire N__25587;
    wire N__25584;
    wire N__25577;
    wire N__25574;
    wire N__25571;
    wire N__25568;
    wire N__25565;
    wire N__25562;
    wire N__25559;
    wire N__25556;
    wire N__25553;
    wire N__25550;
    wire N__25547;
    wire N__25544;
    wire N__25541;
    wire N__25538;
    wire N__25537;
    wire N__25532;
    wire N__25531;
    wire N__25530;
    wire N__25529;
    wire N__25528;
    wire N__25525;
    wire N__25524;
    wire N__25521;
    wire N__25516;
    wire N__25513;
    wire N__25510;
    wire N__25505;
    wire N__25502;
    wire N__25495;
    wire N__25492;
    wire N__25489;
    wire N__25484;
    wire N__25483;
    wire N__25480;
    wire N__25477;
    wire N__25474;
    wire N__25471;
    wire N__25470;
    wire N__25469;
    wire N__25464;
    wire N__25459;
    wire N__25458;
    wire N__25457;
    wire N__25454;
    wire N__25451;
    wire N__25446;
    wire N__25439;
    wire N__25438;
    wire N__25437;
    wire N__25434;
    wire N__25431;
    wire N__25428;
    wire N__25423;
    wire N__25420;
    wire N__25419;
    wire N__25418;
    wire N__25417;
    wire N__25416;
    wire N__25413;
    wire N__25410;
    wire N__25407;
    wire N__25400;
    wire N__25397;
    wire N__25388;
    wire N__25385;
    wire N__25382;
    wire N__25379;
    wire N__25376;
    wire N__25373;
    wire N__25370;
    wire N__25367;
    wire N__25366;
    wire N__25365;
    wire N__25364;
    wire N__25363;
    wire N__25360;
    wire N__25359;
    wire N__25358;
    wire N__25355;
    wire N__25350;
    wire N__25349;
    wire N__25348;
    wire N__25347;
    wire N__25344;
    wire N__25341;
    wire N__25340;
    wire N__25339;
    wire N__25336;
    wire N__25333;
    wire N__25330;
    wire N__25327;
    wire N__25324;
    wire N__25321;
    wire N__25316;
    wire N__25313;
    wire N__25308;
    wire N__25301;
    wire N__25286;
    wire N__25283;
    wire N__25280;
    wire N__25277;
    wire N__25274;
    wire N__25271;
    wire N__25268;
    wire N__25267;
    wire N__25264;
    wire N__25261;
    wire N__25260;
    wire N__25259;
    wire N__25258;
    wire N__25257;
    wire N__25256;
    wire N__25255;
    wire N__25254;
    wire N__25253;
    wire N__25250;
    wire N__25249;
    wire N__25248;
    wire N__25245;
    wire N__25242;
    wire N__25237;
    wire N__25234;
    wire N__25231;
    wire N__25228;
    wire N__25225;
    wire N__25222;
    wire N__25219;
    wire N__25214;
    wire N__25207;
    wire N__25202;
    wire N__25187;
    wire N__25184;
    wire N__25181;
    wire N__25178;
    wire N__25175;
    wire N__25172;
    wire N__25169;
    wire N__25166;
    wire N__25163;
    wire N__25160;
    wire N__25157;
    wire N__25154;
    wire N__25151;
    wire N__25148;
    wire N__25145;
    wire N__25142;
    wire N__25141;
    wire N__25138;
    wire N__25135;
    wire N__25132;
    wire N__25129;
    wire N__25126;
    wire N__25123;
    wire N__25120;
    wire N__25117;
    wire N__25112;
    wire N__25109;
    wire N__25106;
    wire N__25105;
    wire N__25102;
    wire N__25099;
    wire N__25096;
    wire N__25093;
    wire N__25088;
    wire N__25085;
    wire N__25082;
    wire N__25079;
    wire N__25076;
    wire N__25073;
    wire N__25070;
    wire N__25067;
    wire N__25064;
    wire N__25061;
    wire N__25058;
    wire N__25057;
    wire N__25054;
    wire N__25051;
    wire N__25048;
    wire N__25045;
    wire N__25042;
    wire N__25039;
    wire N__25034;
    wire N__25031;
    wire N__25028;
    wire N__25025;
    wire N__25022;
    wire N__25019;
    wire N__25016;
    wire N__25013;
    wire N__25010;
    wire N__25009;
    wire N__25006;
    wire N__25003;
    wire N__25000;
    wire N__24995;
    wire N__24992;
    wire N__24989;
    wire N__24986;
    wire N__24983;
    wire N__24980;
    wire N__24977;
    wire N__24976;
    wire N__24973;
    wire N__24970;
    wire N__24967;
    wire N__24964;
    wire N__24961;
    wire N__24958;
    wire N__24955;
    wire N__24952;
    wire N__24947;
    wire N__24944;
    wire N__24943;
    wire N__24940;
    wire N__24937;
    wire N__24932;
    wire N__24929;
    wire N__24926;
    wire N__24923;
    wire N__24920;
    wire N__24917;
    wire N__24914;
    wire N__24911;
    wire N__24908;
    wire N__24907;
    wire N__24904;
    wire N__24901;
    wire N__24898;
    wire N__24893;
    wire N__24890;
    wire N__24887;
    wire N__24884;
    wire N__24881;
    wire N__24880;
    wire N__24877;
    wire N__24874;
    wire N__24871;
    wire N__24866;
    wire N__24863;
    wire N__24860;
    wire N__24857;
    wire N__24854;
    wire N__24851;
    wire N__24848;
    wire N__24845;
    wire N__24842;
    wire N__24839;
    wire N__24836;
    wire N__24835;
    wire N__24832;
    wire N__24829;
    wire N__24826;
    wire N__24823;
    wire N__24820;
    wire N__24815;
    wire N__24812;
    wire N__24809;
    wire N__24806;
    wire N__24803;
    wire N__24800;
    wire N__24797;
    wire N__24794;
    wire N__24791;
    wire N__24790;
    wire N__24787;
    wire N__24784;
    wire N__24779;
    wire N__24776;
    wire N__24773;
    wire N__24770;
    wire N__24767;
    wire N__24764;
    wire N__24763;
    wire N__24760;
    wire N__24757;
    wire N__24754;
    wire N__24751;
    wire N__24746;
    wire N__24743;
    wire N__24740;
    wire N__24737;
    wire N__24734;
    wire N__24731;
    wire N__24728;
    wire N__24727;
    wire N__24724;
    wire N__24721;
    wire N__24718;
    wire N__24715;
    wire N__24710;
    wire N__24707;
    wire N__24704;
    wire N__24701;
    wire N__24698;
    wire N__24695;
    wire N__24692;
    wire N__24689;
    wire N__24686;
    wire N__24683;
    wire N__24680;
    wire N__24677;
    wire N__24674;
    wire N__24671;
    wire N__24668;
    wire N__24665;
    wire N__24662;
    wire N__24661;
    wire N__24660;
    wire N__24659;
    wire N__24658;
    wire N__24653;
    wire N__24650;
    wire N__24647;
    wire N__24644;
    wire N__24639;
    wire N__24634;
    wire N__24629;
    wire N__24626;
    wire N__24623;
    wire N__24620;
    wire N__24617;
    wire N__24614;
    wire N__24611;
    wire N__24608;
    wire N__24605;
    wire N__24602;
    wire N__24599;
    wire N__24596;
    wire N__24593;
    wire N__24592;
    wire N__24591;
    wire N__24590;
    wire N__24587;
    wire N__24584;
    wire N__24581;
    wire N__24578;
    wire N__24575;
    wire N__24570;
    wire N__24567;
    wire N__24560;
    wire N__24559;
    wire N__24558;
    wire N__24551;
    wire N__24550;
    wire N__24549;
    wire N__24548;
    wire N__24545;
    wire N__24540;
    wire N__24537;
    wire N__24530;
    wire N__24527;
    wire N__24524;
    wire N__24523;
    wire N__24522;
    wire N__24521;
    wire N__24516;
    wire N__24515;
    wire N__24514;
    wire N__24513;
    wire N__24508;
    wire N__24505;
    wire N__24500;
    wire N__24497;
    wire N__24488;
    wire N__24487;
    wire N__24484;
    wire N__24481;
    wire N__24478;
    wire N__24477;
    wire N__24476;
    wire N__24475;
    wire N__24470;
    wire N__24467;
    wire N__24466;
    wire N__24463;
    wire N__24460;
    wire N__24457;
    wire N__24452;
    wire N__24449;
    wire N__24446;
    wire N__24437;
    wire N__24434;
    wire N__24431;
    wire N__24428;
    wire N__24425;
    wire N__24422;
    wire N__24421;
    wire N__24418;
    wire N__24415;
    wire N__24412;
    wire N__24409;
    wire N__24404;
    wire N__24401;
    wire N__24398;
    wire N__24395;
    wire N__24392;
    wire N__24389;
    wire N__24388;
    wire N__24385;
    wire N__24382;
    wire N__24379;
    wire N__24376;
    wire N__24371;
    wire N__24368;
    wire N__24365;
    wire N__24362;
    wire N__24359;
    wire N__24356;
    wire N__24353;
    wire N__24350;
    wire N__24347;
    wire N__24344;
    wire N__24343;
    wire N__24340;
    wire N__24335;
    wire N__24332;
    wire N__24329;
    wire N__24326;
    wire N__24323;
    wire N__24320;
    wire N__24317;
    wire N__24314;
    wire N__24311;
    wire N__24308;
    wire N__24305;
    wire N__24302;
    wire N__24299;
    wire N__24296;
    wire N__24293;
    wire N__24290;
    wire N__24287;
    wire N__24284;
    wire N__24281;
    wire N__24280;
    wire N__24277;
    wire N__24276;
    wire N__24275;
    wire N__24274;
    wire N__24273;
    wire N__24270;
    wire N__24267;
    wire N__24258;
    wire N__24257;
    wire N__24256;
    wire N__24255;
    wire N__24254;
    wire N__24251;
    wire N__24246;
    wire N__24237;
    wire N__24230;
    wire N__24227;
    wire N__24226;
    wire N__24223;
    wire N__24220;
    wire N__24217;
    wire N__24214;
    wire N__24209;
    wire N__24206;
    wire N__24205;
    wire N__24202;
    wire N__24199;
    wire N__24196;
    wire N__24193;
    wire N__24188;
    wire N__24185;
    wire N__24182;
    wire N__24181;
    wire N__24180;
    wire N__24179;
    wire N__24176;
    wire N__24173;
    wire N__24170;
    wire N__24167;
    wire N__24162;
    wire N__24159;
    wire N__24156;
    wire N__24153;
    wire N__24150;
    wire N__24147;
    wire N__24144;
    wire N__24137;
    wire N__24134;
    wire N__24131;
    wire N__24128;
    wire N__24125;
    wire N__24122;
    wire N__24119;
    wire N__24116;
    wire N__24113;
    wire N__24110;
    wire N__24107;
    wire N__24104;
    wire N__24101;
    wire N__24098;
    wire N__24095;
    wire N__24092;
    wire N__24089;
    wire N__24088;
    wire N__24085;
    wire N__24082;
    wire N__24079;
    wire N__24076;
    wire N__24073;
    wire N__24070;
    wire N__24067;
    wire N__24064;
    wire N__24059;
    wire N__24056;
    wire N__24053;
    wire N__24050;
    wire N__24047;
    wire N__24044;
    wire N__24041;
    wire N__24038;
    wire N__24035;
    wire N__24032;
    wire N__24029;
    wire N__24026;
    wire N__24023;
    wire N__24020;
    wire N__24017;
    wire N__24014;
    wire N__24011;
    wire N__24008;
    wire N__24005;
    wire N__24002;
    wire N__23999;
    wire N__23996;
    wire N__23993;
    wire N__23990;
    wire N__23987;
    wire N__23984;
    wire N__23981;
    wire N__23978;
    wire N__23977;
    wire N__23976;
    wire N__23973;
    wire N__23970;
    wire N__23969;
    wire N__23968;
    wire N__23967;
    wire N__23966;
    wire N__23963;
    wire N__23960;
    wire N__23951;
    wire N__23950;
    wire N__23949;
    wire N__23948;
    wire N__23945;
    wire N__23942;
    wire N__23939;
    wire N__23936;
    wire N__23929;
    wire N__23926;
    wire N__23921;
    wire N__23916;
    wire N__23915;
    wire N__23914;
    wire N__23913;
    wire N__23912;
    wire N__23909;
    wire N__23904;
    wire N__23899;
    wire N__23894;
    wire N__23885;
    wire N__23882;
    wire N__23879;
    wire N__23876;
    wire N__23875;
    wire N__23874;
    wire N__23873;
    wire N__23872;
    wire N__23871;
    wire N__23870;
    wire N__23869;
    wire N__23868;
    wire N__23867;
    wire N__23866;
    wire N__23865;
    wire N__23862;
    wire N__23847;
    wire N__23838;
    wire N__23835;
    wire N__23828;
    wire N__23825;
    wire N__23822;
    wire N__23819;
    wire N__23818;
    wire N__23815;
    wire N__23812;
    wire N__23809;
    wire N__23804;
    wire N__23801;
    wire N__23800;
    wire N__23799;
    wire N__23796;
    wire N__23793;
    wire N__23790;
    wire N__23785;
    wire N__23782;
    wire N__23779;
    wire N__23774;
    wire N__23771;
    wire N__23768;
    wire N__23765;
    wire N__23764;
    wire N__23763;
    wire N__23756;
    wire N__23753;
    wire N__23750;
    wire N__23749;
    wire N__23748;
    wire N__23745;
    wire N__23742;
    wire N__23739;
    wire N__23736;
    wire N__23733;
    wire N__23726;
    wire N__23723;
    wire N__23720;
    wire N__23719;
    wire N__23718;
    wire N__23715;
    wire N__23710;
    wire N__23705;
    wire N__23704;
    wire N__23701;
    wire N__23698;
    wire N__23695;
    wire N__23692;
    wire N__23687;
    wire N__23684;
    wire N__23681;
    wire N__23678;
    wire N__23675;
    wire N__23674;
    wire N__23671;
    wire N__23668;
    wire N__23665;
    wire N__23662;
    wire N__23659;
    wire N__23654;
    wire N__23653;
    wire N__23650;
    wire N__23647;
    wire N__23644;
    wire N__23641;
    wire N__23638;
    wire N__23635;
    wire N__23632;
    wire N__23629;
    wire N__23626;
    wire N__23621;
    wire N__23618;
    wire N__23615;
    wire N__23612;
    wire N__23609;
    wire N__23606;
    wire N__23603;
    wire N__23600;
    wire N__23597;
    wire N__23594;
    wire N__23591;
    wire N__23588;
    wire N__23585;
    wire N__23582;
    wire N__23579;
    wire N__23576;
    wire N__23573;
    wire N__23570;
    wire N__23567;
    wire N__23564;
    wire N__23561;
    wire N__23558;
    wire N__23555;
    wire N__23552;
    wire N__23549;
    wire N__23546;
    wire N__23543;
    wire N__23540;
    wire N__23537;
    wire N__23534;
    wire N__23531;
    wire N__23528;
    wire N__23525;
    wire N__23522;
    wire N__23519;
    wire N__23516;
    wire N__23513;
    wire N__23512;
    wire N__23509;
    wire N__23506;
    wire N__23501;
    wire N__23498;
    wire N__23497;
    wire N__23496;
    wire N__23493;
    wire N__23488;
    wire N__23483;
    wire N__23480;
    wire N__23477;
    wire N__23474;
    wire N__23471;
    wire N__23468;
    wire N__23465;
    wire N__23462;
    wire N__23459;
    wire N__23458;
    wire N__23455;
    wire N__23452;
    wire N__23451;
    wire N__23450;
    wire N__23447;
    wire N__23440;
    wire N__23435;
    wire N__23432;
    wire N__23431;
    wire N__23430;
    wire N__23427;
    wire N__23424;
    wire N__23423;
    wire N__23420;
    wire N__23417;
    wire N__23410;
    wire N__23405;
    wire N__23404;
    wire N__23401;
    wire N__23398;
    wire N__23395;
    wire N__23392;
    wire N__23389;
    wire N__23386;
    wire N__23383;
    wire N__23380;
    wire N__23377;
    wire N__23372;
    wire N__23371;
    wire N__23368;
    wire N__23365;
    wire N__23362;
    wire N__23359;
    wire N__23356;
    wire N__23353;
    wire N__23350;
    wire N__23347;
    wire N__23344;
    wire N__23341;
    wire N__23336;
    wire N__23333;
    wire N__23332;
    wire N__23329;
    wire N__23326;
    wire N__23323;
    wire N__23320;
    wire N__23317;
    wire N__23314;
    wire N__23311;
    wire N__23308;
    wire N__23305;
    wire N__23300;
    wire N__23299;
    wire N__23298;
    wire N__23297;
    wire N__23296;
    wire N__23293;
    wire N__23288;
    wire N__23285;
    wire N__23282;
    wire N__23273;
    wire N__23272;
    wire N__23269;
    wire N__23268;
    wire N__23265;
    wire N__23262;
    wire N__23259;
    wire N__23256;
    wire N__23249;
    wire N__23248;
    wire N__23245;
    wire N__23242;
    wire N__23239;
    wire N__23234;
    wire N__23233;
    wire N__23230;
    wire N__23227;
    wire N__23224;
    wire N__23219;
    wire N__23216;
    wire N__23215;
    wire N__23212;
    wire N__23209;
    wire N__23206;
    wire N__23201;
    wire N__23200;
    wire N__23197;
    wire N__23194;
    wire N__23189;
    wire N__23186;
    wire N__23185;
    wire N__23182;
    wire N__23179;
    wire N__23176;
    wire N__23171;
    wire N__23170;
    wire N__23167;
    wire N__23164;
    wire N__23159;
    wire N__23156;
    wire N__23153;
    wire N__23152;
    wire N__23149;
    wire N__23146;
    wire N__23141;
    wire N__23138;
    wire N__23135;
    wire N__23132;
    wire N__23131;
    wire N__23128;
    wire N__23125;
    wire N__23120;
    wire N__23117;
    wire N__23116;
    wire N__23113;
    wire N__23110;
    wire N__23107;
    wire N__23104;
    wire N__23099;
    wire N__23096;
    wire N__23093;
    wire N__23092;
    wire N__23089;
    wire N__23086;
    wire N__23081;
    wire N__23078;
    wire N__23075;
    wire N__23074;
    wire N__23071;
    wire N__23068;
    wire N__23065;
    wire N__23060;
    wire N__23057;
    wire N__23056;
    wire N__23055;
    wire N__23052;
    wire N__23047;
    wire N__23042;
    wire N__23039;
    wire N__23036;
    wire N__23033;
    wire N__23030;
    wire N__23027;
    wire N__23024;
    wire N__23021;
    wire N__23018;
    wire N__23017;
    wire N__23016;
    wire N__23015;
    wire N__23014;
    wire N__23011;
    wire N__23006;
    wire N__23005;
    wire N__23004;
    wire N__23001;
    wire N__23000;
    wire N__22997;
    wire N__22996;
    wire N__22995;
    wire N__22994;
    wire N__22993;
    wire N__22992;
    wire N__22989;
    wire N__22986;
    wire N__22979;
    wire N__22972;
    wire N__22969;
    wire N__22968;
    wire N__22963;
    wire N__22960;
    wire N__22951;
    wire N__22946;
    wire N__22937;
    wire N__22936;
    wire N__22933;
    wire N__22930;
    wire N__22925;
    wire N__22924;
    wire N__22923;
    wire N__22920;
    wire N__22917;
    wire N__22916;
    wire N__22915;
    wire N__22912;
    wire N__22909;
    wire N__22908;
    wire N__22907;
    wire N__22904;
    wire N__22897;
    wire N__22894;
    wire N__22893;
    wire N__22890;
    wire N__22887;
    wire N__22884;
    wire N__22881;
    wire N__22878;
    wire N__22875;
    wire N__22872;
    wire N__22869;
    wire N__22864;
    wire N__22863;
    wire N__22862;
    wire N__22859;
    wire N__22856;
    wire N__22853;
    wire N__22848;
    wire N__22843;
    wire N__22832;
    wire N__22831;
    wire N__22830;
    wire N__22829;
    wire N__22828;
    wire N__22827;
    wire N__22826;
    wire N__22823;
    wire N__22820;
    wire N__22817;
    wire N__22816;
    wire N__22813;
    wire N__22812;
    wire N__22809;
    wire N__22804;
    wire N__22801;
    wire N__22796;
    wire N__22793;
    wire N__22790;
    wire N__22787;
    wire N__22786;
    wire N__22785;
    wire N__22782;
    wire N__22777;
    wire N__22770;
    wire N__22767;
    wire N__22762;
    wire N__22759;
    wire N__22756;
    wire N__22753;
    wire N__22748;
    wire N__22739;
    wire N__22738;
    wire N__22737;
    wire N__22734;
    wire N__22733;
    wire N__22728;
    wire N__22725;
    wire N__22724;
    wire N__22721;
    wire N__22720;
    wire N__22717;
    wire N__22714;
    wire N__22713;
    wire N__22710;
    wire N__22707;
    wire N__22704;
    wire N__22701;
    wire N__22698;
    wire N__22695;
    wire N__22690;
    wire N__22685;
    wire N__22676;
    wire N__22673;
    wire N__22670;
    wire N__22667;
    wire N__22664;
    wire N__22661;
    wire N__22658;
    wire N__22655;
    wire N__22652;
    wire N__22649;
    wire N__22646;
    wire N__22643;
    wire N__22642;
    wire N__22639;
    wire N__22638;
    wire N__22635;
    wire N__22634;
    wire N__22631;
    wire N__22628;
    wire N__22627;
    wire N__22626;
    wire N__22625;
    wire N__22624;
    wire N__22621;
    wire N__22620;
    wire N__22619;
    wire N__22616;
    wire N__22611;
    wire N__22608;
    wire N__22601;
    wire N__22598;
    wire N__22593;
    wire N__22590;
    wire N__22583;
    wire N__22580;
    wire N__22577;
    wire N__22574;
    wire N__22573;
    wire N__22570;
    wire N__22567;
    wire N__22564;
    wire N__22561;
    wire N__22558;
    wire N__22555;
    wire N__22544;
    wire N__22541;
    wire N__22538;
    wire N__22535;
    wire N__22532;
    wire N__22531;
    wire N__22528;
    wire N__22527;
    wire N__22526;
    wire N__22525;
    wire N__22524;
    wire N__22523;
    wire N__22520;
    wire N__22515;
    wire N__22512;
    wire N__22511;
    wire N__22508;
    wire N__22505;
    wire N__22502;
    wire N__22501;
    wire N__22500;
    wire N__22499;
    wire N__22494;
    wire N__22491;
    wire N__22488;
    wire N__22481;
    wire N__22476;
    wire N__22473;
    wire N__22460;
    wire N__22457;
    wire N__22454;
    wire N__22451;
    wire N__22448;
    wire N__22445;
    wire N__22444;
    wire N__22443;
    wire N__22440;
    wire N__22439;
    wire N__22438;
    wire N__22435;
    wire N__22432;
    wire N__22431;
    wire N__22430;
    wire N__22429;
    wire N__22426;
    wire N__22421;
    wire N__22420;
    wire N__22415;
    wire N__22410;
    wire N__22407;
    wire N__22406;
    wire N__22405;
    wire N__22404;
    wire N__22399;
    wire N__22396;
    wire N__22389;
    wire N__22386;
    wire N__22381;
    wire N__22370;
    wire N__22367;
    wire N__22364;
    wire N__22361;
    wire N__22358;
    wire N__22355;
    wire N__22352;
    wire N__22349;
    wire N__22346;
    wire N__22343;
    wire N__22340;
    wire N__22337;
    wire N__22334;
    wire N__22331;
    wire N__22328;
    wire N__22325;
    wire N__22322;
    wire N__22319;
    wire N__22316;
    wire N__22313;
    wire N__22310;
    wire N__22307;
    wire N__22304;
    wire N__22301;
    wire N__22298;
    wire N__22295;
    wire N__22292;
    wire N__22289;
    wire N__22286;
    wire N__22283;
    wire N__22280;
    wire N__22277;
    wire N__22274;
    wire N__22271;
    wire N__22270;
    wire N__22267;
    wire N__22266;
    wire N__22259;
    wire N__22256;
    wire N__22253;
    wire N__22250;
    wire N__22249;
    wire N__22248;
    wire N__22245;
    wire N__22238;
    wire N__22237;
    wire N__22234;
    wire N__22231;
    wire N__22228;
    wire N__22225;
    wire N__22222;
    wire N__22217;
    wire N__22214;
    wire N__22211;
    wire N__22208;
    wire N__22205;
    wire N__22202;
    wire N__22199;
    wire N__22196;
    wire N__22195;
    wire N__22192;
    wire N__22189;
    wire N__22188;
    wire N__22187;
    wire N__22186;
    wire N__22183;
    wire N__22180;
    wire N__22177;
    wire N__22174;
    wire N__22171;
    wire N__22170;
    wire N__22169;
    wire N__22166;
    wire N__22163;
    wire N__22160;
    wire N__22157;
    wire N__22154;
    wire N__22151;
    wire N__22150;
    wire N__22149;
    wire N__22146;
    wire N__22139;
    wire N__22136;
    wire N__22131;
    wire N__22128;
    wire N__22125;
    wire N__22122;
    wire N__22109;
    wire N__22108;
    wire N__22107;
    wire N__22106;
    wire N__22097;
    wire N__22096;
    wire N__22095;
    wire N__22092;
    wire N__22089;
    wire N__22088;
    wire N__22087;
    wire N__22086;
    wire N__22085;
    wire N__22082;
    wire N__22077;
    wire N__22070;
    wire N__22067;
    wire N__22058;
    wire N__22057;
    wire N__22056;
    wire N__22053;
    wire N__22050;
    wire N__22047;
    wire N__22046;
    wire N__22043;
    wire N__22040;
    wire N__22037;
    wire N__22034;
    wire N__22033;
    wire N__22030;
    wire N__22027;
    wire N__22022;
    wire N__22019;
    wire N__22016;
    wire N__22011;
    wire N__22008;
    wire N__22001;
    wire N__21998;
    wire N__21995;
    wire N__21992;
    wire N__21989;
    wire N__21986;
    wire N__21983;
    wire N__21980;
    wire N__21977;
    wire N__21974;
    wire N__21971;
    wire N__21968;
    wire N__21965;
    wire N__21962;
    wire N__21959;
    wire N__21956;
    wire N__21953;
    wire N__21950;
    wire N__21947;
    wire N__21944;
    wire N__21941;
    wire N__21938;
    wire N__21935;
    wire N__21932;
    wire N__21931;
    wire N__21928;
    wire N__21925;
    wire N__21920;
    wire N__21917;
    wire N__21914;
    wire N__21911;
    wire N__21908;
    wire N__21905;
    wire N__21902;
    wire N__21899;
    wire N__21896;
    wire N__21893;
    wire N__21892;
    wire N__21891;
    wire N__21890;
    wire N__21889;
    wire N__21888;
    wire N__21883;
    wire N__21882;
    wire N__21879;
    wire N__21878;
    wire N__21871;
    wire N__21868;
    wire N__21865;
    wire N__21864;
    wire N__21863;
    wire N__21860;
    wire N__21857;
    wire N__21854;
    wire N__21851;
    wire N__21848;
    wire N__21845;
    wire N__21842;
    wire N__21827;
    wire N__21824;
    wire N__21821;
    wire N__21818;
    wire N__21815;
    wire N__21812;
    wire N__21809;
    wire N__21806;
    wire N__21803;
    wire N__21800;
    wire N__21797;
    wire N__21794;
    wire N__21791;
    wire N__21788;
    wire N__21785;
    wire N__21782;
    wire N__21779;
    wire N__21776;
    wire N__21773;
    wire N__21770;
    wire N__21767;
    wire N__21764;
    wire N__21761;
    wire N__21758;
    wire N__21755;
    wire N__21752;
    wire N__21749;
    wire N__21746;
    wire N__21743;
    wire N__21740;
    wire N__21737;
    wire N__21734;
    wire N__21731;
    wire N__21728;
    wire N__21725;
    wire N__21722;
    wire N__21719;
    wire N__21718;
    wire N__21717;
    wire N__21714;
    wire N__21711;
    wire N__21710;
    wire N__21709;
    wire N__21708;
    wire N__21707;
    wire N__21706;
    wire N__21705;
    wire N__21704;
    wire N__21701;
    wire N__21698;
    wire N__21695;
    wire N__21692;
    wire N__21687;
    wire N__21678;
    wire N__21665;
    wire N__21664;
    wire N__21663;
    wire N__21662;
    wire N__21655;
    wire N__21654;
    wire N__21651;
    wire N__21648;
    wire N__21645;
    wire N__21642;
    wire N__21637;
    wire N__21636;
    wire N__21635;
    wire N__21634;
    wire N__21633;
    wire N__21632;
    wire N__21631;
    wire N__21628;
    wire N__21625;
    wire N__21622;
    wire N__21619;
    wire N__21610;
    wire N__21599;
    wire N__21596;
    wire N__21595;
    wire N__21592;
    wire N__21589;
    wire N__21586;
    wire N__21583;
    wire N__21580;
    wire N__21577;
    wire N__21574;
    wire N__21571;
    wire N__21568;
    wire N__21565;
    wire N__21562;
    wire N__21559;
    wire N__21556;
    wire N__21553;
    wire N__21550;
    wire N__21547;
    wire N__21544;
    wire N__21541;
    wire N__21538;
    wire N__21535;
    wire N__21532;
    wire N__21529;
    wire N__21526;
    wire N__21523;
    wire N__21520;
    wire N__21517;
    wire N__21514;
    wire N__21511;
    wire N__21506;
    wire N__21503;
    wire N__21500;
    wire N__21497;
    wire N__21494;
    wire N__21491;
    wire N__21488;
    wire N__21485;
    wire N__21482;
    wire N__21479;
    wire N__21476;
    wire N__21473;
    wire N__21470;
    wire N__21469;
    wire N__21468;
    wire N__21467;
    wire N__21464;
    wire N__21461;
    wire N__21458;
    wire N__21457;
    wire N__21456;
    wire N__21455;
    wire N__21454;
    wire N__21453;
    wire N__21450;
    wire N__21449;
    wire N__21448;
    wire N__21447;
    wire N__21440;
    wire N__21437;
    wire N__21434;
    wire N__21431;
    wire N__21428;
    wire N__21427;
    wire N__21426;
    wire N__21423;
    wire N__21420;
    wire N__21417;
    wire N__21414;
    wire N__21411;
    wire N__21410;
    wire N__21403;
    wire N__21398;
    wire N__21395;
    wire N__21392;
    wire N__21391;
    wire N__21388;
    wire N__21381;
    wire N__21378;
    wire N__21375;
    wire N__21368;
    wire N__21365;
    wire N__21362;
    wire N__21359;
    wire N__21352;
    wire N__21349;
    wire N__21344;
    wire N__21341;
    wire N__21338;
    wire N__21335;
    wire N__21332;
    wire N__21327;
    wire N__21324;
    wire N__21319;
    wire N__21314;
    wire N__21313;
    wire N__21312;
    wire N__21309;
    wire N__21304;
    wire N__21303;
    wire N__21302;
    wire N__21299;
    wire N__21296;
    wire N__21293;
    wire N__21290;
    wire N__21287;
    wire N__21284;
    wire N__21281;
    wire N__21278;
    wire N__21269;
    wire N__21266;
    wire N__21265;
    wire N__21262;
    wire N__21259;
    wire N__21258;
    wire N__21255;
    wire N__21254;
    wire N__21253;
    wire N__21252;
    wire N__21251;
    wire N__21250;
    wire N__21249;
    wire N__21244;
    wire N__21241;
    wire N__21236;
    wire N__21229;
    wire N__21226;
    wire N__21223;
    wire N__21218;
    wire N__21209;
    wire N__21206;
    wire N__21203;
    wire N__21200;
    wire N__21197;
    wire N__21194;
    wire N__21191;
    wire N__21190;
    wire N__21185;
    wire N__21182;
    wire N__21181;
    wire N__21178;
    wire N__21175;
    wire N__21170;
    wire N__21167;
    wire N__21166;
    wire N__21165;
    wire N__21160;
    wire N__21157;
    wire N__21154;
    wire N__21151;
    wire N__21150;
    wire N__21147;
    wire N__21146;
    wire N__21145;
    wire N__21142;
    wire N__21139;
    wire N__21136;
    wire N__21131;
    wire N__21122;
    wire N__21119;
    wire N__21116;
    wire N__21113;
    wire N__21112;
    wire N__21111;
    wire N__21110;
    wire N__21109;
    wire N__21108;
    wire N__21105;
    wire N__21102;
    wire N__21097;
    wire N__21092;
    wire N__21083;
    wire N__21082;
    wire N__21079;
    wire N__21078;
    wire N__21077;
    wire N__21076;
    wire N__21073;
    wire N__21068;
    wire N__21067;
    wire N__21064;
    wire N__21061;
    wire N__21058;
    wire N__21055;
    wire N__21052;
    wire N__21049;
    wire N__21046;
    wire N__21043;
    wire N__21040;
    wire N__21035;
    wire N__21026;
    wire N__21023;
    wire N__21022;
    wire N__21019;
    wire N__21018;
    wire N__21011;
    wire N__21008;
    wire N__21005;
    wire N__21002;
    wire N__20999;
    wire N__20996;
    wire N__20993;
    wire N__20990;
    wire N__20987;
    wire N__20986;
    wire N__20983;
    wire N__20980;
    wire N__20975;
    wire N__20972;
    wire N__20969;
    wire N__20968;
    wire N__20965;
    wire N__20964;
    wire N__20961;
    wire N__20958;
    wire N__20955;
    wire N__20948;
    wire N__20947;
    wire N__20946;
    wire N__20943;
    wire N__20942;
    wire N__20939;
    wire N__20936;
    wire N__20933;
    wire N__20930;
    wire N__20927;
    wire N__20918;
    wire N__20915;
    wire N__20912;
    wire N__20909;
    wire N__20906;
    wire N__20903;
    wire N__20902;
    wire N__20899;
    wire N__20896;
    wire N__20891;
    wire N__20888;
    wire N__20885;
    wire N__20882;
    wire N__20879;
    wire N__20876;
    wire N__20873;
    wire N__20870;
    wire N__20867;
    wire N__20864;
    wire N__20861;
    wire N__20858;
    wire N__20855;
    wire N__20852;
    wire N__20849;
    wire N__20846;
    wire N__20843;
    wire N__20840;
    wire N__20837;
    wire N__20834;
    wire N__20831;
    wire N__20828;
    wire N__20825;
    wire N__20822;
    wire N__20819;
    wire N__20816;
    wire N__20813;
    wire N__20810;
    wire N__20807;
    wire N__20804;
    wire N__20801;
    wire N__20798;
    wire N__20795;
    wire N__20792;
    wire N__20789;
    wire N__20786;
    wire N__20783;
    wire N__20780;
    wire N__20779;
    wire N__20776;
    wire N__20773;
    wire N__20770;
    wire N__20767;
    wire N__20764;
    wire N__20761;
    wire N__20756;
    wire N__20753;
    wire N__20750;
    wire N__20747;
    wire N__20744;
    wire N__20741;
    wire N__20738;
    wire N__20735;
    wire N__20734;
    wire N__20731;
    wire N__20728;
    wire N__20723;
    wire N__20720;
    wire N__20717;
    wire N__20714;
    wire N__20711;
    wire N__20708;
    wire N__20705;
    wire N__20702;
    wire N__20701;
    wire N__20698;
    wire N__20695;
    wire N__20690;
    wire N__20689;
    wire N__20686;
    wire N__20685;
    wire N__20684;
    wire N__20683;
    wire N__20682;
    wire N__20681;
    wire N__20680;
    wire N__20679;
    wire N__20672;
    wire N__20659;
    wire N__20656;
    wire N__20653;
    wire N__20648;
    wire N__20647;
    wire N__20646;
    wire N__20645;
    wire N__20644;
    wire N__20643;
    wire N__20642;
    wire N__20641;
    wire N__20640;
    wire N__20639;
    wire N__20638;
    wire N__20627;
    wire N__20614;
    wire N__20611;
    wire N__20606;
    wire N__20603;
    wire N__20602;
    wire N__20599;
    wire N__20596;
    wire N__20591;
    wire N__20588;
    wire N__20585;
    wire N__20582;
    wire N__20579;
    wire N__20576;
    wire N__20573;
    wire N__20570;
    wire N__20567;
    wire N__20564;
    wire N__20561;
    wire N__20558;
    wire N__20555;
    wire N__20552;
    wire N__20549;
    wire N__20546;
    wire N__20543;
    wire N__20540;
    wire N__20537;
    wire N__20534;
    wire N__20533;
    wire N__20530;
    wire N__20527;
    wire N__20524;
    wire N__20521;
    wire N__20518;
    wire N__20515;
    wire N__20512;
    wire N__20509;
    wire N__20506;
    wire N__20503;
    wire N__20500;
    wire N__20497;
    wire N__20494;
    wire N__20491;
    wire N__20488;
    wire N__20485;
    wire N__20482;
    wire N__20479;
    wire N__20476;
    wire N__20473;
    wire N__20470;
    wire N__20467;
    wire N__20464;
    wire N__20461;
    wire N__20458;
    wire N__20455;
    wire N__20452;
    wire N__20449;
    wire N__20444;
    wire N__20441;
    wire N__20438;
    wire N__20435;
    wire N__20432;
    wire N__20429;
    wire N__20426;
    wire N__20425;
    wire N__20422;
    wire N__20419;
    wire N__20416;
    wire N__20413;
    wire N__20410;
    wire N__20407;
    wire N__20404;
    wire N__20401;
    wire N__20396;
    wire N__20393;
    wire N__20390;
    wire N__20387;
    wire N__20384;
    wire N__20381;
    wire N__20378;
    wire N__20375;
    wire N__20372;
    wire N__20369;
    wire N__20366;
    wire N__20363;
    wire N__20360;
    wire N__20357;
    wire N__20354;
    wire N__20351;
    wire N__20350;
    wire N__20349;
    wire N__20346;
    wire N__20341;
    wire N__20338;
    wire N__20337;
    wire N__20334;
    wire N__20331;
    wire N__20328;
    wire N__20321;
    wire N__20320;
    wire N__20317;
    wire N__20314;
    wire N__20311;
    wire N__20310;
    wire N__20307;
    wire N__20304;
    wire N__20301;
    wire N__20298;
    wire N__20293;
    wire N__20288;
    wire N__20285;
    wire N__20282;
    wire N__20279;
    wire N__20276;
    wire N__20273;
    wire N__20270;
    wire N__20269;
    wire N__20266;
    wire N__20261;
    wire N__20260;
    wire N__20257;
    wire N__20254;
    wire N__20249;
    wire N__20248;
    wire N__20245;
    wire N__20242;
    wire N__20241;
    wire N__20236;
    wire N__20233;
    wire N__20228;
    wire N__20225;
    wire N__20222;
    wire N__20219;
    wire N__20216;
    wire N__20213;
    wire N__20212;
    wire N__20211;
    wire N__20210;
    wire N__20205;
    wire N__20200;
    wire N__20195;
    wire N__20192;
    wire N__20189;
    wire N__20186;
    wire N__20183;
    wire N__20180;
    wire N__20177;
    wire N__20174;
    wire N__20171;
    wire N__20168;
    wire N__20165;
    wire N__20162;
    wire N__20159;
    wire N__20156;
    wire N__20153;
    wire N__20150;
    wire N__20149;
    wire N__20146;
    wire N__20143;
    wire N__20140;
    wire N__20137;
    wire N__20134;
    wire N__20131;
    wire N__20128;
    wire N__20125;
    wire N__20122;
    wire N__20119;
    wire N__20116;
    wire N__20113;
    wire N__20110;
    wire N__20107;
    wire N__20104;
    wire N__20101;
    wire N__20098;
    wire N__20095;
    wire N__20092;
    wire N__20089;
    wire N__20086;
    wire N__20083;
    wire N__20080;
    wire N__20077;
    wire N__20074;
    wire N__20071;
    wire N__20068;
    wire N__20065;
    wire N__20062;
    wire N__20059;
    wire N__20056;
    wire N__20053;
    wire N__20048;
    wire N__20045;
    wire N__20042;
    wire N__20039;
    wire N__20036;
    wire N__20033;
    wire N__20030;
    wire N__20027;
    wire N__20024;
    wire N__20021;
    wire N__20018;
    wire N__20017;
    wire N__20014;
    wire N__20011;
    wire N__20008;
    wire N__20005;
    wire N__20002;
    wire N__19999;
    wire N__19996;
    wire N__19993;
    wire N__19990;
    wire N__19987;
    wire N__19984;
    wire N__19981;
    wire N__19978;
    wire N__19975;
    wire N__19972;
    wire N__19969;
    wire N__19966;
    wire N__19963;
    wire N__19960;
    wire N__19957;
    wire N__19954;
    wire N__19951;
    wire N__19948;
    wire N__19945;
    wire N__19942;
    wire N__19939;
    wire N__19936;
    wire N__19933;
    wire N__19928;
    wire N__19925;
    wire N__19922;
    wire N__19919;
    wire N__19916;
    wire N__19913;
    wire N__19910;
    wire N__19907;
    wire N__19904;
    wire N__19901;
    wire N__19900;
    wire N__19897;
    wire N__19894;
    wire N__19891;
    wire N__19888;
    wire N__19885;
    wire N__19882;
    wire N__19879;
    wire N__19876;
    wire N__19873;
    wire N__19870;
    wire N__19867;
    wire N__19864;
    wire N__19861;
    wire N__19858;
    wire N__19855;
    wire N__19852;
    wire N__19849;
    wire N__19846;
    wire N__19843;
    wire N__19840;
    wire N__19837;
    wire N__19834;
    wire N__19831;
    wire N__19828;
    wire N__19825;
    wire N__19822;
    wire N__19819;
    wire N__19816;
    wire N__19811;
    wire N__19808;
    wire N__19805;
    wire N__19802;
    wire N__19799;
    wire N__19796;
    wire N__19793;
    wire N__19790;
    wire N__19787;
    wire N__19784;
    wire N__19781;
    wire N__19778;
    wire N__19775;
    wire N__19772;
    wire N__19769;
    wire N__19766;
    wire N__19763;
    wire N__19760;
    wire N__19757;
    wire N__19754;
    wire N__19751;
    wire N__19748;
    wire N__19745;
    wire N__19742;
    wire N__19739;
    wire N__19736;
    wire N__19733;
    wire N__19730;
    wire N__19729;
    wire N__19728;
    wire N__19725;
    wire N__19720;
    wire N__19715;
    wire N__19712;
    wire N__19709;
    wire N__19706;
    wire N__19703;
    wire N__19700;
    wire N__19697;
    wire N__19694;
    wire N__19693;
    wire N__19692;
    wire N__19691;
    wire N__19688;
    wire N__19685;
    wire N__19682;
    wire N__19679;
    wire N__19676;
    wire N__19671;
    wire N__19664;
    wire N__19661;
    wire N__19658;
    wire N__19655;
    wire N__19652;
    wire N__19651;
    wire N__19648;
    wire N__19645;
    wire N__19642;
    wire N__19639;
    wire N__19636;
    wire N__19633;
    wire N__19630;
    wire N__19627;
    wire N__19624;
    wire N__19621;
    wire N__19618;
    wire N__19615;
    wire N__19612;
    wire N__19609;
    wire N__19606;
    wire N__19603;
    wire N__19600;
    wire N__19597;
    wire N__19594;
    wire N__19591;
    wire N__19588;
    wire N__19585;
    wire N__19582;
    wire N__19579;
    wire N__19576;
    wire N__19573;
    wire N__19570;
    wire N__19565;
    wire N__19562;
    wire N__19559;
    wire N__19556;
    wire N__19553;
    wire N__19550;
    wire N__19547;
    wire N__19544;
    wire N__19541;
    wire N__19538;
    wire N__19535;
    wire N__19532;
    wire N__19529;
    wire N__19526;
    wire N__19525;
    wire N__19522;
    wire N__19519;
    wire N__19516;
    wire N__19511;
    wire N__19508;
    wire N__19505;
    wire N__19502;
    wire N__19499;
    wire N__19496;
    wire N__19493;
    wire N__19490;
    wire N__19487;
    wire N__19484;
    wire N__19481;
    wire N__19478;
    wire N__19475;
    wire N__19472;
    wire N__19471;
    wire N__19468;
    wire N__19465;
    wire N__19462;
    wire N__19459;
    wire N__19456;
    wire N__19453;
    wire N__19450;
    wire N__19447;
    wire N__19444;
    wire N__19441;
    wire N__19438;
    wire N__19435;
    wire N__19432;
    wire N__19429;
    wire N__19426;
    wire N__19423;
    wire N__19420;
    wire N__19417;
    wire N__19414;
    wire N__19411;
    wire N__19408;
    wire N__19405;
    wire N__19402;
    wire N__19399;
    wire N__19394;
    wire N__19391;
    wire N__19388;
    wire N__19385;
    wire N__19382;
    wire N__19379;
    wire N__19376;
    wire N__19373;
    wire N__19370;
    wire N__19367;
    wire N__19364;
    wire N__19361;
    wire N__19358;
    wire N__19355;
    wire N__19352;
    wire N__19349;
    wire N__19346;
    wire N__19343;
    wire N__19340;
    wire N__19337;
    wire N__19334;
    wire N__19331;
    wire N__19328;
    wire N__19325;
    wire N__19322;
    wire N__19319;
    wire N__19316;
    wire N__19313;
    wire N__19310;
    wire N__19307;
    wire N__19304;
    wire N__19301;
    wire N__19298;
    wire N__19295;
    wire N__19292;
    wire N__19289;
    wire N__19286;
    wire N__19283;
    wire N__19282;
    wire N__19279;
    wire N__19276;
    wire N__19275;
    wire N__19270;
    wire N__19267;
    wire N__19264;
    wire N__19261;
    wire N__19256;
    wire N__19253;
    wire N__19250;
    wire N__19249;
    wire N__19248;
    wire N__19247;
    wire N__19246;
    wire N__19245;
    wire N__19244;
    wire N__19243;
    wire N__19242;
    wire N__19241;
    wire N__19236;
    wire N__19229;
    wire N__19218;
    wire N__19211;
    wire N__19210;
    wire N__19207;
    wire N__19204;
    wire N__19201;
    wire N__19200;
    wire N__19195;
    wire N__19192;
    wire N__19189;
    wire N__19186;
    wire N__19181;
    wire N__19180;
    wire N__19179;
    wire N__19178;
    wire N__19175;
    wire N__19172;
    wire N__19169;
    wire N__19168;
    wire N__19167;
    wire N__19166;
    wire N__19165;
    wire N__19164;
    wire N__19159;
    wire N__19156;
    wire N__19151;
    wire N__19142;
    wire N__19139;
    wire N__19130;
    wire N__19127;
    wire N__19124;
    wire N__19123;
    wire N__19120;
    wire N__19117;
    wire N__19112;
    wire N__19111;
    wire N__19108;
    wire N__19105;
    wire N__19104;
    wire N__19101;
    wire N__19098;
    wire N__19095;
    wire N__19092;
    wire N__19089;
    wire N__19086;
    wire N__19079;
    wire N__19076;
    wire N__19073;
    wire N__19070;
    wire N__19067;
    wire N__19064;
    wire N__19061;
    wire N__19060;
    wire N__19059;
    wire N__19056;
    wire N__19053;
    wire N__19050;
    wire N__19043;
    wire N__19040;
    wire N__19037;
    wire N__19036;
    wire N__19035;
    wire N__19032;
    wire N__19029;
    wire N__19026;
    wire N__19019;
    wire N__19016;
    wire N__19013;
    wire N__19010;
    wire N__19007;
    wire N__19004;
    wire N__19001;
    wire N__18998;
    wire N__18997;
    wire N__18994;
    wire N__18991;
    wire N__18986;
    wire N__18983;
    wire N__18980;
    wire N__18979;
    wire N__18976;
    wire N__18973;
    wire N__18968;
    wire N__18967;
    wire N__18966;
    wire N__18961;
    wire N__18958;
    wire N__18953;
    wire N__18950;
    wire N__18949;
    wire N__18948;
    wire N__18943;
    wire N__18940;
    wire N__18935;
    wire N__18932;
    wire N__18929;
    wire N__18926;
    wire N__18923;
    wire N__18920;
    wire N__18917;
    wire N__18914;
    wire N__18911;
    wire N__18908;
    wire N__18905;
    wire N__18902;
    wire N__18899;
    wire N__18896;
    wire N__18893;
    wire N__18890;
    wire N__18887;
    wire N__18884;
    wire N__18881;
    wire N__18878;
    wire N__18875;
    wire N__18874;
    wire N__18871;
    wire N__18868;
    wire N__18865;
    wire N__18862;
    wire N__18859;
    wire N__18856;
    wire N__18853;
    wire N__18850;
    wire N__18845;
    wire N__18842;
    wire N__18841;
    wire N__18838;
    wire N__18835;
    wire N__18834;
    wire N__18831;
    wire N__18828;
    wire N__18825;
    wire N__18820;
    wire N__18817;
    wire N__18812;
    wire N__18809;
    wire N__18808;
    wire N__18805;
    wire N__18802;
    wire N__18797;
    wire N__18796;
    wire N__18793;
    wire N__18790;
    wire N__18785;
    wire N__18784;
    wire N__18781;
    wire N__18780;
    wire N__18777;
    wire N__18774;
    wire N__18771;
    wire N__18768;
    wire N__18765;
    wire N__18762;
    wire N__18759;
    wire N__18754;
    wire N__18749;
    wire N__18746;
    wire N__18743;
    wire N__18740;
    wire N__18737;
    wire N__18734;
    wire N__18731;
    wire N__18728;
    wire N__18725;
    wire N__18724;
    wire N__18721;
    wire N__18718;
    wire N__18715;
    wire N__18712;
    wire N__18709;
    wire N__18706;
    wire N__18703;
    wire N__18700;
    wire N__18697;
    wire N__18694;
    wire N__18691;
    wire N__18688;
    wire N__18685;
    wire N__18682;
    wire N__18679;
    wire N__18676;
    wire N__18673;
    wire N__18670;
    wire N__18667;
    wire N__18664;
    wire N__18661;
    wire N__18658;
    wire N__18655;
    wire N__18652;
    wire N__18649;
    wire N__18646;
    wire N__18643;
    wire N__18640;
    wire N__18635;
    wire N__18632;
    wire N__18629;
    wire N__18626;
    wire N__18623;
    wire N__18620;
    wire N__18617;
    wire N__18614;
    wire N__18611;
    wire N__18608;
    wire N__18605;
    wire N__18602;
    wire N__18599;
    wire N__18596;
    wire N__18593;
    wire N__18590;
    wire N__18587;
    wire N__18584;
    wire N__18581;
    wire N__18578;
    wire N__18575;
    wire N__18572;
    wire N__18569;
    wire N__18566;
    wire N__18563;
    wire N__18560;
    wire N__18557;
    wire N__18554;
    wire N__18551;
    wire N__18548;
    wire N__18545;
    wire N__18542;
    wire N__18539;
    wire N__18536;
    wire N__18533;
    wire N__18530;
    wire N__18527;
    wire N__18524;
    wire N__18521;
    wire N__18518;
    wire N__18515;
    wire N__18512;
    wire N__18509;
    wire N__18506;
    wire N__18503;
    wire N__18500;
    wire N__18497;
    wire N__18494;
    wire N__18491;
    wire N__18488;
    wire N__18485;
    wire N__18482;
    wire N__18479;
    wire N__18476;
    wire N__18473;
    wire N__18470;
    wire N__18469;
    wire N__18466;
    wire N__18463;
    wire N__18460;
    wire N__18457;
    wire N__18454;
    wire N__18451;
    wire N__18448;
    wire N__18445;
    wire N__18442;
    wire N__18439;
    wire N__18436;
    wire N__18433;
    wire N__18430;
    wire N__18427;
    wire N__18424;
    wire N__18421;
    wire N__18418;
    wire N__18415;
    wire N__18412;
    wire N__18409;
    wire N__18406;
    wire N__18403;
    wire N__18400;
    wire N__18397;
    wire N__18394;
    wire N__18391;
    wire N__18388;
    wire N__18385;
    wire N__18382;
    wire N__18377;
    wire N__18374;
    wire N__18371;
    wire N__18368;
    wire N__18365;
    wire N__18362;
    wire N__18361;
    wire N__18358;
    wire N__18355;
    wire N__18352;
    wire N__18351;
    wire N__18348;
    wire N__18345;
    wire N__18342;
    wire N__18335;
    wire N__18332;
    wire N__18329;
    wire N__18326;
    wire N__18325;
    wire N__18324;
    wire N__18323;
    wire N__18322;
    wire N__18319;
    wire N__18318;
    wire N__18315;
    wire N__18314;
    wire N__18313;
    wire N__18310;
    wire N__18307;
    wire N__18306;
    wire N__18303;
    wire N__18300;
    wire N__18295;
    wire N__18288;
    wire N__18285;
    wire N__18280;
    wire N__18269;
    wire N__18266;
    wire N__18263;
    wire N__18262;
    wire N__18261;
    wire N__18260;
    wire N__18259;
    wire N__18258;
    wire N__18257;
    wire N__18256;
    wire N__18255;
    wire N__18254;
    wire N__18253;
    wire N__18250;
    wire N__18247;
    wire N__18242;
    wire N__18227;
    wire N__18218;
    wire N__18215;
    wire N__18212;
    wire N__18209;
    wire N__18208;
    wire N__18205;
    wire N__18204;
    wire N__18203;
    wire N__18200;
    wire N__18197;
    wire N__18194;
    wire N__18191;
    wire N__18188;
    wire N__18183;
    wire N__18180;
    wire N__18177;
    wire N__18174;
    wire N__18167;
    wire N__18166;
    wire N__18161;
    wire N__18158;
    wire N__18155;
    wire N__18152;
    wire N__18149;
    wire N__18146;
    wire N__18143;
    wire N__18140;
    wire N__18139;
    wire N__18134;
    wire N__18131;
    wire N__18128;
    wire N__18125;
    wire N__18122;
    wire N__18119;
    wire N__18116;
    wire N__18113;
    wire N__18112;
    wire N__18109;
    wire N__18106;
    wire N__18103;
    wire N__18100;
    wire N__18097;
    wire N__18094;
    wire N__18089;
    wire N__18086;
    wire N__18083;
    wire N__18080;
    wire N__18077;
    wire N__18074;
    wire N__18071;
    wire N__18068;
    wire N__18065;
    wire N__18062;
    wire N__18059;
    wire N__18056;
    wire N__18053;
    wire N__18050;
    wire N__18047;
    wire N__18044;
    wire N__18041;
    wire N__18038;
    wire N__18035;
    wire N__18032;
    wire N__18029;
    wire N__18026;
    wire N__18023;
    wire N__18020;
    wire N__18017;
    wire N__18014;
    wire N__18013;
    wire N__18010;
    wire N__18007;
    wire N__18002;
    wire N__17999;
    wire N__17998;
    wire N__17995;
    wire N__17992;
    wire N__17987;
    wire N__17986;
    wire N__17983;
    wire N__17980;
    wire N__17977;
    wire N__17974;
    wire N__17971;
    wire N__17966;
    wire N__17963;
    wire N__17960;
    wire N__17957;
    wire N__17954;
    wire N__17951;
    wire N__17948;
    wire N__17945;
    wire N__17942;
    wire N__17939;
    wire N__17936;
    wire N__17933;
    wire N__17930;
    wire N__17927;
    wire N__17924;
    wire N__17921;
    wire N__17920;
    wire N__17917;
    wire N__17914;
    wire N__17911;
    wire N__17906;
    wire N__17903;
    wire N__17900;
    wire N__17897;
    wire N__17894;
    wire N__17891;
    wire N__17888;
    wire N__17885;
    wire N__17882;
    wire N__17879;
    wire N__17876;
    wire N__17873;
    wire N__17870;
    wire N__17867;
    wire N__17864;
    wire N__17861;
    wire N__17858;
    wire N__17857;
    wire N__17854;
    wire N__17851;
    wire N__17848;
    wire N__17843;
    wire N__17840;
    wire N__17837;
    wire N__17834;
    wire N__17831;
    wire N__17828;
    wire N__17825;
    wire N__17822;
    wire N__17821;
    wire N__17818;
    wire N__17815;
    wire N__17812;
    wire N__17809;
    wire N__17806;
    wire N__17803;
    wire N__17798;
    wire N__17795;
    wire N__17792;
    wire N__17789;
    wire N__17786;
    wire N__17783;
    wire N__17782;
    wire N__17779;
    wire N__17776;
    wire N__17773;
    wire N__17770;
    wire N__17765;
    wire N__17764;
    wire N__17761;
    wire N__17758;
    wire N__17755;
    wire N__17752;
    wire N__17749;
    wire N__17746;
    wire N__17743;
    wire N__17738;
    wire N__17735;
    wire N__17732;
    wire N__17731;
    wire N__17730;
    wire N__17729;
    wire N__17728;
    wire N__17727;
    wire N__17724;
    wire N__17723;
    wire N__17722;
    wire N__17715;
    wire N__17714;
    wire N__17713;
    wire N__17710;
    wire N__17709;
    wire N__17706;
    wire N__17705;
    wire N__17702;
    wire N__17699;
    wire N__17696;
    wire N__17695;
    wire N__17692;
    wire N__17689;
    wire N__17686;
    wire N__17685;
    wire N__17682;
    wire N__17677;
    wire N__17674;
    wire N__17671;
    wire N__17668;
    wire N__17665;
    wire N__17662;
    wire N__17659;
    wire N__17656;
    wire N__17653;
    wire N__17650;
    wire N__17645;
    wire N__17636;
    wire N__17621;
    wire N__17620;
    wire N__17617;
    wire N__17614;
    wire N__17613;
    wire N__17612;
    wire N__17611;
    wire N__17610;
    wire N__17605;
    wire N__17602;
    wire N__17599;
    wire N__17598;
    wire N__17595;
    wire N__17594;
    wire N__17593;
    wire N__17592;
    wire N__17589;
    wire N__17584;
    wire N__17581;
    wire N__17578;
    wire N__17575;
    wire N__17572;
    wire N__17569;
    wire N__17566;
    wire N__17565;
    wire N__17562;
    wire N__17559;
    wire N__17552;
    wire N__17549;
    wire N__17544;
    wire N__17541;
    wire N__17538;
    wire N__17525;
    wire N__17524;
    wire N__17521;
    wire N__17518;
    wire N__17513;
    wire N__17510;
    wire N__17509;
    wire N__17506;
    wire N__17503;
    wire N__17502;
    wire N__17501;
    wire N__17500;
    wire N__17497;
    wire N__17494;
    wire N__17491;
    wire N__17490;
    wire N__17485;
    wire N__17484;
    wire N__17483;
    wire N__17476;
    wire N__17473;
    wire N__17470;
    wire N__17467;
    wire N__17464;
    wire N__17461;
    wire N__17456;
    wire N__17447;
    wire N__17446;
    wire N__17445;
    wire N__17444;
    wire N__17441;
    wire N__17438;
    wire N__17437;
    wire N__17436;
    wire N__17433;
    wire N__17432;
    wire N__17431;
    wire N__17428;
    wire N__17423;
    wire N__17420;
    wire N__17417;
    wire N__17414;
    wire N__17411;
    wire N__17408;
    wire N__17405;
    wire N__17402;
    wire N__17397;
    wire N__17394;
    wire N__17381;
    wire N__17380;
    wire N__17377;
    wire N__17376;
    wire N__17373;
    wire N__17370;
    wire N__17365;
    wire N__17360;
    wire N__17357;
    wire N__17354;
    wire N__17351;
    wire N__17348;
    wire N__17345;
    wire N__17342;
    wire N__17339;
    wire N__17336;
    wire N__17333;
    wire N__17330;
    wire N__17327;
    wire N__17324;
    wire N__17321;
    wire N__17318;
    wire N__17315;
    wire N__17314;
    wire N__17311;
    wire N__17308;
    wire N__17303;
    wire N__17302;
    wire N__17301;
    wire N__17300;
    wire N__17299;
    wire N__17294;
    wire N__17291;
    wire N__17290;
    wire N__17289;
    wire N__17286;
    wire N__17285;
    wire N__17282;
    wire N__17279;
    wire N__17276;
    wire N__17273;
    wire N__17270;
    wire N__17267;
    wire N__17264;
    wire N__17261;
    wire N__17254;
    wire N__17247;
    wire N__17242;
    wire N__17239;
    wire N__17234;
    wire N__17231;
    wire N__17228;
    wire N__17225;
    wire N__17222;
    wire N__17221;
    wire N__17218;
    wire N__17217;
    wire N__17214;
    wire N__17209;
    wire N__17206;
    wire N__17201;
    wire N__17198;
    wire N__17195;
    wire N__17192;
    wire N__17189;
    wire N__17186;
    wire N__17185;
    wire N__17182;
    wire N__17179;
    wire N__17176;
    wire N__17173;
    wire N__17170;
    wire N__17167;
    wire N__17164;
    wire N__17161;
    wire N__17156;
    wire N__17153;
    wire N__17150;
    wire N__17149;
    wire N__17146;
    wire N__17143;
    wire N__17140;
    wire N__17137;
    wire N__17134;
    wire N__17131;
    wire N__17128;
    wire N__17125;
    wire N__17120;
    wire N__17117;
    wire N__17114;
    wire N__17111;
    wire N__17108;
    wire N__17105;
    wire N__17104;
    wire N__17101;
    wire N__17098;
    wire N__17095;
    wire N__17092;
    wire N__17087;
    wire N__17084;
    wire N__17081;
    wire N__17078;
    wire N__17075;
    wire N__17072;
    wire N__17069;
    wire N__17066;
    wire N__17063;
    wire N__17060;
    wire N__17057;
    wire N__17056;
    wire N__17055;
    wire N__17054;
    wire N__17049;
    wire N__17048;
    wire N__17047;
    wire N__17046;
    wire N__17043;
    wire N__17042;
    wire N__17041;
    wire N__17038;
    wire N__17035;
    wire N__17028;
    wire N__17021;
    wire N__17012;
    wire N__17011;
    wire N__17010;
    wire N__17009;
    wire N__17006;
    wire N__17001;
    wire N__17000;
    wire N__16999;
    wire N__16998;
    wire N__16997;
    wire N__16996;
    wire N__16995;
    wire N__16992;
    wire N__16987;
    wire N__16982;
    wire N__16973;
    wire N__16964;
    wire N__16961;
    wire N__16958;
    wire N__16955;
    wire N__16952;
    wire N__16949;
    wire N__16946;
    wire N__16943;
    wire N__16940;
    wire N__16937;
    wire N__16934;
    wire N__16931;
    wire N__16928;
    wire N__16925;
    wire N__16922;
    wire N__16919;
    wire N__16916;
    wire N__16913;
    wire N__16910;
    wire N__16907;
    wire N__16906;
    wire N__16905;
    wire N__16904;
    wire N__16903;
    wire N__16902;
    wire N__16901;
    wire N__16898;
    wire N__16893;
    wire N__16890;
    wire N__16887;
    wire N__16882;
    wire N__16879;
    wire N__16876;
    wire N__16865;
    wire N__16862;
    wire N__16859;
    wire N__16856;
    wire N__16853;
    wire N__16852;
    wire N__16849;
    wire N__16848;
    wire N__16847;
    wire N__16844;
    wire N__16843;
    wire N__16842;
    wire N__16839;
    wire N__16836;
    wire N__16833;
    wire N__16828;
    wire N__16825;
    wire N__16824;
    wire N__16823;
    wire N__16822;
    wire N__16821;
    wire N__16816;
    wire N__16813;
    wire N__16810;
    wire N__16807;
    wire N__16800;
    wire N__16797;
    wire N__16794;
    wire N__16789;
    wire N__16784;
    wire N__16775;
    wire N__16772;
    wire N__16769;
    wire N__16766;
    wire N__16763;
    wire N__16760;
    wire N__16757;
    wire N__16756;
    wire N__16753;
    wire N__16752;
    wire N__16749;
    wire N__16748;
    wire N__16747;
    wire N__16746;
    wire N__16745;
    wire N__16744;
    wire N__16741;
    wire N__16738;
    wire N__16735;
    wire N__16728;
    wire N__16727;
    wire N__16724;
    wire N__16721;
    wire N__16716;
    wire N__16711;
    wire N__16708;
    wire N__16703;
    wire N__16700;
    wire N__16697;
    wire N__16688;
    wire N__16685;
    wire N__16682;
    wire N__16679;
    wire N__16676;
    wire N__16673;
    wire N__16670;
    wire N__16667;
    wire N__16664;
    wire N__16661;
    wire N__16658;
    wire N__16655;
    wire N__16652;
    wire N__16649;
    wire N__16646;
    wire N__16643;
    wire N__16640;
    wire N__16639;
    wire N__16638;
    wire N__16633;
    wire N__16632;
    wire N__16631;
    wire N__16630;
    wire N__16629;
    wire N__16628;
    wire N__16627;
    wire N__16624;
    wire N__16621;
    wire N__16618;
    wire N__16615;
    wire N__16612;
    wire N__16609;
    wire N__16606;
    wire N__16603;
    wire N__16596;
    wire N__16583;
    wire N__16580;
    wire N__16577;
    wire N__16574;
    wire N__16571;
    wire N__16568;
    wire N__16565;
    wire N__16562;
    wire N__16559;
    wire N__16556;
    wire N__16553;
    wire N__16550;
    wire N__16547;
    wire N__16544;
    wire N__16541;
    wire N__16540;
    wire N__16537;
    wire N__16536;
    wire N__16533;
    wire N__16530;
    wire N__16527;
    wire N__16524;
    wire N__16517;
    wire N__16514;
    wire N__16511;
    wire N__16508;
    wire N__16505;
    wire N__16502;
    wire N__16501;
    wire N__16500;
    wire N__16499;
    wire N__16498;
    wire N__16495;
    wire N__16494;
    wire N__16491;
    wire N__16488;
    wire N__16485;
    wire N__16482;
    wire N__16479;
    wire N__16476;
    wire N__16475;
    wire N__16474;
    wire N__16473;
    wire N__16470;
    wire N__16465;
    wire N__16458;
    wire N__16453;
    wire N__16450;
    wire N__16447;
    wire N__16442;
    wire N__16439;
    wire N__16430;
    wire N__16429;
    wire N__16426;
    wire N__16425;
    wire N__16424;
    wire N__16423;
    wire N__16420;
    wire N__16417;
    wire N__16414;
    wire N__16411;
    wire N__16410;
    wire N__16409;
    wire N__16408;
    wire N__16407;
    wire N__16404;
    wire N__16399;
    wire N__16394;
    wire N__16387;
    wire N__16384;
    wire N__16379;
    wire N__16376;
    wire N__16373;
    wire N__16364;
    wire N__16363;
    wire N__16362;
    wire N__16359;
    wire N__16358;
    wire N__16355;
    wire N__16354;
    wire N__16351;
    wire N__16350;
    wire N__16347;
    wire N__16344;
    wire N__16341;
    wire N__16340;
    wire N__16339;
    wire N__16338;
    wire N__16335;
    wire N__16332;
    wire N__16329;
    wire N__16326;
    wire N__16323;
    wire N__16320;
    wire N__16313;
    wire N__16306;
    wire N__16301;
    wire N__16296;
    wire N__16289;
    wire N__16286;
    wire N__16283;
    wire N__16280;
    wire N__16277;
    wire N__16274;
    wire N__16271;
    wire N__16268;
    wire N__16267;
    wire N__16266;
    wire N__16263;
    wire N__16260;
    wire N__16257;
    wire N__16250;
    wire N__16247;
    wire N__16246;
    wire N__16245;
    wire N__16242;
    wire N__16239;
    wire N__16236;
    wire N__16233;
    wire N__16230;
    wire N__16225;
    wire N__16220;
    wire N__16217;
    wire N__16216;
    wire N__16215;
    wire N__16212;
    wire N__16209;
    wire N__16206;
    wire N__16203;
    wire N__16200;
    wire N__16193;
    wire N__16190;
    wire N__16187;
    wire N__16184;
    wire N__16181;
    wire N__16178;
    wire N__16175;
    wire N__16172;
    wire N__16169;
    wire N__16166;
    wire N__16163;
    wire N__16160;
    wire N__16159;
    wire N__16156;
    wire N__16151;
    wire N__16150;
    wire N__16147;
    wire N__16144;
    wire N__16139;
    wire N__16136;
    wire N__16133;
    wire N__16130;
    wire N__16127;
    wire N__16124;
    wire N__16121;
    wire N__16118;
    wire N__16115;
    wire N__16112;
    wire N__16109;
    wire N__16106;
    wire N__16103;
    wire N__16100;
    wire N__16097;
    wire N__16094;
    wire N__16091;
    wire N__16088;
    wire N__16085;
    wire N__16082;
    wire N__16079;
    wire N__16076;
    wire N__16073;
    wire N__16072;
    wire N__16071;
    wire N__16068;
    wire N__16065;
    wire N__16062;
    wire N__16059;
    wire N__16056;
    wire N__16049;
    wire N__16046;
    wire N__16043;
    wire N__16040;
    wire N__16037;
    wire N__16034;
    wire N__16031;
    wire N__16028;
    wire N__16025;
    wire N__16022;
    wire N__16019;
    wire N__16016;
    wire N__16015;
    wire N__16012;
    wire N__16009;
    wire N__16004;
    wire N__16003;
    wire N__16002;
    wire N__15999;
    wire N__15994;
    wire N__15989;
    wire N__15986;
    wire N__15983;
    wire N__15980;
    wire N__15977;
    wire N__15976;
    wire N__15973;
    wire N__15970;
    wire N__15967;
    wire N__15964;
    wire N__15961;
    wire N__15958;
    wire N__15955;
    wire N__15952;
    wire N__15949;
    wire N__15946;
    wire N__15943;
    wire N__15940;
    wire N__15937;
    wire N__15934;
    wire N__15931;
    wire N__15928;
    wire N__15925;
    wire N__15922;
    wire N__15919;
    wire N__15916;
    wire N__15913;
    wire N__15910;
    wire N__15907;
    wire N__15904;
    wire N__15901;
    wire N__15898;
    wire N__15895;
    wire N__15892;
    wire N__15887;
    wire N__15884;
    wire N__15881;
    wire N__15878;
    wire N__15877;
    wire N__15876;
    wire N__15875;
    wire N__15872;
    wire N__15869;
    wire N__15866;
    wire N__15863;
    wire N__15860;
    wire N__15859;
    wire N__15854;
    wire N__15849;
    wire N__15848;
    wire N__15845;
    wire N__15842;
    wire N__15839;
    wire N__15834;
    wire N__15827;
    wire N__15826;
    wire N__15825;
    wire N__15824;
    wire N__15821;
    wire N__15818;
    wire N__15813;
    wire N__15808;
    wire N__15807;
    wire N__15802;
    wire N__15801;
    wire N__15798;
    wire N__15795;
    wire N__15792;
    wire N__15789;
    wire N__15782;
    wire N__15779;
    wire N__15778;
    wire N__15775;
    wire N__15774;
    wire N__15773;
    wire N__15770;
    wire N__15767;
    wire N__15764;
    wire N__15761;
    wire N__15758;
    wire N__15755;
    wire N__15752;
    wire N__15749;
    wire N__15744;
    wire N__15741;
    wire N__15734;
    wire N__15731;
    wire N__15730;
    wire N__15729;
    wire N__15726;
    wire N__15725;
    wire N__15722;
    wire N__15719;
    wire N__15716;
    wire N__15713;
    wire N__15710;
    wire N__15707;
    wire N__15704;
    wire N__15699;
    wire N__15696;
    wire N__15693;
    wire N__15690;
    wire N__15683;
    wire N__15682;
    wire N__15681;
    wire N__15678;
    wire N__15675;
    wire N__15674;
    wire N__15671;
    wire N__15668;
    wire N__15665;
    wire N__15662;
    wire N__15659;
    wire N__15654;
    wire N__15649;
    wire N__15646;
    wire N__15641;
    wire N__15638;
    wire N__15635;
    wire N__15634;
    wire N__15631;
    wire N__15628;
    wire N__15625;
    wire N__15622;
    wire N__15617;
    wire N__15616;
    wire N__15613;
    wire N__15610;
    wire N__15609;
    wire N__15606;
    wire N__15603;
    wire N__15600;
    wire N__15599;
    wire N__15598;
    wire N__15597;
    wire N__15596;
    wire N__15593;
    wire N__15588;
    wire N__15585;
    wire N__15582;
    wire N__15577;
    wire N__15566;
    wire N__15565;
    wire N__15564;
    wire N__15561;
    wire N__15558;
    wire N__15555;
    wire N__15552;
    wire N__15549;
    wire N__15548;
    wire N__15547;
    wire N__15546;
    wire N__15543;
    wire N__15538;
    wire N__15533;
    wire N__15530;
    wire N__15529;
    wire N__15526;
    wire N__15521;
    wire N__15518;
    wire N__15515;
    wire N__15506;
    wire N__15503;
    wire N__15502;
    wire N__15501;
    wire N__15500;
    wire N__15499;
    wire N__15496;
    wire N__15495;
    wire N__15492;
    wire N__15487;
    wire N__15484;
    wire N__15481;
    wire N__15478;
    wire N__15477;
    wire N__15474;
    wire N__15471;
    wire N__15468;
    wire N__15463;
    wire N__15460;
    wire N__15455;
    wire N__15450;
    wire N__15443;
    wire N__15440;
    wire N__15437;
    wire N__15434;
    wire N__15431;
    wire N__15428;
    wire N__15425;
    wire N__15422;
    wire N__15419;
    wire N__15416;
    wire N__15413;
    wire N__15410;
    wire N__15409;
    wire N__15406;
    wire N__15403;
    wire N__15398;
    wire N__15397;
    wire N__15396;
    wire N__15393;
    wire N__15392;
    wire N__15387;
    wire N__15384;
    wire N__15381;
    wire N__15378;
    wire N__15377;
    wire N__15376;
    wire N__15371;
    wire N__15368;
    wire N__15363;
    wire N__15356;
    wire N__15353;
    wire N__15352;
    wire N__15349;
    wire N__15346;
    wire N__15345;
    wire N__15344;
    wire N__15343;
    wire N__15342;
    wire N__15337;
    wire N__15332;
    wire N__15327;
    wire N__15320;
    wire N__15319;
    wire N__15316;
    wire N__15313;
    wire N__15310;
    wire N__15307;
    wire N__15306;
    wire N__15305;
    wire N__15302;
    wire N__15299;
    wire N__15294;
    wire N__15287;
    wire N__15284;
    wire N__15281;
    wire N__15280;
    wire N__15277;
    wire N__15274;
    wire N__15273;
    wire N__15272;
    wire N__15271;
    wire N__15266;
    wire N__15263;
    wire N__15262;
    wire N__15257;
    wire N__15254;
    wire N__15251;
    wire N__15248;
    wire N__15239;
    wire N__15238;
    wire N__15237;
    wire N__15236;
    wire N__15233;
    wire N__15230;
    wire N__15227;
    wire N__15226;
    wire N__15225;
    wire N__15220;
    wire N__15215;
    wire N__15212;
    wire N__15209;
    wire N__15200;
    wire N__15199;
    wire N__15198;
    wire N__15197;
    wire N__15194;
    wire N__15193;
    wire N__15190;
    wire N__15187;
    wire N__15184;
    wire N__15181;
    wire N__15178;
    wire N__15175;
    wire N__15172;
    wire N__15171;
    wire N__15166;
    wire N__15163;
    wire N__15158;
    wire N__15155;
    wire N__15152;
    wire N__15147;
    wire N__15140;
    wire N__15139;
    wire N__15136;
    wire N__15133;
    wire N__15132;
    wire N__15127;
    wire N__15124;
    wire N__15123;
    wire N__15122;
    wire N__15121;
    wire N__15118;
    wire N__15115;
    wire N__15108;
    wire N__15101;
    wire N__15098;
    wire N__15095;
    wire N__15092;
    wire N__15089;
    wire N__15088;
    wire N__15087;
    wire N__15084;
    wire N__15081;
    wire N__15078;
    wire N__15073;
    wire N__15068;
    wire N__15065;
    wire N__15062;
    wire N__15059;
    wire N__15056;
    wire N__15053;
    wire N__15050;
    wire N__15047;
    wire N__15044;
    wire N__15043;
    wire N__15042;
    wire N__15041;
    wire N__15038;
    wire N__15035;
    wire N__15030;
    wire N__15023;
    wire N__15020;
    wire N__15019;
    wire N__15018;
    wire N__15017;
    wire N__15014;
    wire N__15007;
    wire N__15002;
    wire N__14999;
    wire N__14996;
    wire N__14993;
    wire N__14990;
    wire N__14987;
    wire N__14984;
    wire N__14981;
    wire N__14978;
    wire N__14975;
    wire N__14972;
    wire N__14969;
    wire N__14966;
    wire N__14963;
    wire N__14960;
    wire N__14957;
    wire N__14954;
    wire N__14951;
    wire N__14948;
    wire N__14945;
    wire N__14942;
    wire N__14939;
    wire N__14936;
    wire N__14933;
    wire N__14930;
    wire N__14927;
    wire N__14924;
    wire N__14921;
    wire N__14918;
    wire N__14915;
    wire N__14912;
    wire N__14909;
    wire N__14906;
    wire N__14903;
    wire N__14900;
    wire N__14897;
    wire N__14896;
    wire N__14895;
    wire N__14892;
    wire N__14889;
    wire N__14886;
    wire N__14881;
    wire N__14876;
    wire N__14875;
    wire N__14872;
    wire N__14869;
    wire N__14866;
    wire N__14865;
    wire N__14864;
    wire N__14861;
    wire N__14858;
    wire N__14853;
    wire N__14846;
    wire N__14843;
    wire N__14840;
    wire N__14837;
    wire N__14834;
    wire N__14833;
    wire N__14832;
    wire N__14825;
    wire N__14822;
    wire N__14819;
    wire N__14816;
    wire N__14813;
    wire N__14812;
    wire N__14811;
    wire N__14808;
    wire N__14803;
    wire N__14800;
    wire N__14797;
    wire N__14792;
    wire N__14791;
    wire N__14790;
    wire N__14789;
    wire N__14788;
    wire N__14787;
    wire N__14786;
    wire N__14785;
    wire N__14784;
    wire N__14783;
    wire N__14780;
    wire N__14779;
    wire N__14778;
    wire N__14777;
    wire N__14774;
    wire N__14771;
    wire N__14768;
    wire N__14765;
    wire N__14762;
    wire N__14755;
    wire N__14754;
    wire N__14753;
    wire N__14752;
    wire N__14751;
    wire N__14740;
    wire N__14737;
    wire N__14734;
    wire N__14731;
    wire N__14726;
    wire N__14723;
    wire N__14714;
    wire N__14711;
    wire N__14708;
    wire N__14705;
    wire N__14698;
    wire N__14687;
    wire N__14684;
    wire N__14683;
    wire N__14680;
    wire N__14677;
    wire N__14674;
    wire N__14671;
    wire N__14666;
    wire N__14663;
    wire N__14660;
    wire N__14657;
    wire N__14654;
    wire N__14651;
    wire N__14648;
    wire N__14645;
    wire N__14642;
    wire N__14641;
    wire N__14640;
    wire N__14637;
    wire N__14632;
    wire N__14629;
    wire N__14626;
    wire N__14621;
    wire N__14618;
    wire N__14617;
    wire N__14616;
    wire N__14613;
    wire N__14610;
    wire N__14607;
    wire N__14604;
    wire N__14601;
    wire N__14594;
    wire N__14591;
    wire N__14590;
    wire N__14587;
    wire N__14584;
    wire N__14583;
    wire N__14580;
    wire N__14577;
    wire N__14574;
    wire N__14571;
    wire N__14568;
    wire N__14561;
    wire N__14558;
    wire N__14557;
    wire N__14554;
    wire N__14551;
    wire N__14548;
    wire N__14543;
    wire N__14540;
    wire N__14539;
    wire N__14536;
    wire N__14533;
    wire N__14528;
    wire N__14525;
    wire N__14522;
    wire N__14519;
    wire N__14516;
    wire N__14513;
    wire N__14510;
    wire N__14507;
    wire N__14504;
    wire N__14501;
    wire N__14498;
    wire N__14495;
    wire N__14492;
    wire N__14489;
    wire N__14486;
    wire N__14483;
    wire N__14480;
    wire N__14477;
    wire N__14474;
    wire N__14471;
    wire N__14468;
    wire N__14465;
    wire N__14462;
    wire N__14459;
    wire N__14456;
    wire N__14453;
    wire N__14452;
    wire N__14449;
    wire N__14446;
    wire N__14443;
    wire N__14440;
    wire N__14437;
    wire N__14434;
    wire N__14431;
    wire N__14428;
    wire N__14425;
    wire N__14422;
    wire N__14419;
    wire N__14416;
    wire N__14413;
    wire N__14410;
    wire N__14407;
    wire N__14404;
    wire N__14401;
    wire N__14398;
    wire N__14395;
    wire N__14392;
    wire N__14389;
    wire N__14386;
    wire N__14383;
    wire N__14380;
    wire N__14377;
    wire N__14374;
    wire N__14371;
    wire N__14368;
    wire N__14365;
    wire N__14360;
    wire N__14357;
    wire N__14356;
    wire N__14353;
    wire N__14350;
    wire N__14347;
    wire N__14344;
    wire N__14341;
    wire N__14338;
    wire N__14335;
    wire N__14332;
    wire N__14329;
    wire N__14326;
    wire N__14323;
    wire N__14320;
    wire N__14317;
    wire N__14314;
    wire N__14311;
    wire N__14308;
    wire N__14305;
    wire N__14302;
    wire N__14299;
    wire N__14296;
    wire N__14293;
    wire N__14290;
    wire N__14287;
    wire N__14284;
    wire N__14281;
    wire N__14278;
    wire N__14275;
    wire N__14272;
    wire N__14269;
    wire N__14264;
    wire N__14263;
    wire N__14260;
    wire N__14257;
    wire N__14254;
    wire N__14251;
    wire N__14248;
    wire N__14245;
    wire N__14242;
    wire N__14239;
    wire N__14236;
    wire N__14233;
    wire N__14230;
    wire N__14227;
    wire N__14224;
    wire N__14221;
    wire N__14218;
    wire N__14215;
    wire N__14212;
    wire N__14209;
    wire N__14206;
    wire N__14203;
    wire N__14200;
    wire N__14197;
    wire N__14194;
    wire N__14191;
    wire N__14188;
    wire N__14185;
    wire N__14182;
    wire N__14179;
    wire N__14176;
    wire N__14171;
    wire N__14170;
    wire N__14167;
    wire N__14164;
    wire N__14161;
    wire N__14158;
    wire N__14155;
    wire N__14152;
    wire N__14149;
    wire N__14146;
    wire N__14143;
    wire N__14140;
    wire N__14137;
    wire N__14134;
    wire N__14131;
    wire N__14128;
    wire N__14125;
    wire N__14122;
    wire N__14119;
    wire N__14116;
    wire N__14113;
    wire N__14110;
    wire N__14107;
    wire N__14104;
    wire N__14101;
    wire N__14098;
    wire N__14095;
    wire N__14092;
    wire N__14089;
    wire N__14086;
    wire N__14081;
    wire N__14078;
    wire N__14075;
    wire N__14072;
    wire N__14069;
    wire N__14068;
    wire N__14063;
    wire N__14060;
    wire N__14057;
    wire N__14054;
    wire N__14051;
    wire N__14048;
    wire N__14045;
    wire N__14042;
    wire N__14039;
    wire N__14036;
    wire N__14033;
    wire N__14032;
    wire N__14029;
    wire N__14026;
    wire N__14021;
    wire N__14018;
    wire N__14015;
    wire N__14012;
    wire N__14009;
    wire N__14008;
    wire N__14005;
    wire N__14002;
    wire N__13997;
    wire N__13994;
    wire N__13991;
    wire N__13988;
    wire N__13987;
    wire N__13982;
    wire N__13979;
    wire N__13976;
    wire N__13973;
    wire N__13970;
    wire N__13969;
    wire N__13964;
    wire N__13961;
    wire N__13958;
    wire N__13955;
    wire N__13952;
    wire N__13949;
    wire N__13948;
    wire N__13945;
    wire N__13942;
    wire N__13937;
    wire N__13934;
    wire N__13931;
    wire N__13928;
    wire N__13925;
    wire N__13922;
    wire N__13919;
    wire N__13918;
    wire N__13915;
    wire N__13914;
    wire N__13907;
    wire N__13904;
    wire N__13901;
    wire N__13898;
    wire N__13895;
    wire N__13892;
    wire N__13889;
    wire N__13886;
    wire N__13883;
    wire N__13880;
    wire N__13877;
    wire N__13874;
    wire N__13871;
    wire N__13868;
    wire N__13865;
    wire N__13862;
    wire N__13859;
    wire N__13856;
    wire N__13853;
    wire N__13852;
    wire N__13851;
    wire N__13850;
    wire N__13849;
    wire N__13848;
    wire N__13847;
    wire N__13846;
    wire N__13845;
    wire N__13844;
    wire N__13823;
    wire N__13820;
    wire N__13817;
    wire N__13814;
    wire N__13811;
    wire N__13808;
    wire N__13805;
    wire N__13802;
    wire N__13801;
    wire N__13798;
    wire N__13795;
    wire N__13790;
    wire N__13787;
    wire N__13784;
    wire N__13781;
    wire N__13778;
    wire N__13775;
    wire N__13774;
    wire N__13771;
    wire N__13768;
    wire N__13763;
    wire N__13760;
    wire N__13759;
    wire N__13758;
    wire N__13755;
    wire N__13752;
    wire N__13749;
    wire N__13748;
    wire N__13747;
    wire N__13744;
    wire N__13743;
    wire N__13740;
    wire N__13737;
    wire N__13732;
    wire N__13729;
    wire N__13726;
    wire N__13721;
    wire N__13712;
    wire N__13709;
    wire N__13706;
    wire N__13703;
    wire N__13700;
    wire N__13697;
    wire N__13694;
    wire N__13691;
    wire N__13690;
    wire N__13689;
    wire N__13682;
    wire N__13679;
    wire N__13676;
    wire N__13675;
    wire N__13672;
    wire N__13671;
    wire N__13664;
    wire N__13661;
    wire N__13658;
    wire N__13657;
    wire N__13656;
    wire N__13655;
    wire N__13652;
    wire N__13645;
    wire N__13642;
    wire N__13639;
    wire N__13634;
    wire N__13631;
    wire N__13630;
    wire N__13627;
    wire N__13624;
    wire N__13621;
    wire N__13616;
    wire N__13613;
    wire N__13612;
    wire N__13609;
    wire N__13606;
    wire N__13605;
    wire N__13602;
    wire N__13597;
    wire N__13592;
    wire N__13589;
    wire N__13586;
    wire N__13583;
    wire N__13580;
    wire N__13577;
    wire N__13574;
    wire N__13571;
    wire N__13568;
    wire N__13565;
    wire N__13562;
    wire N__13559;
    wire N__13556;
    wire N__13553;
    wire N__13550;
    wire N__13547;
    wire N__13544;
    wire N__13541;
    wire N__13538;
    wire N__13535;
    wire N__13532;
    wire N__13529;
    wire N__13526;
    wire N__13523;
    wire N__13520;
    wire N__13517;
    wire N__13514;
    wire N__13511;
    wire N__13508;
    wire N__13505;
    wire N__13502;
    wire N__13499;
    wire N__13496;
    wire N__13493;
    wire N__13490;
    wire N__13487;
    wire N__13484;
    wire N__13481;
    wire N__13478;
    wire N__13475;
    wire N__13472;
    wire N__13469;
    wire N__13466;
    wire N__13465;
    wire N__13462;
    wire N__13459;
    wire N__13454;
    wire N__13451;
    wire N__13448;
    wire N__13445;
    wire N__13444;
    wire N__13441;
    wire N__13438;
    wire N__13433;
    wire N__13430;
    wire N__13427;
    wire N__13424;
    wire N__13421;
    wire N__13418;
    wire N__13415;
    wire N__13412;
    wire N__13409;
    wire N__13406;
    wire N__13403;
    wire N__13400;
    wire N__13397;
    wire N__13394;
    wire N__13393;
    wire N__13392;
    wire N__13389;
    wire N__13384;
    wire N__13379;
    wire N__13376;
    wire N__13375;
    wire N__13374;
    wire N__13371;
    wire N__13368;
    wire N__13365;
    wire N__13362;
    wire N__13355;
    wire N__13352;
    wire N__13349;
    wire N__13346;
    wire N__13343;
    wire N__13340;
    wire N__13337;
    wire N__13334;
    wire N__13331;
    wire N__13328;
    wire N__13325;
    wire N__13322;
    wire N__13319;
    wire N__13316;
    wire N__13313;
    wire N__13310;
    wire N__13307;
    wire N__13304;
    wire N__13301;
    wire N__13298;
    wire N__13295;
    wire N__13292;
    wire N__13289;
    wire N__13286;
    wire N__13283;
    wire N__13280;
    wire N__13277;
    wire N__13274;
    wire N__13271;
    wire N__13268;
    wire N__13265;
    wire N__13262;
    wire N__13259;
    wire N__13256;
    wire N__13253;
    wire N__13250;
    wire N__13247;
    wire N__13244;
    wire N__13241;
    wire N__13238;
    wire N__13235;
    wire N__13232;
    wire N__13229;
    wire N__13226;
    wire N__13223;
    wire N__13220;
    wire N__13217;
    wire N__13214;
    wire N__13211;
    wire N__13208;
    wire N__13205;
    wire N__13202;
    wire N__13199;
    wire N__13196;
    wire N__13193;
    wire N__13190;
    wire N__13187;
    wire N__13184;
    wire N__13181;
    wire N__13178;
    wire N__13175;
    wire N__13172;
    wire N__13169;
    wire N__13166;
    wire N__13163;
    wire N__13162;
    wire N__13161;
    wire N__13156;
    wire N__13153;
    wire N__13148;
    wire N__13145;
    wire N__13142;
    wire N__13141;
    wire N__13140;
    wire N__13133;
    wire N__13130;
    wire N__13129;
    wire N__13126;
    wire N__13125;
    wire N__13122;
    wire N__13115;
    wire N__13112;
    wire N__13109;
    wire N__13106;
    wire N__13103;
    wire N__13100;
    wire N__13097;
    wire N__13096;
    wire N__13095;
    wire N__13088;
    wire N__13085;
    wire VCCG0;
    wire GNDG0;
    wire \b2v_inst.N_4_i_i_a3_0_0_cascade_ ;
    wire \b2v_inst.un4_pix_count_intlto6_d_1_1_cascade_ ;
    wire b2v_inst4_pix_count_int_fast_1;
    wire b2v_inst4_pix_count_int_fast_0;
    wire \b2v_inst.N_13 ;
    wire b2v_inst4_pix_count_int_fast_2;
    wire b2v_inst4_pix_count_int_fast_3;
    wire \b2v_inst.pix_count_anteriorZ0Z_1 ;
    wire \b2v_inst.pix_count_anteriorZ0Z_4 ;
    wire \b2v_inst.un7_pix_count_int_0_I_1_c_RNOZ0 ;
    wire bfn_2_11_0_;
    wire \b2v_inst.un7_pix_count_int_0_data_tmp_0 ;
    wire \b2v_inst.un7_pix_count_int_0_I_15_c_RNOZ0 ;
    wire \b2v_inst.un7_pix_count_int_0_data_tmp_1 ;
    wire \b2v_inst.un7_pix_count_int_0_data_tmp_2 ;
    wire \b2v_inst.un7_pix_count_int_0_data_tmp_3 ;
    wire \b2v_inst.un7_pix_count_int_0_data_tmp_4 ;
    wire \b2v_inst.un7_pix_count_int_0_data_tmp_5 ;
    wire \b2v_inst.un7_pix_count_int_0_data_tmp_6 ;
    wire \b2v_inst.un7_pix_count_int_0_data_tmp_7 ;
    wire bfn_2_12_0_;
    wire \b2v_inst.un7_pix_count_int_0_data_tmp_8 ;
    wire \b2v_inst.un7_pix_count_int_0_N_2 ;
    wire \b2v_inst.un7_pix_count_int_0_I_57_c_RNOZ0 ;
    wire \b2v_inst4.un1_pix_count_int_0_sqmuxa_6 ;
    wire \b2v_inst.un7_pix_count_int_0_I_27_c_RNOZ0 ;
    wire \b2v_inst.pix_count_anteriorZ0Z_2 ;
    wire \b2v_inst.pix_count_anteriorZ0Z_3 ;
    wire \b2v_inst.pix_count_anteriorZ0Z_0 ;
    wire \b2v_inst.pix_count_anteriorZ0Z_5 ;
    wire \b2v_inst.un7_pix_count_int_0_I_33_c_RNOZ0 ;
    wire \b2v_inst.pix_count_anteriorZ0Z_18 ;
    wire \b2v_inst.un7_pix_count_int_0_I_39_c_RNOZ0 ;
    wire \b2v_inst.pix_count_anteriorZ0Z_12 ;
    wire \b2v_inst.pix_count_anteriorZ0Z_13 ;
    wire \b2v_inst.un7_pix_count_int_0_I_45_c_RNOZ0 ;
    wire \b2v_inst.pix_count_anteriorZ0Z_14 ;
    wire \b2v_inst4.un1_pix_count_int_0_sqmuxa_5_cascade_ ;
    wire \b2v_inst.pix_count_anteriorZ0Z_15 ;
    wire \b2v_inst.pix_count_anteriorZ0Z_19 ;
    wire \b2v_inst.pix_count_anteriorZ0Z_16 ;
    wire \b2v_inst.un1_state_36_0_a2_0_2_1_cascade_ ;
    wire \b2v_inst.N_305_2 ;
    wire \b2v_inst.N_305_2_cascade_ ;
    wire \b2v_inst.cuenta_pixelZ0Z_1 ;
    wire bfn_3_10_0_;
    wire \b2v_inst.un1_cuenta_pixel_cry_1 ;
    wire \b2v_inst.un1_cuenta_pixel_cry_2 ;
    wire \b2v_inst.un1_cuenta_pixel_cry_3 ;
    wire \b2v_inst.un1_cuenta_pixel_cry_4 ;
    wire \b2v_inst.cuenta_pixelZ0Z_6 ;
    wire \b2v_inst.un1_cuenta_pixel_cry_5_c_RNIGL1IZ0 ;
    wire \b2v_inst.un1_cuenta_pixel_cry_5 ;
    wire \b2v_inst.cuenta_pixelZ0Z_7 ;
    wire \b2v_inst.un1_cuenta_pixel_cry_6_c_RNIIO2IZ0 ;
    wire \b2v_inst.un1_cuenta_pixel_cry_6 ;
    wire \b2v_inst.cuenta_pixelZ0Z_8 ;
    wire \b2v_inst.un1_cuenta_pixel_cry_7 ;
    wire \b2v_inst.un1_cuenta_pixel_cry_8 ;
    wire \b2v_inst.cuenta_pixelZ0Z_9 ;
    wire bfn_3_11_0_;
    wire \b2v_inst.un1_cuenta_pixel_cry_9 ;
    wire \b2v_inst.cuenta_pixelZ0Z_10 ;
    wire \b2v_inst.pix_count_anteriorZ0Z_9 ;
    wire \b2v_inst.un7_pix_count_int_0_I_51_c_RNOZ0 ;
    wire \b2v_inst.N_1_0_0_cascade_ ;
    wire \b2v_inst.N_4_i_i_o6_2_cascade_ ;
    wire \b2v_inst.N_7 ;
    wire \b2v_inst.un7_pix_count_int_0_I_21_c_RNOZ0 ;
    wire \b2v_inst.pix_count_anteriorZ0Z_6 ;
    wire \b2v_inst.pix_count_anteriorZ0Z_7 ;
    wire \b2v_inst.pix_count_anteriorZ0Z_8 ;
    wire \b2v_inst4.un1_pix_count_int_0_sqmuxa_7 ;
    wire \b2v_inst4.un1_pix_count_int_0_sqmuxa_13 ;
    wire \b2v_inst4.un1_pix_count_int_0_sqmuxa_8_cascade_ ;
    wire \b2v_inst4.un1_pix_count_int_0_sqmuxa_14 ;
    wire \b2v_inst4.un1_pix_count_int_0_sqmuxa_10 ;
    wire \b2v_inst.cuenta_pixel_RNIT0FMZ0Z_1 ;
    wire \b2v_inst.cuenta_pixelZ0Z_0 ;
    wire \b2v_inst.cuenta_pixel_5_i_a2_0_2_5_cascade_ ;
    wire \b2v_inst.cuenta_pixelZ0Z_2 ;
    wire \b2v_inst.cuenta_pixelZ0Z_3 ;
    wire \b2v_inst.un1_cuenta_pixel_cry_1_c_RNI89THZ0 ;
    wire \b2v_inst.un1_cuenta_pixel_cry_2_c_RNIACUHZ0 ;
    wire \b2v_inst.un1_cuenta_pixel_cry_4_c_RNIEI0IZ0 ;
    wire \b2v_inst.cuenta_pixel_5_i_a2_0_2_5 ;
    wire \b2v_inst.cuenta_pixel_5_i_a2_0_1_5 ;
    wire \b2v_inst.cuenta_pixelZ0Z_5 ;
    wire \b2v_inst.un1_cuenta_pixel_cry_3_c_RNICFVHZ0 ;
    wire \b2v_inst.cuenta_pixelZ0Z_4 ;
    wire \b2v_inst.un7_pix_count_int_0_I_9_c_RNOZ0 ;
    wire \b2v_inst.pix_count_anteriorZ0Z_10 ;
    wire \b2v_inst.pix_count_anteriorZ0Z_11 ;
    wire \b2v_inst.pix_count_anteriorZ0Z_17 ;
    wire \b2v_inst.N_305_1_g ;
    wire \b2v_inst.N_4_i_i_a6_1 ;
    wire \b2v_inst4.pix_count_int_RNI0EPTZ0Z_0 ;
    wire bfn_5_13_0_;
    wire \b2v_inst4.un1_pix_count_int_cry_0_c_RNIIC2IZ0 ;
    wire \b2v_inst4.un1_pix_count_int_cry_0 ;
    wire \b2v_inst4.un1_pix_count_int_cry_1_c_RNIKF3IZ0 ;
    wire \b2v_inst4.un1_pix_count_int_cry_1 ;
    wire \b2v_inst4.un1_pix_count_int_cry_2_c_RNIMI4IZ0 ;
    wire \b2v_inst4.un1_pix_count_int_cry_2 ;
    wire \b2v_inst4.un1_pix_count_int_cry_3 ;
    wire \b2v_inst4.un1_pix_count_int_cry_4_c_RNIQO6IZ0 ;
    wire \b2v_inst4.un1_pix_count_int_cry_4 ;
    wire \b2v_inst4.un1_pix_count_int_cry_5_c_RNISR7IZ0 ;
    wire \b2v_inst4.un1_pix_count_int_cry_5 ;
    wire \b2v_inst4.un1_pix_count_int_cry_6 ;
    wire \b2v_inst4.un1_pix_count_int_cry_7 ;
    wire bfn_5_14_0_;
    wire \b2v_inst4.un1_pix_count_int_cry_8 ;
    wire \b2v_inst4.un1_pix_count_int_cry_9 ;
    wire \b2v_inst4.un1_pix_count_int_cry_10 ;
    wire \b2v_inst4.un1_pix_count_int_cry_11_c_RNIMPVJZ0 ;
    wire \b2v_inst4.un1_pix_count_int_cry_11 ;
    wire \b2v_inst4.un1_pix_count_int_cry_12 ;
    wire \b2v_inst4.un1_pix_count_int_cry_13 ;
    wire \b2v_inst4.un1_pix_count_int_cry_14 ;
    wire \b2v_inst4.un1_pix_count_int_cry_15 ;
    wire bfn_5_15_0_;
    wire \b2v_inst4.un1_pix_count_int_cry_16 ;
    wire \b2v_inst4.un1_pix_count_int_cry_17 ;
    wire \b2v_inst4.un1_pix_count_int_cry_18 ;
    wire SYNTHESIZED_WIRE_12_1;
    wire SYNTHESIZED_WIRE_12_7;
    wire SYNTHESIZED_WIRE_12_0;
    wire SYNTHESIZED_WIRE_12_8;
    wire bfn_6_5_0_;
    wire \b2v_inst.un2_dir_mem_3_cry_0 ;
    wire \b2v_inst.un2_dir_mem_3_cry_1 ;
    wire \b2v_inst.un2_dir_mem_3_cry_2 ;
    wire \b2v_inst.un2_dir_mem_3_cry_3 ;
    wire \b2v_inst.un2_dir_mem_3_cry_4 ;
    wire bfn_6_6_0_;
    wire \b2v_inst.un1_indice_cry_1 ;
    wire \b2v_inst.un1_indice_cry_2 ;
    wire \b2v_inst.un1_indice_cry_3 ;
    wire \b2v_inst.un1_indice_cry_4 ;
    wire \b2v_inst.un1_indice_cry_5 ;
    wire \b2v_inst.un1_indice_cry_6 ;
    wire \b2v_inst.un1_indice_cry_7 ;
    wire \b2v_inst.un1_indice_cry_8 ;
    wire bfn_6_7_0_;
    wire \b2v_inst.un1_indice_cry_9 ;
    wire \b2v_inst.un1_indice_cry_10 ;
    wire \b2v_inst.ignorar_ancho_1_RNOZ0Z_1 ;
    wire \b2v_inst.ignorar_ancho_1_RNOZ0Z_2 ;
    wire \b2v_inst4.un1_pix_count_int_cry_9_c_RNIB86JZ0 ;
    wire \b2v_inst4.un1_pix_count_int_cry_8_c_RNI25BIZ0 ;
    wire \b2v_inst4.un1_pix_count_int_0_sqmuxa_0 ;
    wire \b2v_inst4.un1_pix_count_int_cry_10_c_RNIKMUJZ0 ;
    wire \b2v_inst.ignorar_ancho_1_RNOZ0Z_0 ;
    wire \b2v_inst.N_482_cascade_ ;
    wire \b2v_inst.un1_state_34_0 ;
    wire \b2v_inst.un1_cuenta_pixel_cry_8_c_RNIMU4IZ0 ;
    wire \b2v_inst.cuenta_pixel_RNIVBL9Z0Z_10 ;
    wire \b2v_inst.un1_cuenta_pixel_cry_7_c_RNIKR3IZ0 ;
    wire \b2v_inst.cuenta_pixel_5_i_a2_1_1_0_5 ;
    wire \b2v_inst.N_325 ;
    wire \b2v_inst.un1_state_36_0_rn_1 ;
    wire \b2v_inst.un1_state_36_0_sn ;
    wire \b2v_inst.N_325_cascade_ ;
    wire \b2v_inst.N_305_1 ;
    wire \b2v_inst.un1_state_36_0 ;
    wire \b2v_inst4.stateZ0Z_0 ;
    wire SYNTHESIZED_WIRE_9;
    wire \b2v_inst.un1_state_36_0_a2_0_1_mbZ0Z_1 ;
    wire \b2v_inst1.N_40 ;
    wire bfn_7_6_0_;
    wire \b2v_inst.un8_dir_mem_1_cry_0 ;
    wire \b2v_inst.un8_dir_mem_1_cry_1 ;
    wire \b2v_inst.un8_dir_mem_1_cry_2 ;
    wire \b2v_inst.un8_dir_mem_1_cry_3 ;
    wire \b2v_inst.un8_dir_mem_1_cry_4 ;
    wire \b2v_inst.un8_dir_mem_1_cry_5 ;
    wire \b2v_inst.un8_dir_mem_1_cry_6 ;
    wire \b2v_inst.un8_dir_mem_1_cry_7 ;
    wire bfn_7_7_0_;
    wire \b2v_inst.un8_dir_mem_1_cry_8 ;
    wire \b2v_inst.un8_dir_mem_1_cry_9 ;
    wire \b2v_inst.un8_dir_mem_1_cry_10 ;
    wire \b2v_inst.dir_mem_316lt6_0_cascade_ ;
    wire \b2v_inst.dir_mem_316lt7 ;
    wire \b2v_inst.un1_indice_cry_1_c_RNIUSJGZ0 ;
    wire SYNTHESIZED_WIRE_4_fast_10;
    wire SYNTHESIZED_WIRE_4_fast_9;
    wire \b2v_inst.N_9_cascade_ ;
    wire b2v_inst4_pix_count_int_fast_5;
    wire b2v_inst4_pix_count_int_fast_6;
    wire \b2v_inst.un4_pix_count_intlto6_1_xZ0Z1 ;
    wire \b2v_inst.un4_pix_count_intlto6_1_xZ0Z0 ;
    wire \b2v_inst.un4_pix_count_intlto6_dZ0Z_1 ;
    wire \b2v_inst.un4_pix_count_intlto10_1_0Z0Z_0 ;
    wire \b2v_inst.un4_pix_count_intlt8_cascade_ ;
    wire \b2v_inst.un4_pix_count_intlto15_1_aZ0Z0 ;
    wire \b2v_inst.un4_pix_count_intlt16 ;
    wire SYNTHESIZED_WIRE_4_12;
    wire SYNTHESIZED_WIRE_4_11;
    wire SYNTHESIZED_WIRE_4_9_rep1;
    wire \b2v_inst1.r_RX_Bytece_0_4_cascade_ ;
    wire \b2v_inst.un4_pix_count_intlto10_1_d_0_xZ0Z1_cascade_ ;
    wire SYNTHESIZED_WIRE_4_0;
    wire SYNTHESIZED_WIRE_4_3;
    wire SYNTHESIZED_WIRE_4_1;
    wire SYNTHESIZED_WIRE_4_2;
    wire SYNTHESIZED_WIRE_4_6;
    wire SYNTHESIZED_WIRE_4_5;
    wire \b2v_inst.un4_pix_count_intlto6_d_1_0_cascade_ ;
    wire SYNTHESIZED_WIRE_4_10_rep1;
    wire b2v_inst4_pix_count_int_fast_11;
    wire b2v_inst4_pix_count_int_fast_12;
    wire b2v_inst_un4_pix_count_intlto12_0;
    wire SYNTHESIZED_WIRE_4_10;
    wire SYNTHESIZED_WIRE_4_9;
    wire b2v_inst_un4_pix_count_intlto12_0_cascade_;
    wire SYNTHESIZED_WIRE_4_8;
    wire N_457_i;
    wire \b2v_inst1.N_48 ;
    wire \b2v_inst1.N_44_cascade_ ;
    wire \b2v_inst.N_8 ;
    wire \b2v_inst1.N_42 ;
    wire \b2v_inst1.r_SM_Main_d_4 ;
    wire \b2v_inst1.N_47 ;
    wire \b2v_inst1.r_SM_Main_d_4_cascade_ ;
    wire \b2v_inst1.N_51 ;
    wire SYNTHESIZED_WIRE_12_9;
    wire bfn_8_5_0_;
    wire \b2v_inst.un2_dir_mem_1_cry_0 ;
    wire \b2v_inst.un2_dir_mem_1_cry_1 ;
    wire \b2v_inst.un2_dir_mem_1_cry_2 ;
    wire \b2v_inst.un2_dir_mem_1_cry_3 ;
    wire \b2v_inst.un2_dir_mem_1_cry_4 ;
    wire \b2v_inst.un2_dir_mem_1_cry_5 ;
    wire \b2v_inst.un2_dir_mem_1_cry_6 ;
    wire \b2v_inst.un2_dir_mem_1_cry_7 ;
    wire bfn_8_6_0_;
    wire \b2v_inst.un2_dir_mem_1_cry_8 ;
    wire \b2v_inst.un1_indice_cry_10_THRU_CO ;
    wire \b2v_inst.dir_mem_3_RNO_0Z0Z_10 ;
    wire \b2v_inst.dir_mem_3_RNO_0Z0Z_7 ;
    wire \b2v_inst.dir_mem_3_RNO_0Z0Z_8 ;
    wire \b2v_inst.dir_mem_3_RNO_0Z0Z_9 ;
    wire \b2v_inst.un1_indice_cry_2_c_RNI00LGZ0 ;
    wire \b2v_inst.indice_RNIJFHBZ0Z_0 ;
    wire \b2v_inst.un1_indice_cry_5_c_RNI69OGZ0 ;
    wire \b2v_inst.dir_mem_3_RNO_0Z0Z_6 ;
    wire bfn_8_9_0_;
    wire \b2v_inst.un3_dir_mem_cry_0 ;
    wire \b2v_inst.un3_dir_mem_cry_1 ;
    wire \b2v_inst.un3_dir_mem_cry_2 ;
    wire \b2v_inst.un3_dir_mem_cry_3 ;
    wire \b2v_inst.un3_dir_mem_cry_4 ;
    wire \b2v_inst.un3_dir_mem_cry_5 ;
    wire \b2v_inst.un3_dir_mem_cry_6 ;
    wire \b2v_inst.un3_dir_mem_cry_7 ;
    wire bfn_8_10_0_;
    wire \b2v_inst.un3_dir_mem_cry_8 ;
    wire \b2v_inst.un3_dir_mem_cry_9 ;
    wire SYNTHESIZED_WIRE_4_13;
    wire SYNTHESIZED_WIRE_4_15;
    wire SYNTHESIZED_WIRE_4_14;
    wire \b2v_inst.state_RNO_25Z0Z_29 ;
    wire \b2v_inst.g2_1_0 ;
    wire \b2v_inst.m29_2_cascade_ ;
    wire \b2v_inst.un4_pix_count_intlto10_1_d_0 ;
    wire \b2v_inst1.N_96_cascade_ ;
    wire \b2v_inst.g0_0_i_a4Z0Z_0 ;
    wire \b2v_inst.g0_0_iZ0Z_2 ;
    wire \b2v_inst.g2Z0Z_1 ;
    wire \b2v_inst1.N_58_i_cascade_ ;
    wire \b2v_inst1.un22_r_clk_count_ac0_3 ;
    wire \b2v_inst1.r_RX_Bytece_0_6 ;
    wire \b2v_inst1.r_Clk_CountZ0Z_2 ;
    wire \b2v_inst1.m16_0_o2_cascade_ ;
    wire \b2v_inst.g0_1_0_0 ;
    wire SYNTHESIZED_WIRE_4_7;
    wire \b2v_inst.un4_pix_count_intlto6_d_1_2 ;
    wire SYNTHESIZED_WIRE_4_4;
    wire \b2v_inst.g1_0_0 ;
    wire \b2v_inst.g1_0_0Z0Z_2 ;
    wire \b2v_inst.g1_0_a4Z0Z_0 ;
    wire swit_c_9;
    wire \b2v_inst.addr_ram_energia_m0_9 ;
    wire \b2v_inst1.N_38_cascade_ ;
    wire \b2v_inst1.r_Bit_IndexZ0Z_2 ;
    wire \b2v_inst1.N_44 ;
    wire \b2v_inst1.N_36_cascade_ ;
    wire \b2v_inst1.r_Bit_IndexZ0Z_1 ;
    wire \b2v_inst1.r_Bit_IndexZ0Z_0 ;
    wire \b2v_inst1.N_50 ;
    wire \b2v_inst1.r_RX_Bytece_0_5 ;
    wire N_460_i;
    wire N_459_i;
    wire bfn_9_5_0_;
    wire \b2v_inst.un8_dir_mem_2_cry_1 ;
    wire \b2v_inst.un8_dir_mem_2_cry_2 ;
    wire \b2v_inst.un8_dir_mem_2_cry_3 ;
    wire \b2v_inst.un8_dir_mem_2_cry_4 ;
    wire \b2v_inst.un8_dir_mem_2_cry_5 ;
    wire \b2v_inst.un8_dir_mem_2_cry_6 ;
    wire \b2v_inst.un8_dir_mem_2_cry_7 ;
    wire \b2v_inst.un8_dir_mem_2_cry_8 ;
    wire bfn_9_6_0_;
    wire \b2v_inst.un8_dir_mem_2_cry_9 ;
    wire \b2v_inst.dir_mem_215lt6_0 ;
    wire leds_c_4;
    wire leds_c_5;
    wire \b2v_inst.dir_mem_115lt6_0 ;
    wire \b2v_inst.g0_1_0_cascade_ ;
    wire \b2v_inst.un7_pix_count_int_0_N_2_THRU_CO ;
    wire \b2v_inst.g0_6_cascade_ ;
    wire \b2v_inst.o2 ;
    wire \b2v_inst.G_40_i_6_cascade_ ;
    wire \b2v_inst.state_ns_i_0_a2_11_a2_0_3_3 ;
    wire \b2v_inst.N_618_5 ;
    wire \b2v_inst1.N_49 ;
    wire \b2v_inst1.r_RX_Byte_1_sqmuxa ;
    wire \b2v_inst.N_618_3 ;
    wire \b2v_inst.state_ns_i_0_a2_11_o2_4_0_3_3 ;
    wire \b2v_inst.un4_pix_count_intlto19_0_0 ;
    wire \b2v_inst.G_40_i_2 ;
    wire \b2v_inst.G_40_i_3 ;
    wire SYNTHESIZED_WIRE_4_19;
    wire SYNTHESIZED_WIRE_4_16;
    wire \b2v_inst.N_5 ;
    wire \b2v_inst.N_430_i_1_cascade_ ;
    wire SYNTHESIZED_WIRE_4_18;
    wire SYNTHESIZED_WIRE_4_17;
    wire \b2v_inst.g1Z0Z_0 ;
    wire \b2v_inst.pix_count_anterior5 ;
    wire \b2v_inst.state_ns_0_i_o2_6_23_cascade_ ;
    wire \b2v_inst.state_ns_0_i_o2_7_23 ;
    wire \b2v_inst.N_512_cascade_ ;
    wire \b2v_inst.N_430_tz ;
    wire \b2v_inst.g0_4_4_cascade_ ;
    wire \b2v_inst.g3_0_0 ;
    wire \b2v_inst.un4_pix_count_intlto18Z0Z_0 ;
    wire \b2v_inst.g0_0_cascade_ ;
    wire \b2v_inst.g3_0 ;
    wire \b2v_inst.g0_4_5 ;
    wire leds_c_10;
    wire leds_c_11;
    wire leds_c_7;
    wire \b2v_inst.un8_dir_mem_1_cry_2_c_RNI82QCZ0 ;
    wire \b2v_inst.un8_dir_mem_1_cry_3_c_RNIA5RCZ0 ;
    wire \b2v_inst.un8_dir_mem_1_cry_5_c_RNIEBTCZ0 ;
    wire \b2v_inst.dir_mem_1_RNO_0Z0Z_6 ;
    wire \b2v_inst.dir_mem_215lt7 ;
    wire \b2v_inst.dir_mem_115lt7 ;
    wire \b2v_inst.dir_mem_1_RNO_0Z0Z_10 ;
    wire \b2v_inst.dir_mem_115lt11_cascade_ ;
    wire \b2v_inst.dir_mem_115lto7 ;
    wire \b2v_inst.dir_mem_1_RNO_0Z0Z_7 ;
    wire \b2v_inst.un8_dir_mem_1_cry_7_c_RNIIHVCZ0 ;
    wire \b2v_inst.dir_mem_1_RNO_0Z0Z_8 ;
    wire \b2v_inst.un8_dir_mem_1_cry_8_c_RNIKK0DZ0 ;
    wire \b2v_inst.dir_mem_1_RNO_0Z0Z_9 ;
    wire \b2v_inst.un8_dir_mem_1_cry_4_c_RNIC8SCZ0 ;
    wire \b2v_inst.dir_mem_1_RNO_0Z0Z_5 ;
    wire \b2v_inst.dir_mem_1Z0Z_6 ;
    wire \b2v_inst.dir_mem_3Z0Z_6 ;
    wire \b2v_inst.dir_memZ0Z_7 ;
    wire \b2v_inst.N_450_i_1_cascade_ ;
    wire \b2v_inst.dir_memZ0Z_10 ;
    wire \b2v_inst.dir_mem_1Z0Z_5 ;
    wire \b2v_inst.dir_mem_3Z0Z_5 ;
    wire SYNTHESIZED_WIRE_1_5;
    wire \b2v_inst.dir_memZ0Z_4 ;
    wire \b2v_inst.addr_ram_iv_i_0_4_cascade_ ;
    wire indice_RNIN3333_4;
    wire \b2v_inst.dir_mem_1Z0Z_4 ;
    wire \b2v_inst.addr_ram_iv_i_1_4 ;
    wire \b2v_inst.un1_indice_cry_3_c_RNI23MGZ0 ;
    wire \b2v_inst.dir_mem_316lto11_0 ;
    wire \b2v_inst.dir_mem_316lt11 ;
    wire \b2v_inst.dir_mem_3Z0Z_4 ;
    wire \b2v_inst.N_362_i ;
    wire \b2v_inst.state_ns_0_i_a2_0_0_23 ;
    wire \b2v_inst.state_ns_i_0_a2_11_o2_4_0_6_1_3_cascade_ ;
    wire \b2v_inst.state_ns_i_0_a2_11_o2_4_0_1_3 ;
    wire \b2v_inst.N_11 ;
    wire \b2v_inst.N_4_i_i_1_cascade_ ;
    wire \b2v_inst.g3_i_1 ;
    wire swit_c_8;
    wire \b2v_inst.addr_ram_energia_m0_8 ;
    wire \b2v_inst.state_ns_i_0_a2_11_o2_4_0_5_3 ;
    wire \b2v_inst.state_RNO_2Z0Z_29 ;
    wire \b2v_inst.state_ns_i_0_a2_11_o2_4_0_7_3_cascade_ ;
    wire \b2v_inst.state_RNO_1Z0Z_29 ;
    wire \b2v_inst.dir_energia_RNO_0Z0Z_0 ;
    wire swit_c_6;
    wire \b2v_inst.addr_ram_energia_m0_6_cascade_ ;
    wire SYNTHESIZED_WIRE_12_6;
    wire swit_c_7;
    wire \b2v_inst.addr_ram_energia_m0_7 ;
    wire leds_c_12;
    wire \b2v_inst.un1_indice_cry_4_c_RNI46NGZ0 ;
    wire \b2v_inst.un1_indice_cry_8_c_RNICIRGZ0 ;
    wire \b2v_inst.dir_mem_316lto7 ;
    wire \b2v_inst.un8_dir_mem_2_cry_1_c_RNI88LLZ0 ;
    wire \b2v_inst.un8_dir_mem_2_cry_2_c_RNIABMLZ0 ;
    wire \b2v_inst.dir_mem_2Z0Z_4 ;
    wire \b2v_inst.un8_dir_mem_2_cry_3_c_RNICENLZ0 ;
    wire \b2v_inst.un8_dir_mem_2_cry_4_c_RNIEHOLZ0 ;
    wire \b2v_inst.un8_dir_mem_1_cry_10_THRU_CO ;
    wire \b2v_inst.un8_dir_mem_1_cry_9_c_RNITCOLZ0 ;
    wire \b2v_inst.dir_mem_1Z0Z_8 ;
    wire \b2v_inst.dir_mem_3Z0Z_8 ;
    wire \b2v_inst.dir_mem_3Z0Z_1 ;
    wire \b2v_inst.dir_memZ0Z_1 ;
    wire \b2v_inst.dir_mem_2Z0Z_1 ;
    wire \b2v_inst.un8_dir_mem_1_cry_0_c_RNI4SNCZ0 ;
    wire \b2v_inst.dir_mem_1Z0Z_1 ;
    wire \b2v_inst.dir_mem_115lt11 ;
    wire \b2v_inst.indice_RNILHHBZ0Z_2 ;
    wire \b2v_inst.dir_mem_115lto11_0 ;
    wire \b2v_inst.un8_dir_mem_1_cry_1_c_RNI6VOCZ0 ;
    wire \b2v_inst.N_363_i ;
    wire \b2v_inst.dir_mem_2Z0Z_6 ;
    wire \b2v_inst.N_489_cascade_ ;
    wire \b2v_inst.dir_mem_1Z0Z_7 ;
    wire \b2v_inst.dir_mem_3Z0Z_7 ;
    wire \b2v_inst.N_488_cascade_ ;
    wire \b2v_inst.addr_ram_iv_i_0_0_7 ;
    wire \b2v_inst.addr_ram_iv_i_0_1_7_cascade_ ;
    wire indice_RNI6J333_7;
    wire \b2v_inst.state_RNO_0Z0Z_29 ;
    wire \b2v_inst.dir_mem_1Z0Z_0 ;
    wire \b2v_inst.dir_mem_3Z0Z_0 ;
    wire \b2v_inst.dir_mem_2Z0Z_3 ;
    wire \b2v_inst.dir_memZ0Z_3 ;
    wire \b2v_inst.addr_ram_iv_i_0_0_3_cascade_ ;
    wire indice_RNIIU233_3;
    wire \b2v_inst.dir_mem_3Z0Z_3 ;
    wire \b2v_inst.dir_mem_1Z0Z_3 ;
    wire \b2v_inst.addr_ram_iv_i_0_1_3 ;
    wire \b2v_inst.dir_memZ0Z_0 ;
    wire \b2v_inst.N_618_6 ;
    wire \b2v_inst.N_514_cascade_ ;
    wire N_116_i;
    wire \b2v_inst.stateZ0Z_16 ;
    wire N_548_i;
    wire \b2v_inst.stateZ0Z_0 ;
    wire \b2v_inst.N_692_cascade_ ;
    wire \b2v_inst.N_477 ;
    wire swit_c_1;
    wire \b2v_inst.N_494_cascade_ ;
    wire \b2v_inst.addr_ram_energia_m0_1 ;
    wire SYNTHESIZED_WIRE_12_10;
    wire swit_c_2;
    wire \b2v_inst.addr_ram_energia_m0_2_cascade_ ;
    wire SYNTHESIZED_WIRE_12_2;
    wire swit_c_5;
    wire \b2v_inst.addr_ram_energia_m0_5_cascade_ ;
    wire SYNTHESIZED_WIRE_12_5;
    wire swit_c_10;
    wire \b2v_inst.addr_ram_energia_m0_10 ;
    wire swit_c_3;
    wire \b2v_inst.addr_ram_energia_m0_3_cascade_ ;
    wire SYNTHESIZED_WIRE_12_3;
    wire leds_c_6;
    wire swit_c_0;
    wire \b2v_inst.addr_ram_energia_m0_0 ;
    wire N_120_i;
    wire \b2v_inst.N_432_1_cascade_ ;
    wire \b2v_inst.un1_indice_cry_9_c_RNILAJPZ0 ;
    wire \b2v_inst.un1_indice_cry_7_c_RNIAFQGZ0 ;
    wire \b2v_inst.dir_mem_2Z0Z_0 ;
    wire \b2v_inst.un8_dir_mem_2_cry_9_THRU_CO ;
    wire \b2v_inst.un8_dir_mem_2_cry_8_c_RNITIJEZ0 ;
    wire \b2v_inst.dir_mem_2Z0Z_10 ;
    wire \b2v_inst.dir_mem_215lto7 ;
    wire \b2v_inst.dir_mem_2Z0Z_7 ;
    wire \b2v_inst.un8_dir_mem_2_cry_6_c_RNIINQZ0Z5 ;
    wire \b2v_inst.dir_mem_2Z0Z_8 ;
    wire \b2v_inst.un8_dir_mem_2_cry_7_c_RNIKQRZ0Z5 ;
    wire \b2v_inst.dir_mem_215lto11_0 ;
    wire \b2v_inst.dir_mem_215lt11 ;
    wire \b2v_inst.N_463_i ;
    wire \b2v_inst.indice_4_i_a2_0_7_3_1 ;
    wire \b2v_inst.N_432_1_tz ;
    wire N_556_i;
    wire \b2v_inst.indice_4_i_a2_0_7_2_1 ;
    wire N_117_i;
    wire \b2v_inst.dir_mem_1Z0Z_9 ;
    wire \b2v_inst.dir_mem_3Z0Z_9 ;
    wire N_554_i;
    wire \b2v_inst.dir_mem_2Z0Z_2 ;
    wire \b2v_inst.dir_memZ0Z_2 ;
    wire \b2v_inst.dir_mem_2Z0Z_9 ;
    wire \b2v_inst.dir_mem_1Z0Z_2 ;
    wire \b2v_inst.dir_mem_3Z0Z_2 ;
    wire \b2v_inst.N_829_cascade_ ;
    wire \b2v_inst.N_829 ;
    wire \b2v_inst.un1_state_23_i_a2_0_a2_0_a2_0_cascade_ ;
    wire \b2v_inst.stateZ0Z_22 ;
    wire \b2v_inst.stateZ0Z_26 ;
    wire \b2v_inst.un2_cuentalto10_i_a2_6 ;
    wire \b2v_inst1.m16_0_o2 ;
    wire \b2v_inst1.m16_0_a3_0_cascade_ ;
    wire \b2v_inst1.N_119 ;
    wire \b2v_inst1.r_Clk_Count_6_iv_0_a3_1_1_1_cascade_ ;
    wire \b2v_inst1.N_43 ;
    wire \b2v_inst1.r_Clk_Count_6_iv_0_0_1_cascade_ ;
    wire \b2v_inst1.r_Clk_CountZ0Z_0 ;
    wire \b2v_inst1.r_Clk_CountZ0Z_1 ;
    wire \b2v_inst.N_653_cascade_ ;
    wire \b2v_inst.stateZ0Z_17 ;
    wire \b2v_inst.state_ns_i_a2_1_15 ;
    wire \b2v_inst.cuenta_RNIKUJVZ0Z_0_cascade_ ;
    wire \b2v_inst.un20_cuentalto10_5_cascade_ ;
    wire \b2v_inst.un20_cuentalto10_sx ;
    wire \b2v_inst.un20_cuentalto10_sx_cascade_ ;
    wire \b2v_inst.state18_li_0_cascade_ ;
    wire N_130_i;
    wire \b2v_inst.N_512 ;
    wire \b2v_inst.stateZ0Z_30 ;
    wire \b2v_inst.N_828_cascade_ ;
    wire N_552_i;
    wire \b2v_inst.state_ns_0_i_o2_8_23 ;
    wire N_550_i;
    wire \b2v_inst.state_fastZ0Z_32 ;
    wire \b2v_inst.stateZ0Z_5 ;
    wire \b2v_inst.addr_ram_energia_ss0_0_i_o2_i_o2_0 ;
    wire \b2v_inst.dir_mem_RNO_0Z0Z_6 ;
    wire \b2v_inst.dir_memZ0Z_6 ;
    wire \b2v_inst.dir_mem_RNO_0Z0Z_8 ;
    wire \b2v_inst.dir_memZ0Z_8 ;
    wire \b2v_inst.dir_mem_RNO_0Z0Z_9 ;
    wire \b2v_inst.dir_memZ0Z_9 ;
    wire swit_c_4;
    wire \b2v_inst.N_494 ;
    wire \b2v_inst.N_247 ;
    wire \b2v_inst.addr_ram_energia_m0_4_cascade_ ;
    wire SYNTHESIZED_WIRE_12_4;
    wire uart_rx_i_c;
    wire \b2v_inst1.r_RX_Data_RZ0 ;
    wire \b2v_inst.un9_indice_0_a2_2 ;
    wire \b2v_inst.un9_indice_0_a2_3 ;
    wire \b2v_inst.dir_mem_RNO_0Z0Z_5 ;
    wire \b2v_inst.un9_indice_0_a2_2_cascade_ ;
    wire \b2v_inst.stateZ0Z_28 ;
    wire \b2v_inst.N_432_1 ;
    wire bfn_13_6_0_;
    wire \b2v_inst.N_442_i ;
    wire \b2v_inst.un2_dir_mem_2_cry_0_THRU_CO ;
    wire \b2v_inst.un2_dir_mem_2_cry_0 ;
    wire \b2v_inst.dir_mem_2_RNO_0Z0Z_2 ;
    wire \b2v_inst.un2_dir_mem_2_cry_1 ;
    wire \b2v_inst.dir_mem_2_RNO_0Z0Z_3 ;
    wire \b2v_inst.un2_dir_mem_2_cry_2 ;
    wire \b2v_inst.dir_mem_2_RNO_0Z0Z_4 ;
    wire \b2v_inst.un2_dir_mem_2_cry_3 ;
    wire \b2v_inst.dir_mem_2_RNO_0Z0Z_5 ;
    wire \b2v_inst.un2_dir_mem_2_cry_4 ;
    wire \b2v_inst.dir_mem_2_RNO_0Z0Z_6 ;
    wire \b2v_inst.un2_dir_mem_2_cry_5 ;
    wire \b2v_inst.dir_mem_2_RNO_0Z0Z_7 ;
    wire \b2v_inst.un2_dir_mem_2_cry_6 ;
    wire \b2v_inst.un2_dir_mem_2_cry_7 ;
    wire \b2v_inst.dir_mem_2_RNO_0Z0Z_8 ;
    wire bfn_13_7_0_;
    wire \b2v_inst.dir_mem_2_RNO_0Z0Z_9 ;
    wire \b2v_inst.un2_dir_mem_2_cry_8 ;
    wire \b2v_inst.un2_dir_mem_2_cry_9 ;
    wire \b2v_inst.dir_mem_2_RNO_0Z0Z_10 ;
    wire \b2v_inst1.r_SM_MainZ0Z_1 ;
    wire \b2v_inst1.r_RX_DataZ0 ;
    wire \b2v_inst1.r_SM_MainZ0Z_2 ;
    wire \b2v_inst1.m13_i_2 ;
    wire \b2v_inst1.N_95_cascade_ ;
    wire \b2v_inst1.N_96 ;
    wire \b2v_inst1.r_SM_MainZ0Z_0 ;
    wire \b2v_inst.dir_memZ0Z_5 ;
    wire \b2v_inst.N_450_i_1 ;
    wire \b2v_inst.dir_mem_2Z0Z_5 ;
    wire \b2v_inst.N_489 ;
    wire \b2v_inst9.data_to_send_10_0_0_0_5_cascade_ ;
    wire \b2v_inst9.data_to_sendZ0Z_5 ;
    wire \b2v_inst9.data_to_send_10_0_0_0_3_cascade_ ;
    wire \b2v_inst9.data_to_sendZ0Z_6 ;
    wire \b2v_inst.un1_data_a_escribir_0_sqmuxa_3_i_i_a2_0 ;
    wire \b2v_inst.N_655_cascade_ ;
    wire \b2v_inst.state18_li_0 ;
    wire \b2v_inst.cuenta_RNIR03AZ0Z_1 ;
    wire \b2v_inst.cuentaZ0Z_0 ;
    wire \b2v_inst.cuentaZ0Z_1 ;
    wire bfn_13_12_0_;
    wire \b2v_inst.cuentaZ0Z_2 ;
    wire \b2v_inst.un4_cuenta_cry_1_c_RNI9VZ0Z48 ;
    wire \b2v_inst.un4_cuenta_cry_1 ;
    wire \b2v_inst.cuentaZ0Z_3 ;
    wire \b2v_inst.un4_cuenta_cry_2_c_RNIBZ0Z268 ;
    wire \b2v_inst.un4_cuenta_cry_2 ;
    wire \b2v_inst.cuentaZ0Z_4 ;
    wire \b2v_inst.un4_cuenta_cry_3_c_RNIDZ0Z578 ;
    wire \b2v_inst.un4_cuenta_cry_3 ;
    wire \b2v_inst.un4_cuenta_cry_4 ;
    wire \b2v_inst.cuentaZ0Z_6 ;
    wire \b2v_inst.un4_cuenta_cry_5_c_RNIHBZ0Z98 ;
    wire \b2v_inst.un4_cuenta_cry_5 ;
    wire \b2v_inst.cuentaZ0Z_7 ;
    wire \b2v_inst.un4_cuenta_cry_6_c_RNIJEAZ0Z8 ;
    wire \b2v_inst.un4_cuenta_cry_6 ;
    wire \b2v_inst.cuentaZ0Z_8 ;
    wire \b2v_inst.un4_cuenta_cry_7_c_RNILHBZ0Z8 ;
    wire \b2v_inst.un4_cuenta_cry_7 ;
    wire \b2v_inst.un4_cuenta_cry_8 ;
    wire \b2v_inst.cuentaZ0Z_9 ;
    wire \b2v_inst.un4_cuenta_cry_8_c_RNINKCZ0Z8 ;
    wire bfn_13_13_0_;
    wire \b2v_inst.un4_cuenta_cry_9 ;
    wire N_458_i;
    wire b2v_inst_state_4;
    wire b2v_inst_state_8;
    wire leds_c_0;
    wire leds_c_1;
    wire leds_c_13;
    wire leds_c_2;
    wire leds_c_3;
    wire N_546_i;
    wire bfn_13_16_0_;
    wire \b2v_inst.dir_energia_s_1 ;
    wire \b2v_inst.dir_energia_cry_0 ;
    wire \b2v_inst.dir_energia_s_2 ;
    wire \b2v_inst.dir_energia_cry_1 ;
    wire \b2v_inst.dir_energia_s_3 ;
    wire \b2v_inst.dir_energia_cry_2 ;
    wire \b2v_inst.dir_energia_s_4 ;
    wire \b2v_inst.dir_energia_cry_3 ;
    wire \b2v_inst.dir_energia_s_5 ;
    wire \b2v_inst.dir_energia_cry_4 ;
    wire \b2v_inst.dir_energia_s_6 ;
    wire \b2v_inst.dir_energia_cry_5 ;
    wire \b2v_inst.dir_energia_s_7 ;
    wire \b2v_inst.dir_energia_cry_6 ;
    wire \b2v_inst.dir_energia_cry_7 ;
    wire \b2v_inst.dir_energia_s_8 ;
    wire bfn_13_17_0_;
    wire \b2v_inst.dir_energia_s_9 ;
    wire \b2v_inst.dir_energia_cry_8 ;
    wire \b2v_inst.dir_energia_s_10 ;
    wire \b2v_inst.dir_energia_cry_9 ;
    wire \b2v_inst.stateZ0Z_19 ;
    wire \b2v_inst.N_352_0 ;
    wire \b2v_inst.dir_energia_cry_10 ;
    wire \b2v_inst.dir_energiaZ0Z_11 ;
    wire \b2v_inst.N_430_i ;
    wire \b2v_inst.N_648_5 ;
    wire \b2v_inst.un9_indice_0_a2_5_1 ;
    wire \b2v_inst.un4_cuenta_cry_9_c_RNI01TZ0Z9 ;
    wire \b2v_inst.cuentaZ0Z_10 ;
    wire \b2v_inst.N_655 ;
    wire \b2v_inst.un4_cuenta_cry_4_c_RNIFZ0Z888 ;
    wire \b2v_inst.cuentaZ0Z_5 ;
    wire \b2v_inst.N_547_i_0 ;
    wire \b2v_inst9.data_to_send_10_0_0_0_4 ;
    wire \b2v_inst9.data_to_sendZ0Z_4 ;
    wire \b2v_inst9.data_to_send_10_0_0_1_4 ;
    wire \b2v_inst9.data_to_send_10_0_0_1_5 ;
    wire \b2v_inst9.fsm_state_ns_i_i_0_a2_2_2Z0Z_0 ;
    wire \b2v_inst9.N_583_cascade_ ;
    wire reset_c_i;
    wire \b2v_inst9.un2_n_fsm_state_0_sqmuxa_2_0_i_cascade_ ;
    wire \b2v_inst9.data_to_send_10_0_0_0_6 ;
    wire \b2v_inst9.data_to_send_10_0_0_0_7_cascade_ ;
    wire \b2v_inst9.data_to_sendZ0Z_7 ;
    wire \b2v_inst9.data_to_send_10_0_0_2_0 ;
    wire \b2v_inst9.data_to_send_10_0_0_1_0 ;
    wire \b2v_inst9.N_738_cascade_ ;
    wire \b2v_inst9.data_to_send_10_0_0_2_1 ;
    wire \b2v_inst9.data_to_sendZ0Z_1 ;
    wire N_478_cascade_;
    wire \b2v_inst9.data_to_send_10_0_0_0_0 ;
    wire b2v_inst_state_15;
    wire \b2v_inst9.N_832_cascade_ ;
    wire \b2v_inst9.data_to_send_10_0_0_0_1 ;
    wire \b2v_inst9.data_to_send_10_0_0_1_1 ;
    wire \b2v_inst9.data_to_send_10_0_0_2_2_cascade_ ;
    wire \b2v_inst9.data_to_sendZ0Z_2 ;
    wire \b2v_inst9.un2_n_fsm_state_0_sqmuxa_2_0_i_0 ;
    wire \b2v_inst9.N_740 ;
    wire \b2v_inst9.data_to_send_10_0_0_1_2 ;
    wire \b2v_inst9.N_738 ;
    wire \b2v_inst9.N_741 ;
    wire \b2v_inst9.data_to_send_10_0_0_1_3 ;
    wire b2v_inst_energia_temp_0;
    wire \b2v_inst.un14_data_ram_energia_o_axb_0 ;
    wire bfn_14_14_0_;
    wire b2v_inst_energia_temp_1;
    wire \b2v_inst.un14_data_ram_energia_o_cry_0_c_RNIEI4MZ0 ;
    wire \b2v_inst.un14_data_ram_energia_o_cry_0 ;
    wire b2v_inst_energia_temp_2;
    wire \b2v_inst.un14_data_ram_energia_o_cry_1_c_RNIHM5MZ0 ;
    wire \b2v_inst.un14_data_ram_energia_o_cry_1 ;
    wire b2v_inst_energia_temp_3;
    wire \b2v_inst.un14_data_ram_energia_o_cry_2_c_RNIKQ6MZ0 ;
    wire \b2v_inst.un14_data_ram_energia_o_cry_2 ;
    wire \b2v_inst.pix_data_regZ0Z_4 ;
    wire b2v_inst_energia_temp_4;
    wire \b2v_inst.un14_data_ram_energia_o_cry_3_c_RNINU7MZ0 ;
    wire \b2v_inst.un14_data_ram_energia_o_cry_3 ;
    wire b2v_inst_energia_temp_5;
    wire \b2v_inst.un14_data_ram_energia_o_cry_4_c_RNIQ29MZ0 ;
    wire \b2v_inst.un14_data_ram_energia_o_cry_4 ;
    wire b2v_inst_energia_temp_6;
    wire \b2v_inst.un14_data_ram_energia_o_cry_5_c_RNIT6AMZ0 ;
    wire \b2v_inst.un14_data_ram_energia_o_cry_5 ;
    wire b2v_inst_energia_temp_7;
    wire \b2v_inst.un14_data_ram_energia_o_cry_6_c_RNI0BBMZ0 ;
    wire \b2v_inst.un14_data_ram_energia_o_cry_6 ;
    wire \b2v_inst.un14_data_ram_energia_o_cry_7 ;
    wire \b2v_inst.un14_data_ram_energia_o_cry_7_c_RNIN84CZ0 ;
    wire bfn_14_15_0_;
    wire \b2v_inst.un14_data_ram_energia_o_cry_8_c_RNIPB5CZ0 ;
    wire \b2v_inst.un14_data_ram_energia_o_cry_8 ;
    wire b2v_inst_energia_temp_10;
    wire \b2v_inst.un14_data_ram_energia_o_cry_9 ;
    wire b2v_inst_energia_temp_11;
    wire SYNTHESIZED_WIRE_13_11;
    wire \b2v_inst.un14_data_ram_energia_o_cry_10 ;
    wire b2v_inst_energia_temp_12;
    wire SYNTHESIZED_WIRE_13_12;
    wire \b2v_inst.un14_data_ram_energia_o_cry_11 ;
    wire b2v_inst_energia_temp_13;
    wire \b2v_inst.un14_data_ram_energia_o_cry_12 ;
    wire SYNTHESIZED_WIRE_13_13;
    wire leds_c_8;
    wire b2v_inst_energia_temp_8;
    wire \b2v_inst.un14_data_ram_energia_o_cry_9_c_RNI28GBZ0 ;
    wire N_461_i;
    wire bfn_15_8_0_;
    wire \b2v_inst.data_a_escribir11_0 ;
    wire \b2v_inst.data_a_escribir11_2_and ;
    wire \b2v_inst.data_a_escribir11_1 ;
    wire \b2v_inst.data_a_escribir11_2 ;
    wire \b2v_inst.data_a_escribir11_4_and ;
    wire \b2v_inst.data_a_escribir11_3 ;
    wire \b2v_inst.data_a_escribir11_4 ;
    wire \b2v_inst.data_a_escribir11_5 ;
    wire \b2v_inst.data_a_escribir11_6 ;
    wire \b2v_inst.data_a_escribir11_7 ;
    wire bfn_15_9_0_;
    wire \b2v_inst.data_a_escribir11_8 ;
    wire \b2v_inst.data_a_escribir11_9 ;
    wire \b2v_inst.data_a_escribir12 ;
    wire \b2v_inst.data_a_escribir11_9_and ;
    wire \b2v_inst.data_a_escribir11_8_and ;
    wire \b2v_inst.dir_mem_1Z0Z_10 ;
    wire \b2v_inst.N_490 ;
    wire \b2v_inst.dir_mem_3Z0Z_10 ;
    wire \b2v_inst.N_488 ;
    wire bfn_15_10_0_;
    wire \b2v_inst.eventos_cry_0 ;
    wire \b2v_inst.eventos_cry_1 ;
    wire \b2v_inst.eventos_cry_2 ;
    wire \b2v_inst.eventos_cry_3 ;
    wire \b2v_inst.eventos_cry_4 ;
    wire \b2v_inst.eventos_cry_5 ;
    wire \b2v_inst.eventos_cry_6 ;
    wire \b2v_inst.eventos_cry_7 ;
    wire bfn_15_11_0_;
    wire \b2v_inst.eventos_cry_8 ;
    wire \b2v_inst.eventos_cry_9 ;
    wire \b2v_inst.state_ns_a3_i_0_a2_5_1 ;
    wire \b2v_inst.state_ns_a3_i_0_a2_4_1_cascade_ ;
    wire \b2v_inst.stateZ0Z_31 ;
    wire b2v_inst_state_7;
    wire b2v_inst_state_1;
    wire b2v_inst_state_2;
    wire \b2v_inst.stateZ0Z_11 ;
    wire \b2v_inst.stateZ0Z_32 ;
    wire b2v_inst_state_14;
    wire \b2v_inst.state_ns_a3_i_0_a2_6_1 ;
    wire \b2v_inst9.fsm_state_ns_i_0_i_0_1_cascade_ ;
    wire \b2v_inst9.N_832 ;
    wire \b2v_inst9.data_to_sendZ0Z_3 ;
    wire \b2v_inst9.data_to_send_10_0_0_0_2 ;
    wire b2v_inst_state_12;
    wire b2v_inst_state_13;
    wire \b2v_inst9.N_739 ;
    wire \b2v_inst.pix_data_regZ0Z_0 ;
    wire \b2v_inst.pix_data_regZ0Z_1 ;
    wire \b2v_inst.pix_data_regZ0Z_2 ;
    wire \b2v_inst.pix_data_regZ0Z_5 ;
    wire \b2v_inst.pix_data_regZ0Z_6 ;
    wire \b2v_inst.pix_data_regZ0Z_7 ;
    wire \b2v_inst9.N_583 ;
    wire leds_c_9;
    wire b2v_inst_energia_temp_9;
    wire \b2v_inst.N_577_i ;
    wire \b2v_inst9.data_to_sendZ0Z_0 ;
    wire uart_tx_o_c;
    wire \b2v_inst.reg_ancho_1_i_0 ;
    wire bfn_16_6_0_;
    wire \b2v_inst.reg_ancho_1_i_1 ;
    wire \b2v_inst.un2_valor_max1_cry_0 ;
    wire \b2v_inst.reg_ancho_1_i_2 ;
    wire \b2v_inst.un2_valor_max1_cry_1 ;
    wire \b2v_inst.reg_ancho_1_i_3 ;
    wire \b2v_inst.un2_valor_max1_cry_2 ;
    wire \b2v_inst.reg_ancho_1_i_4 ;
    wire \b2v_inst.un2_valor_max1_cry_3 ;
    wire \b2v_inst.reg_ancho_1_i_5 ;
    wire \b2v_inst.un2_valor_max1_cry_4 ;
    wire \b2v_inst.reg_ancho_1_i_6 ;
    wire \b2v_inst.un2_valor_max1_cry_5 ;
    wire \b2v_inst.reg_ancho_1_i_7 ;
    wire \b2v_inst.un2_valor_max1_cry_6 ;
    wire \b2v_inst.un2_valor_max1_cry_7 ;
    wire \b2v_inst.reg_ancho_1_i_8 ;
    wire bfn_16_7_0_;
    wire \b2v_inst.reg_ancho_1_i_9 ;
    wire \b2v_inst.un2_valor_max1_cry_8 ;
    wire \b2v_inst.reg_ancho_1_i_10 ;
    wire \b2v_inst.un2_valor_max1_cry_9 ;
    wire \b2v_inst.un2_valor_max1 ;
    wire \b2v_inst.ignorar_anchoZ0Z_1 ;
    wire \b2v_inst.stateZ0Z_25 ;
    wire \b2v_inst.data_a_escribir11_0_and ;
    wire \b2v_inst.eventosZ0Z_0 ;
    wire \b2v_inst.data_a_escribir_RNO_2Z0Z_0_cascade_ ;
    wire \b2v_inst.un1_reg_anterior_0_i_1_0_cascade_ ;
    wire \b2v_inst.eventosZ0Z_1 ;
    wire \b2v_inst.data_a_escribir_RNO_2Z0Z_1_cascade_ ;
    wire \b2v_inst.un1_reg_anterior_0_i_1_1_cascade_ ;
    wire \b2v_inst.eventosZ0Z_10 ;
    wire \b2v_inst.N_269 ;
    wire \b2v_inst.un1_reg_anterior_iv_0_0_10_cascade_ ;
    wire \b2v_inst.eventosZ0Z_6 ;
    wire \b2v_inst.un1_reg_anterior_iv_0_0_6_cascade_ ;
    wire \b2v_inst.N_272 ;
    wire \b2v_inst.data_a_escribir_1_sqmuxa ;
    wire \b2v_inst.data_a_escribir11_1_and ;
    wire \b2v_inst.eventosZ0Z_4 ;
    wire \b2v_inst.un1_reg_anterior_iv_0_0_4_cascade_ ;
    wire \b2v_inst.un1_reg_anterior_iv_0_1_4_cascade_ ;
    wire \b2v_inst.N_274 ;
    wire \b2v_inst.N_268 ;
    wire \b2v_inst.un1_reg_anterior_iv_0_1_10 ;
    wire SYNTHESIZED_WIRE_10_3;
    wire SYNTHESIZED_WIRE_10_4;
    wire SYNTHESIZED_WIRE_10_6;
    wire SYNTHESIZED_WIRE_10_7;
    wire SYNTHESIZED_WIRE_10_0;
    wire SYNTHESIZED_WIRE_5_0;
    wire SYNTHESIZED_WIRE_5_4;
    wire \b2v_inst.un12_pix_count_intlto7_N_2LZ0Z1_cascade_ ;
    wire \b2v_inst.un13_pix_count_int_li_0 ;
    wire \b2v_inst.un13_pix_count_int_li_0_cascade_ ;
    wire SYNTHESIZED_WIRE_10_1;
    wire SYNTHESIZED_WIRE_5_1;
    wire SYNTHESIZED_WIRE_10_2;
    wire SYNTHESIZED_WIRE_5_2;
    wire \b2v_inst.state_fastZ0Z_19 ;
    wire \b2v_inst9.fsm_state_srsts_1_0 ;
    wire \b2v_inst9.N_522 ;
    wire \b2v_inst9.N_522_cascade_ ;
    wire \b2v_inst9.fsm_stateZ0Z_0 ;
    wire \b2v_inst9.fsm_stateZ0Z_1 ;
    wire \b2v_inst9.N_84_2_cascade_ ;
    wire \b2v_inst9.N_582 ;
    wire bfn_17_5_0_;
    wire \b2v_inst.valor_max_final4_2_cry_0 ;
    wire \b2v_inst.valor_max_final4_2_cry_1 ;
    wire \b2v_inst.valor_max_final4_2_cry_2 ;
    wire \b2v_inst.valor_max_final4_2_cry_3 ;
    wire \b2v_inst.valor_max_final4_2_cry_4 ;
    wire \b2v_inst.valor_max_final4_2_cry_5 ;
    wire \b2v_inst.valor_max_final4_2_cry_6 ;
    wire \b2v_inst.valor_max_final4_2_cry_7 ;
    wire bfn_17_6_0_;
    wire \b2v_inst.valor_max_final4_2_cry_8 ;
    wire \b2v_inst.valor_max_final4_2_cry_9 ;
    wire \b2v_inst.valor_max_final42 ;
    wire \b2v_inst.data_a_escribir11_7_and ;
    wire SYNTHESIZED_WIRE_3_7;
    wire SYNTHESIZED_WIRE_3_8;
    wire SYNTHESIZED_WIRE_3_0;
    wire \b2v_inst.reg_ancho_2Z0Z_0 ;
    wire bfn_17_8_0_;
    wire \b2v_inst.valor_max_final4_3_cry_0 ;
    wire \b2v_inst.valor_max_final4_3_cry_1 ;
    wire \b2v_inst.valor_max_final4_3_cry_2 ;
    wire \b2v_inst.valor_max_final4_3_cry_3 ;
    wire \b2v_inst.reg_ancho_2Z0Z_5 ;
    wire \b2v_inst.valor_max_final4_3_cry_4 ;
    wire \b2v_inst.reg_ancho_2Z0Z_6 ;
    wire \b2v_inst.valor_max_final4_3_cry_5 ;
    wire \b2v_inst.reg_ancho_2Z0Z_7 ;
    wire \b2v_inst.valor_max_final4_3_cry_6 ;
    wire \b2v_inst.valor_max_final4_3_cry_7 ;
    wire bfn_17_9_0_;
    wire \b2v_inst.valor_max_final4_3_cry_8 ;
    wire \b2v_inst.valor_max_final4_3_cry_9 ;
    wire \b2v_inst.valor_max_final43 ;
    wire \b2v_inst.data_a_escribir_RNO_0Z0Z_0 ;
    wire \b2v_inst.data_a_escribir_RNO_0Z0Z_1 ;
    wire \b2v_inst.eventosZ0Z_5 ;
    wire \b2v_inst.reg_anterior_i_0 ;
    wire bfn_17_10_0_;
    wire \b2v_inst.reg_anterior_i_1 ;
    wire \b2v_inst.valor_max_final4_1_cry_0 ;
    wire \b2v_inst.reg_anterior_i_2 ;
    wire \b2v_inst.valor_max_final4_1_cry_1 ;
    wire \b2v_inst.reg_anterior_i_3 ;
    wire \b2v_inst.valor_max_final4_1_cry_2 ;
    wire \b2v_inst.reg_anterior_i_4 ;
    wire \b2v_inst.valor_max_final4_1_cry_3 ;
    wire \b2v_inst.reg_anterior_i_5 ;
    wire \b2v_inst.valor_max_final4_1_cry_4 ;
    wire \b2v_inst.reg_anterior_i_6 ;
    wire \b2v_inst.valor_max_final4_1_cry_5 ;
    wire \b2v_inst.reg_anterior_i_7 ;
    wire \b2v_inst.valor_max_final4_1_cry_6 ;
    wire \b2v_inst.valor_max_final4_1_cry_7 ;
    wire \b2v_inst.reg_anterior_i_8 ;
    wire bfn_17_11_0_;
    wire \b2v_inst.reg_anterior_i_9 ;
    wire \b2v_inst.valor_max_final4_1_cry_8 ;
    wire \b2v_inst.reg_anterior_i_10 ;
    wire \b2v_inst.valor_max_final4_1_cry_9 ;
    wire \b2v_inst.valor_max_final43_THRU_CO ;
    wire \b2v_inst.m54_ns_1 ;
    wire \b2v_inst.valor_max_final41 ;
    wire \b2v_inst.stateZ0Z_6 ;
    wire \b2v_inst.stateZ0Z_10 ;
    wire \b2v_inst.stateZ0Z_29 ;
    wire \b2v_inst.state_ns_a3_i_0_a2_1_4_1 ;
    wire b2v_inst_state_3;
    wire \b2v_inst.N_694 ;
    wire \b2v_inst.N_695_cascade_ ;
    wire \b2v_inst.state_ns_a3_i_0_1_1 ;
    wire \b2v_inst.un2_cuentalto10_i_a2_8 ;
    wire \b2v_inst.un2_cuentalto10_i_a2_7 ;
    wire \b2v_inst.state_32_repZ0Z1 ;
    wire reset_c;
    wire \b2v_inst.N_654_2 ;
    wire \b2v_inst.un1_reset_inv_0_0_tz_cascade_ ;
    wire \b2v_inst.N_482 ;
    wire \b2v_inst.eventosZ0Z_7 ;
    wire \b2v_inst.data_a_escribir_RNO_2Z0Z_7 ;
    wire bfn_17_13_0_;
    wire \b2v_inst9.un1_cycle_counter_2_cry_0 ;
    wire \b2v_inst9.un1_cycle_counter_2_cry_1 ;
    wire \b2v_inst9.un1_cycle_counter_2_cry_2 ;
    wire \b2v_inst9.cycle_counterZ0Z_3 ;
    wire \b2v_inst9.cycle_counter_RNIQAGDZ0Z_3_cascade_ ;
    wire \b2v_inst9.un1_cycle_counter_2_cry_0_THRU_CO ;
    wire \b2v_inst9.cycle_counterZ0Z_1 ;
    wire SYNTHESIZED_WIRE_5_7;
    wire SYNTHESIZED_WIRE_5_6;
    wire \b2v_inst.un12_pix_count_intlto7_N_3LZ0Z3 ;
    wire SYNTHESIZED_WIRE_10_5;
    wire SYNTHESIZED_WIRE_5_5;
    wire \b2v_inst4.pix_count_int_0_sqmuxa ;
    wire \b2v_inst9.N_175_i ;
    wire \b2v_inst9.bit_counterZ0Z_0 ;
    wire bfn_17_16_0_;
    wire \b2v_inst9.bit_counterZ1Z_1 ;
    wire \b2v_inst9.un1_bit_counter_3_cry_0 ;
    wire \b2v_inst9.bit_counterZ0Z_2 ;
    wire \b2v_inst9.un1_bit_counter_3_cry_1 ;
    wire \b2v_inst9.fsm_state_RNIND1P1Z0Z_0 ;
    wire \b2v_inst9.un1_bit_counter_3_cry_2 ;
    wire \b2v_inst9.bit_counterZ0Z_3 ;
    wire \b2v_inst.reg_anteriorZ0Z_0 ;
    wire bfn_18_6_0_;
    wire \b2v_inst.reg_anteriorZ0Z_1 ;
    wire \b2v_inst.un2_valor_max2_cry_0 ;
    wire \b2v_inst.un2_valor_max2_cry_1 ;
    wire \b2v_inst.un2_valor_max2_cry_2 ;
    wire \b2v_inst.un2_valor_max2_cry_3 ;
    wire \b2v_inst.un2_valor_max2_cry_4 ;
    wire \b2v_inst.un2_valor_max2_cry_5 ;
    wire \b2v_inst.un2_valor_max2_cry_6 ;
    wire \b2v_inst.un2_valor_max2_cry_7 ;
    wire bfn_18_7_0_;
    wire \b2v_inst.un2_valor_max2_cry_8 ;
    wire \b2v_inst.un2_valor_max2_cry_9 ;
    wire \b2v_inst.un2_valor_max2 ;
    wire \b2v_inst.reg_anteriorZ0Z_3 ;
    wire \b2v_inst.data_a_escribir_RNO_0Z0Z_3 ;
    wire \b2v_inst.reg_anteriorZ0Z_5 ;
    wire \b2v_inst.reg_ancho_1Z0Z_0 ;
    wire \b2v_inst.reg_ancho_3_i_0 ;
    wire bfn_18_8_0_;
    wire \b2v_inst.reg_ancho_1Z0Z_1 ;
    wire \b2v_inst.reg_ancho_3_i_1 ;
    wire \b2v_inst.valor_max_final4_0_cry_0 ;
    wire \b2v_inst.reg_ancho_3_i_2 ;
    wire \b2v_inst.valor_max_final4_0_cry_1 ;
    wire \b2v_inst.reg_ancho_3_i_3 ;
    wire \b2v_inst.valor_max_final4_0_cry_2 ;
    wire \b2v_inst.reg_ancho_1Z0Z_4 ;
    wire \b2v_inst.reg_ancho_3_i_4 ;
    wire \b2v_inst.valor_max_final4_0_cry_3 ;
    wire \b2v_inst.reg_ancho_1Z0Z_5 ;
    wire \b2v_inst.reg_ancho_3_i_5 ;
    wire \b2v_inst.valor_max_final4_0_cry_4 ;
    wire \b2v_inst.reg_ancho_1Z0Z_6 ;
    wire \b2v_inst.reg_ancho_3Z0Z_6 ;
    wire \b2v_inst.reg_ancho_3_i_6 ;
    wire \b2v_inst.valor_max_final4_0_cry_5 ;
    wire \b2v_inst.reg_ancho_1Z0Z_7 ;
    wire \b2v_inst.reg_ancho_3_i_7 ;
    wire \b2v_inst.valor_max_final4_0_cry_6 ;
    wire \b2v_inst.valor_max_final4_0_cry_7 ;
    wire \b2v_inst.reg_ancho_3_i_8 ;
    wire bfn_18_9_0_;
    wire \b2v_inst.reg_ancho_3_i_9 ;
    wire \b2v_inst.valor_max_final4_0_cry_8 ;
    wire \b2v_inst.reg_ancho_1Z0Z_10 ;
    wire \b2v_inst.reg_ancho_3_i_10 ;
    wire \b2v_inst.valor_max_final4_0_cry_9 ;
    wire \b2v_inst.valor_max_final40 ;
    wire \b2v_inst.valor_max_final40_THRU_CO ;
    wire \b2v_inst.reg_ancho_1Z0Z_9 ;
    wire \b2v_inst.reg_ancho_1Z0Z_8 ;
    wire \b2v_inst.reg_ancho_2Z0Z_8 ;
    wire \b2v_inst.eventosZ0Z_3 ;
    wire \b2v_inst.un1_reg_anterior_0_i_1_3 ;
    wire \b2v_inst.reg_anteriorZ0Z_2 ;
    wire \b2v_inst.data_a_escribir11_6_and ;
    wire \b2v_inst.N_273 ;
    wire \b2v_inst.un1_reg_anterior_iv_0_0_5 ;
    wire \b2v_inst.N_267 ;
    wire \b2v_inst.un1_reg_anterior_iv_0_1_5_cascade_ ;
    wire \b2v_inst.data_a_escribir_RNO_0Z0Z_2 ;
    wire \b2v_inst.reg_ancho_2Z0Z_9 ;
    wire \b2v_inst.reg_ancho_3Z0Z_1 ;
    wire \b2v_inst.reg_ancho_3Z0Z_0 ;
    wire \b2v_inst.data_a_escribir11_5_and ;
    wire \b2v_inst.reg_ancho_3Z0Z_9 ;
    wire \b2v_inst.eventosZ0Z_9 ;
    wire \b2v_inst.N_545 ;
    wire \b2v_inst.un1_reg_anterior_iv_0_0_0_9_cascade_ ;
    wire \b2v_inst.N_543 ;
    wire \b2v_inst.un1_reg_anterior_iv_0_0_1_9_cascade_ ;
    wire \b2v_inst.valor_max2_6 ;
    wire \b2v_inst.un1_reg_anterior_iv_0_1_6 ;
    wire \b2v_inst.data_a_escribir11_10_and ;
    wire \b2v_inst.eventosZ0Z_8 ;
    wire \b2v_inst.un1_reg_anterior_iv_0_0_0_8_cascade_ ;
    wire \b2v_inst.N_542 ;
    wire \b2v_inst.un1_reg_anterior_iv_0_0_1_8_cascade_ ;
    wire \b2v_inst.reg_anteriorZ0Z_8 ;
    wire \b2v_inst.reg_ancho_3Z0Z_8 ;
    wire \b2v_inst.N_544 ;
    wire \b2v_inst.reg_ancho_3Z0Z_7 ;
    wire \b2v_inst.reg_anteriorZ0Z_7 ;
    wire \b2v_inst.un1_reg_anterior_0_i_1_7 ;
    wire \b2v_inst.data_a_escribir_RNO_0Z0Z_7_cascade_ ;
    wire \b2v_inst.N_711 ;
    wire \b2v_inst.un1_reset_inv_0 ;
    wire \b2v_inst9.un1_cycle_counter_2_cry_1_THRU_CO ;
    wire \b2v_inst9.cycle_counterZ0Z_2 ;
    wire \b2v_inst9.cycle_counter_RNIQAGDZ0Z_3 ;
    wire N_478;
    wire \b2v_inst9.cycle_counterZ0Z_0 ;
    wire SYNTHESIZED_WIRE_5_3;
    wire \b2v_inst.pix_data_regZ0Z_3 ;
    wire \b2v_inst.stateZ0Z_24 ;
    wire SYNTHESIZED_WIRE_1_2;
    wire \b2v_inst.reg_anteriorZ0Z_4 ;
    wire SYNTHESIZED_WIRE_3_6;
    wire \b2v_inst.reg_anteriorZ0Z_6 ;
    wire \b2v_inst.reg_ancho_2Z0Z_10 ;
    wire \b2v_inst.reg_ancho_3Z0Z_4 ;
    wire \b2v_inst.data_a_escribir11_3_and ;
    wire SYNTHESIZED_WIRE_3_1;
    wire \b2v_inst.reg_ancho_2Z0Z_1 ;
    wire \b2v_inst.reg_ancho_2Z0Z_2 ;
    wire \b2v_inst.reg_ancho_1Z0Z_2 ;
    wire \b2v_inst.eventosZ0Z_2 ;
    wire \b2v_inst.data_a_escribir_RNO_2Z0Z_2_cascade_ ;
    wire \b2v_inst.data_a_escribir12_THRU_CO ;
    wire \b2v_inst.un1_reg_anterior_0_i_1_2 ;
    wire \b2v_inst.reg_ancho_1Z0Z_3 ;
    wire \b2v_inst.stateZ0Z_20 ;
    wire \b2v_inst.un2_valor_max1_THRU_CO ;
    wire \b2v_inst.data_a_escribir_RNO_2Z0Z_3 ;
    wire \b2v_inst.reg_ancho_2Z0Z_3 ;
    wire \b2v_inst.un2_valor_max2_THRU_CO ;
    wire \b2v_inst.N_264 ;
    wire \b2v_inst.reg_ancho_3Z0Z_10 ;
    wire SYNTHESIZED_WIRE_3_3;
    wire \b2v_inst.reg_ancho_3Z0Z_3 ;
    wire SYNTHESIZED_WIRE_3_2;
    wire \b2v_inst.reg_ancho_3Z0Z_2 ;
    wire SYNTHESIZED_WIRE_3_5;
    wire \b2v_inst.reg_ancho_3Z0Z_5 ;
    wire \b2v_inst.stateZ0Z_21 ;
    wire SYNTHESIZED_WIRE_3_9;
    wire \b2v_inst.reg_anteriorZ0Z_9 ;
    wire \b2v_inst.ignorar_anteriorZ0 ;
    wire SYNTHESIZED_WIRE_3_10;
    wire \b2v_inst.reg_anteriorZ0Z_10 ;
    wire \b2v_inst.stateZ0Z_27 ;
    wire SYNTHESIZED_WIRE_1_0;
    wire SYNTHESIZED_WIRE_1_1;
    wire SYNTHESIZED_WIRE_1_4;
    wire bfn_19_14_0_;
    wire b2v_inst_cantidad_temp_2;
    wire \b2v_inst.un16_data_ram_cantidad_o_cry_1 ;
    wire \b2v_inst.un16_data_ram_cantidad_o_cry_2 ;
    wire b2v_inst_cantidad_temp_4;
    wire \b2v_inst.un16_data_ram_cantidad_o_cry_3 ;
    wire b2v_inst_cantidad_temp_5;
    wire \b2v_inst.un16_data_ram_cantidad_o_cry_4 ;
    wire \b2v_inst.un16_data_ram_cantidad_o_cry_1_c_RNI77COZ0 ;
    wire N_553_i;
    wire \b2v_inst.un16_data_ram_cantidad_o_cry_3_c_RNIBDEOZ0 ;
    wire b2v_inst_data_a_escribir_4;
    wire N_549_i;
    wire \b2v_inst.un16_data_ram_cantidad_o_cry_2_c_RNI9ADOZ0 ;
    wire b2v_inst_data_a_escribir_3;
    wire N_551_i;
    wire \b2v_inst.N_481 ;
    wire N_121_i;
    wire b2v_inst_data_a_escribir_2;
    wire N_118_i;
    wire SYNTHESIZED_WIRE_3_4;
    wire \b2v_inst.reg_ancho_2Z0Z_4 ;
    wire \b2v_inst.stateZ0Z_23 ;
    wire b2v_inst_data_a_escribir_9;
    wire N_111_i;
    wire \b2v_inst.addr_ram_iv_i_1_6 ;
    wire \b2v_inst.addr_ram_iv_i_0_6 ;
    wire N_298;
    wire \b2v_inst.addr_ram_iv_i_0_5 ;
    wire \b2v_inst.addr_ram_iv_i_1_5 ;
    wire indice_RNIS8333_5;
    wire \b2v_inst.addr_ram_iv_i_0_8 ;
    wire \b2v_inst.addr_ram_iv_i_1_8 ;
    wire indice_RNIBO333_8;
    wire \b2v_inst.addr_ram_iv_i_0_9 ;
    wire \b2v_inst.addr_ram_iv_i_1_9 ;
    wire indice_RNIGT333_9;
    wire N_115_i;
    wire b2v_inst_data_a_escribir_10;
    wire N_110_i;
    wire \b2v_inst.addr_ram_iv_i_0_0 ;
    wire \b2v_inst.addr_ram_iv_i_1_0 ;
    wire indice_RNI3F233_0;
    wire \b2v_inst.addr_ram_iv_i_0_10 ;
    wire \b2v_inst.addr_ram_iv_i_1_10 ;
    wire N_37;
    wire b2v_inst_data_a_escribir_8;
    wire N_112_i;
    wire b2v_inst_data_a_escribir_7;
    wire N_113_i;
    wire \b2v_inst.addr_ram_iv_i_0_0_1 ;
    wire \b2v_inst.addr_ram_iv_i_0_1_1 ;
    wire indice_RNI8K233_1;
    wire b2v_inst_data_a_escribir_6;
    wire N_114_i;
    wire \b2v_inst.addr_ram_iv_i_0_2 ;
    wire \b2v_inst.N_480 ;
    wire \b2v_inst.addr_ram_iv_i_1_2 ;
    wire indice_RNIDP233_2;
    wire b2v_inst_data_a_escribir_0;
    wire N_557_i;
    wire b2v_inst_cantidad_temp_0;
    wire b2v_inst_cantidad_temp_1;
    wire b2v_inst_data_a_escribir_1;
    wire \b2v_inst.cantidad_temp_RNILL3KZ0Z_1_cascade_ ;
    wire N_555_i;
    wire \b2v_inst.stateZ0Z_18 ;
    wire SYNTHESIZED_WIRE_1_3;
    wire \b2v_inst.stateZ0Z_9 ;
    wire b2v_inst_cantidad_temp_3;
    wire clk_c_g;
    wire reset_c_i_g;
    wire \b2v_inst.N_828 ;
    wire \b2v_inst.un16_data_ram_cantidad_o_cry_4_c_RNIDGFOZ0 ;
    wire b2v_inst_data_a_escribir_5;
    wire \b2v_inst.N_514 ;
    wire N_547_i;
    wire CONSTANT_ONE_NET;
    wire \b2v_inst.dir_energiaZ0Z_10 ;
    wire \b2v_inst.indiceZ0Z_10 ;
    wire N_445_i;
    wire \b2v_inst.indiceZ0Z_3 ;
    wire \b2v_inst.dir_energiaZ0Z_3 ;
    wire N_357_i;
    wire \b2v_inst.indiceZ0Z_4 ;
    wire \b2v_inst.dir_energiaZ0Z_4 ;
    wire N_356_i;
    wire \b2v_inst.dir_energiaZ0Z_2 ;
    wire \b2v_inst.indiceZ0Z_2 ;
    wire N_358_i;
    wire \b2v_inst.indiceZ0Z_9 ;
    wire \b2v_inst.dir_energiaZ0Z_9 ;
    wire N_444_i;
    wire \b2v_inst.indiceZ0Z_5 ;
    wire \b2v_inst.dir_energiaZ0Z_5 ;
    wire N_355_i;
    wire \b2v_inst.dir_energiaZ0Z_0 ;
    wire \b2v_inst.indiceZ0Z_0 ;
    wire N_360_i;
    wire \b2v_inst.dir_energiaZ0Z_8 ;
    wire \b2v_inst.indiceZ0Z_8 ;
    wire N_443_i;
    wire \b2v_inst.dir_energiaZ0Z_7 ;
    wire \b2v_inst.indiceZ0Z_7 ;
    wire N_353_i;
    wire \b2v_inst.dir_energiaZ0Z_1 ;
    wire \b2v_inst.indiceZ0Z_1 ;
    wire N_359_i;
    wire \b2v_inst.N_645 ;
    wire \b2v_inst.dir_energiaZ0Z_6 ;
    wire \b2v_inst.indiceZ0Z_6 ;
    wire \b2v_inst.N_484 ;
    wire N_354_i;
    wire _gnd_net_;

    defparam \b2v_inst2.mem_mem_0_0_physical .WRITE_MODE=3;
    defparam \b2v_inst2.mem_mem_0_0_physical .READ_MODE=3;
    SB_RAM40_4K \b2v_inst2.mem_mem_0_0_physical  (
            .RDATA({dangling_wire_0,dangling_wire_1,dangling_wire_2,dangling_wire_3,SYNTHESIZED_WIRE_3_1,dangling_wire_4,dangling_wire_5,dangling_wire_6,dangling_wire_7,dangling_wire_8,dangling_wire_9,dangling_wire_10,SYNTHESIZED_WIRE_3_0,dangling_wire_11,dangling_wire_12,dangling_wire_13}),
            .RADDR({N__33476,N__33778,N__33892,N__19472,N__32785,N__34009,N__18469,N__19651,N__35057,N__35410,N__33590}),
            .WADDR({N__33475,N__33779,N__33893,N__19471,N__32786,N__34010,N__18473,N__19658,N__35056,N__35411,N__33589}),
            .MASK({dangling_wire_14,dangling_wire_15,dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29}),
            .WDATA({dangling_wire_30,dangling_wire_31,dangling_wire_32,dangling_wire_33,N__20372,dangling_wire_34,dangling_wire_35,dangling_wire_36,dangling_wire_37,dangling_wire_38,dangling_wire_39,dangling_wire_40,N__33146,dangling_wire_41,dangling_wire_42,dangling_wire_43}),
            .RCLKE(),
            .RCLK(N__34435),
            .RE(N__37212),
            .WCLKE(N__21473),
            .WCLK(N__34436),
            .WE(N__37292));
    defparam \b2v_inst8.mem_mem_0_0_physical .WRITE_MODE=3;
    defparam \b2v_inst8.mem_mem_0_0_physical .READ_MODE=3;
    SB_RAM40_4K \b2v_inst8.mem_mem_0_0_physical  (
            .RDATA({dangling_wire_44,dangling_wire_45,dangling_wire_46,dangling_wire_47,SYNTHESIZED_WIRE_1_1,dangling_wire_48,dangling_wire_49,dangling_wire_50,dangling_wire_51,dangling_wire_52,dangling_wire_53,dangling_wire_54,SYNTHESIZED_WIRE_1_0,dangling_wire_55,dangling_wire_56,dangling_wire_57}),
            .RADDR({N__36625,N__35770,N__38969,N__38756,N__38198,N__35548,N__36208,N__36421,N__35998,N__38510,N__39188}),
            .WADDR({N__36629,N__35771,N__38968,N__38755,N__38197,N__35549,N__36209,N__36422,N__35999,N__38509,N__39187}),
            .MASK({dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,dangling_wire_62,dangling_wire_63,dangling_wire_64,dangling_wire_65,dangling_wire_66,dangling_wire_67,dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71,dangling_wire_72,dangling_wire_73}),
            .WDATA({dangling_wire_74,dangling_wire_75,dangling_wire_76,dangling_wire_77,N__34772,dangling_wire_78,dangling_wire_79,dangling_wire_80,dangling_wire_81,dangling_wire_82,dangling_wire_83,dangling_wire_84,N__34916,dangling_wire_85,dangling_wire_86,dangling_wire_87}),
            .RCLKE(),
            .RCLK(N__34376),
            .RE(N__36996),
            .WCLKE(N__21453),
            .WCLK(N__34377),
            .WE(N__36847));
    defparam \b2v_inst7.mem_mem_0_2_physical .WRITE_MODE=3;
    defparam \b2v_inst7.mem_mem_0_2_physical .READ_MODE=3;
    SB_RAM40_4K \b2v_inst7.mem_mem_0_2_physical  (
            .RDATA({dangling_wire_88,dangling_wire_89,dangling_wire_90,dangling_wire_91,leds_c_5,dangling_wire_92,dangling_wire_93,dangling_wire_94,dangling_wire_95,dangling_wire_96,dangling_wire_97,dangling_wire_98,leds_c_4,dangling_wire_99,dangling_wire_100,dangling_wire_101}),
            .RADDR({N__20128,N__15955,N__14149,N__14332,N__18703,N__19879,N__21574,N__20512,N__19996,N__14428,N__14239}),
            .WADDR({N__20125,N__15952,N__14146,N__14341,N__18700,N__19876,N__21571,N__20509,N__19993,N__14431,N__14242}),
            .MASK({dangling_wire_102,dangling_wire_103,dangling_wire_104,dangling_wire_105,dangling_wire_106,dangling_wire_107,dangling_wire_108,dangling_wire_109,dangling_wire_110,dangling_wire_111,dangling_wire_112,dangling_wire_113,dangling_wire_114,dangling_wire_115,dangling_wire_116,dangling_wire_117}),
            .WDATA({dangling_wire_118,dangling_wire_119,dangling_wire_120,dangling_wire_121,N__23621,dangling_wire_122,dangling_wire_123,dangling_wire_124,dangling_wire_125,dangling_wire_126,dangling_wire_127,dangling_wire_128,N__19715,dangling_wire_129,dangling_wire_130,dangling_wire_131}),
            .RCLKE(),
            .RCLK(N__34486),
            .RE(N__37231),
            .WCLKE(N__21447),
            .WCLK(N__34487),
            .WE(N__37242));
    defparam \b2v_inst2.mem_mem_0_2_physical .WRITE_MODE=3;
    defparam \b2v_inst2.mem_mem_0_2_physical .READ_MODE=3;
    SB_RAM40_4K \b2v_inst2.mem_mem_0_2_physical  (
            .RDATA({dangling_wire_132,dangling_wire_133,dangling_wire_134,dangling_wire_135,SYNTHESIZED_WIRE_3_5,dangling_wire_136,dangling_wire_137,dangling_wire_138,dangling_wire_139,dangling_wire_140,dangling_wire_141,dangling_wire_142,SYNTHESIZED_WIRE_3_4,dangling_wire_143,dangling_wire_144,dangling_wire_145}),
            .RADDR({N__33454,N__33754,N__33868,N__19450,N__32761,N__33985,N__18445,N__19627,N__35035,N__35386,N__33568}),
            .WADDR({N__33451,N__33757,N__33871,N__19447,N__32764,N__33988,N__18454,N__19642,N__35032,N__35389,N__33565}),
            .MASK({dangling_wire_146,dangling_wire_147,dangling_wire_148,dangling_wire_149,dangling_wire_150,dangling_wire_151,dangling_wire_152,dangling_wire_153,dangling_wire_154,dangling_wire_155,dangling_wire_156,dangling_wire_157,dangling_wire_158,dangling_wire_159,dangling_wire_160,dangling_wire_161}),
            .WDATA({dangling_wire_162,dangling_wire_163,dangling_wire_164,dangling_wire_165,N__33698,dangling_wire_166,dangling_wire_167,dangling_wire_168,dangling_wire_169,dangling_wire_170,dangling_wire_171,dangling_wire_172,N__19754,dangling_wire_173,dangling_wire_174,dangling_wire_175}),
            .RCLKE(),
            .RCLK(N__34400),
            .RE(N__37129),
            .WCLKE(N__21468),
            .WCLK(N__34401),
            .WE(N__37198));
    defparam \b2v_inst2.mem_mem_0_1_physical .WRITE_MODE=3;
    defparam \b2v_inst2.mem_mem_0_1_physical .READ_MODE=3;
    SB_RAM40_4K \b2v_inst2.mem_mem_0_1_physical  (
            .RDATA({dangling_wire_176,dangling_wire_177,dangling_wire_178,dangling_wire_179,SYNTHESIZED_WIRE_3_3,dangling_wire_180,dangling_wire_181,dangling_wire_182,dangling_wire_183,dangling_wire_184,dangling_wire_185,dangling_wire_186,SYNTHESIZED_WIRE_3_2,dangling_wire_187,dangling_wire_188,dangling_wire_189}),
            .RADDR({N__33466,N__33766,N__33880,N__19462,N__32773,N__33997,N__18457,N__19639,N__35047,N__35398,N__33580}),
            .WADDR({N__33463,N__33769,N__33883,N__19459,N__32776,N__34000,N__18466,N__19652,N__35044,N__35401,N__33577}),
            .MASK({dangling_wire_190,dangling_wire_191,dangling_wire_192,dangling_wire_193,dangling_wire_194,dangling_wire_195,dangling_wire_196,dangling_wire_197,dangling_wire_198,dangling_wire_199,dangling_wire_200,dangling_wire_201,dangling_wire_202,dangling_wire_203,dangling_wire_204,dangling_wire_205}),
            .WDATA({dangling_wire_206,dangling_wire_207,dangling_wire_208,dangling_wire_209,N__20555,dangling_wire_210,dangling_wire_211,dangling_wire_212,dangling_wire_213,dangling_wire_214,dangling_wire_215,dangling_wire_216,N__33071,dangling_wire_217,dangling_wire_218,dangling_wire_219}),
            .RCLKE(),
            .RCLK(N__34419),
            .RE(N__37256),
            .WCLKE(N__21469),
            .WCLK(N__34418),
            .WE(N__37199));
    defparam \b2v_inst8.mem_mem_0_1_physical .WRITE_MODE=3;
    defparam \b2v_inst8.mem_mem_0_1_physical .READ_MODE=3;
    SB_RAM40_4K \b2v_inst8.mem_mem_0_1_physical  (
            .RDATA({dangling_wire_220,dangling_wire_221,dangling_wire_222,dangling_wire_223,SYNTHESIZED_WIRE_1_3,dangling_wire_224,dangling_wire_225,dangling_wire_226,dangling_wire_227,dangling_wire_228,dangling_wire_229,dangling_wire_230,SYNTHESIZED_WIRE_1_2,dangling_wire_231,dangling_wire_232,dangling_wire_233}),
            .RADDR({N__36613,N__35758,N__38959,N__38746,N__38188,N__35536,N__36196,N__36409,N__35986,N__38500,N__39178}),
            .WADDR({N__36622,N__35761,N__38956,N__38743,N__38185,N__35539,N__36199,N__36412,N__35989,N__38497,N__39175}),
            .MASK({dangling_wire_234,dangling_wire_235,dangling_wire_236,dangling_wire_237,dangling_wire_238,dangling_wire_239,dangling_wire_240,dangling_wire_241,dangling_wire_242,dangling_wire_243,dangling_wire_244,dangling_wire_245,dangling_wire_246,dangling_wire_247,dangling_wire_248,dangling_wire_249}),
            .WDATA({dangling_wire_250,dangling_wire_251,dangling_wire_252,dangling_wire_253,N__33197,dangling_wire_254,dangling_wire_255,dangling_wire_256,dangling_wire_257,dangling_wire_258,dangling_wire_259,dangling_wire_260,N__32558,dangling_wire_261,dangling_wire_262,dangling_wire_263}),
            .RCLKE(),
            .RCLK(N__34389),
            .RE(N__36836),
            .WCLKE(N__21454),
            .WCLK(N__34390),
            .WE(N__36837));
    defparam \b2v_inst7.mem_mem_0_4_physical .WRITE_MODE=3;
    defparam \b2v_inst7.mem_mem_0_4_physical .READ_MODE=3;
    SB_RAM40_4K \b2v_inst7.mem_mem_0_4_physical  (
            .RDATA({dangling_wire_264,dangling_wire_265,dangling_wire_266,dangling_wire_267,leds_c_9,dangling_wire_268,dangling_wire_269,dangling_wire_270,dangling_wire_271,dangling_wire_272,dangling_wire_273,dangling_wire_274,leds_c_8,dangling_wire_275,dangling_wire_276,dangling_wire_277}),
            .RADDR({N__20104,N__15931,N__14125,N__14308,N__18679,N__19855,N__21550,N__20488,N__19972,N__14404,N__14215}),
            .WADDR({N__20101,N__15928,N__14122,N__14317,N__18676,N__19852,N__21547,N__20485,N__19969,N__14407,N__14218}),
            .MASK({dangling_wire_278,dangling_wire_279,dangling_wire_280,dangling_wire_281,dangling_wire_282,dangling_wire_283,dangling_wire_284,dangling_wire_285,dangling_wire_286,dangling_wire_287,dangling_wire_288,dangling_wire_289,dangling_wire_290,dangling_wire_291,dangling_wire_292,dangling_wire_293}),
            .WDATA({dangling_wire_294,dangling_wire_295,dangling_wire_296,dangling_wire_297,N__16949,dangling_wire_298,dangling_wire_299,dangling_wire_300,dangling_wire_301,dangling_wire_302,dangling_wire_303,dangling_wire_304,N__16940,dangling_wire_305,dangling_wire_306,dangling_wire_307}),
            .RCLKE(),
            .RCLK(N__34520),
            .RE(N__37213),
            .WCLKE(N__21448),
            .WCLK(N__34521),
            .WE(N__37226));
    defparam \b2v_inst7.mem_mem_0_1_physical .WRITE_MODE=3;
    defparam \b2v_inst7.mem_mem_0_1_physical .READ_MODE=3;
    SB_RAM40_4K \b2v_inst7.mem_mem_0_1_physical  (
            .RDATA({dangling_wire_308,dangling_wire_309,dangling_wire_310,dangling_wire_311,leds_c_3,dangling_wire_312,dangling_wire_313,dangling_wire_314,dangling_wire_315,dangling_wire_316,dangling_wire_317,dangling_wire_318,leds_c_2,dangling_wire_319,dangling_wire_320,dangling_wire_321}),
            .RADDR({N__20140,N__15967,N__14161,N__14344,N__18715,N__19891,N__21586,N__20524,N__20008,N__14440,N__14251}),
            .WADDR({N__20137,N__15964,N__14158,N__14353,N__18712,N__19888,N__21583,N__20521,N__20005,N__14443,N__14254}),
            .MASK({dangling_wire_322,dangling_wire_323,dangling_wire_324,dangling_wire_325,dangling_wire_326,dangling_wire_327,dangling_wire_328,dangling_wire_329,dangling_wire_330,dangling_wire_331,dangling_wire_332,dangling_wire_333,dangling_wire_334,dangling_wire_335,dangling_wire_336,dangling_wire_337}),
            .WDATA({dangling_wire_338,dangling_wire_339,dangling_wire_340,dangling_wire_341,N__21917,dangling_wire_342,dangling_wire_343,dangling_wire_344,dangling_wire_345,dangling_wire_346,dangling_wire_347,dangling_wire_348,N__21206,dangling_wire_349,dangling_wire_350,dangling_wire_351}),
            .RCLKE(),
            .RCLK(N__34504),
            .RE(N__37286),
            .WCLKE(N__21391),
            .WCLK(N__34505),
            .WE(N__37249));
    defparam \b2v_inst2.mem_mem_0_4_physical .WRITE_MODE=3;
    defparam \b2v_inst2.mem_mem_0_4_physical .READ_MODE=3;
    SB_RAM40_4K \b2v_inst2.mem_mem_0_4_physical  (
            .RDATA({dangling_wire_352,dangling_wire_353,dangling_wire_354,dangling_wire_355,SYNTHESIZED_WIRE_3_9,dangling_wire_356,dangling_wire_357,dangling_wire_358,dangling_wire_359,dangling_wire_360,dangling_wire_361,dangling_wire_362,SYNTHESIZED_WIRE_3_8,dangling_wire_363,dangling_wire_364,dangling_wire_365}),
            .RADDR({N__33430,N__33730,N__33844,N__19426,N__32737,N__33961,N__18421,N__19603,N__35011,N__35362,N__33544}),
            .WADDR({N__33427,N__33733,N__33847,N__19423,N__32740,N__33964,N__18430,N__19618,N__35008,N__35365,N__33541}),
            .MASK({dangling_wire_366,dangling_wire_367,dangling_wire_368,dangling_wire_369,dangling_wire_370,dangling_wire_371,dangling_wire_372,dangling_wire_373,dangling_wire_374,dangling_wire_375,dangling_wire_376,dangling_wire_377,dangling_wire_378,dangling_wire_379,dangling_wire_380,dangling_wire_381}),
            .WDATA({dangling_wire_382,dangling_wire_383,dangling_wire_384,dangling_wire_385,N__32825,dangling_wire_386,dangling_wire_387,dangling_wire_388,dangling_wire_389,dangling_wire_390,dangling_wire_391,dangling_wire_392,N__33356,dangling_wire_393,dangling_wire_394,dangling_wire_395}),
            .RCLKE(),
            .RCLK(N__34374),
            .RE(N__37014),
            .WCLKE(N__21456),
            .WCLK(N__34375),
            .WE(N__37015));
    defparam \b2v_inst2.mem_mem_0_3_physical .WRITE_MODE=3;
    defparam \b2v_inst2.mem_mem_0_3_physical .READ_MODE=3;
    SB_RAM40_4K \b2v_inst2.mem_mem_0_3_physical  (
            .RDATA({dangling_wire_396,dangling_wire_397,dangling_wire_398,dangling_wire_399,SYNTHESIZED_WIRE_3_7,dangling_wire_400,dangling_wire_401,dangling_wire_402,dangling_wire_403,dangling_wire_404,dangling_wire_405,dangling_wire_406,SYNTHESIZED_WIRE_3_6,dangling_wire_407,dangling_wire_408,dangling_wire_409}),
            .RADDR({N__33442,N__33742,N__33856,N__19438,N__32749,N__33973,N__18433,N__19615,N__35023,N__35374,N__33556}),
            .WADDR({N__33439,N__33745,N__33859,N__19435,N__32752,N__33976,N__18442,N__19630,N__35020,N__35377,N__33553}),
            .MASK({dangling_wire_410,dangling_wire_411,dangling_wire_412,dangling_wire_413,dangling_wire_414,dangling_wire_415,dangling_wire_416,dangling_wire_417,dangling_wire_418,dangling_wire_419,dangling_wire_420,dangling_wire_421,dangling_wire_422,dangling_wire_423,dangling_wire_424,dangling_wire_425}),
            .WDATA({dangling_wire_426,dangling_wire_427,dangling_wire_428,dangling_wire_429,N__35462,dangling_wire_430,dangling_wire_431,dangling_wire_432,dangling_wire_433,dangling_wire_434,dangling_wire_435,dangling_wire_436,N__35270,dangling_wire_437,dangling_wire_438,dangling_wire_439}),
            .RCLKE(),
            .RCLK(N__34387),
            .RE(N__37112),
            .WCLKE(N__21457),
            .WCLK(N__34388),
            .WE(N__37029));
    defparam \b2v_inst7.mem_mem_0_6_physical .WRITE_MODE=3;
    defparam \b2v_inst7.mem_mem_0_6_physical .READ_MODE=3;
    SB_RAM40_4K \b2v_inst7.mem_mem_0_6_physical  (
            .RDATA({dangling_wire_440,dangling_wire_441,dangling_wire_442,dangling_wire_443,leds_c_13,dangling_wire_444,dangling_wire_445,dangling_wire_446,dangling_wire_447,dangling_wire_448,dangling_wire_449,dangling_wire_450,leds_c_12,dangling_wire_451,dangling_wire_452,dangling_wire_453}),
            .RADDR({N__20080,N__15907,N__14101,N__14284,N__18655,N__19831,N__21526,N__20464,N__19948,N__14380,N__14191}),
            .WADDR({N__20077,N__15904,N__14098,N__14293,N__18652,N__19828,N__21523,N__20461,N__19945,N__14383,N__14194}),
            .MASK({dangling_wire_454,dangling_wire_455,dangling_wire_456,dangling_wire_457,dangling_wire_458,dangling_wire_459,dangling_wire_460,dangling_wire_461,dangling_wire_462,dangling_wire_463,dangling_wire_464,dangling_wire_465,dangling_wire_466,dangling_wire_467,dangling_wire_468,dangling_wire_469}),
            .WDATA({dangling_wire_470,dangling_wire_471,dangling_wire_472,dangling_wire_473,N__24992,dangling_wire_474,dangling_wire_475,dangling_wire_476,dangling_wire_477,dangling_wire_478,dangling_wire_479,dangling_wire_480,N__25034,dangling_wire_481,dangling_wire_482,dangling_wire_483}),
            .RCLKE(),
            .RCLK(N__34528),
            .RE(N__37282),
            .WCLKE(N__21467),
            .WCLK(N__34529),
            .WE(N__37285));
    defparam \b2v_inst8.mem_mem_0_2_physical .WRITE_MODE=3;
    defparam \b2v_inst8.mem_mem_0_2_physical .READ_MODE=3;
    SB_RAM40_4K \b2v_inst8.mem_mem_0_2_physical  (
            .RDATA({dangling_wire_484,dangling_wire_485,dangling_wire_486,dangling_wire_487,SYNTHESIZED_WIRE_1_5,dangling_wire_488,dangling_wire_489,dangling_wire_490,dangling_wire_491,dangling_wire_492,dangling_wire_493,dangling_wire_494,SYNTHESIZED_WIRE_1_4,dangling_wire_495,dangling_wire_496,dangling_wire_497}),
            .RADDR({N__36601,N__35746,N__38947,N__38734,N__38176,N__35524,N__36184,N__36397,N__35974,N__38488,N__39166}),
            .WADDR({N__36610,N__35749,N__38944,N__38731,N__38173,N__35527,N__36187,N__36400,N__35977,N__38485,N__39163}),
            .MASK({dangling_wire_498,dangling_wire_499,dangling_wire_500,dangling_wire_501,dangling_wire_502,dangling_wire_503,dangling_wire_504,dangling_wire_505,dangling_wire_506,dangling_wire_507,dangling_wire_508,dangling_wire_509,dangling_wire_510,dangling_wire_511,dangling_wire_512,dangling_wire_513}),
            .WDATA({dangling_wire_514,dangling_wire_515,dangling_wire_516,dangling_wire_517,N__37316,dangling_wire_518,dangling_wire_519,dangling_wire_520,dangling_wire_521,dangling_wire_522,dangling_wire_523,dangling_wire_524,N__33275,dangling_wire_525,dangling_wire_526,dangling_wire_527}),
            .RCLKE(),
            .RCLK(N__34402),
            .RE(N__36921),
            .WCLKE(N__21455),
            .WCLK(N__34403),
            .WE(N__37012));
    defparam \b2v_inst7.mem_mem_0_3_physical .WRITE_MODE=3;
    defparam \b2v_inst7.mem_mem_0_3_physical .READ_MODE=3;
    SB_RAM40_4K \b2v_inst7.mem_mem_0_3_physical  (
            .RDATA({dangling_wire_528,dangling_wire_529,dangling_wire_530,dangling_wire_531,leds_c_7,dangling_wire_532,dangling_wire_533,dangling_wire_534,dangling_wire_535,dangling_wire_536,dangling_wire_537,dangling_wire_538,leds_c_6,dangling_wire_539,dangling_wire_540,dangling_wire_541}),
            .RADDR({N__20116,N__15943,N__14137,N__14320,N__18691,N__19867,N__21562,N__20500,N__19984,N__14416,N__14227}),
            .WADDR({N__20113,N__15940,N__14134,N__14329,N__18688,N__19864,N__21559,N__20497,N__19981,N__14419,N__14230}),
            .MASK({dangling_wire_542,dangling_wire_543,dangling_wire_544,dangling_wire_545,dangling_wire_546,dangling_wire_547,dangling_wire_548,dangling_wire_549,dangling_wire_550,dangling_wire_551,dangling_wire_552,dangling_wire_553,dangling_wire_554,dangling_wire_555,dangling_wire_556,dangling_wire_557}),
            .WDATA({dangling_wire_558,dangling_wire_559,dangling_wire_560,dangling_wire_561,N__23477,dangling_wire_562,dangling_wire_563,dangling_wire_564,dangling_wire_565,dangling_wire_566,dangling_wire_567,dangling_wire_568,N__15443,dangling_wire_569,dangling_wire_570,dangling_wire_571}),
            .RCLKE(),
            .RCLK(N__34506),
            .RE(N__37160),
            .WCLKE(N__21410),
            .WCLK(N__34507),
            .WE(N__37235));
    defparam \b2v_inst7.mem_mem_0_0_physical .WRITE_MODE=3;
    defparam \b2v_inst7.mem_mem_0_0_physical .READ_MODE=3;
    SB_RAM40_4K \b2v_inst7.mem_mem_0_0_physical  (
            .RDATA({dangling_wire_572,dangling_wire_573,dangling_wire_574,dangling_wire_575,leds_c_1,dangling_wire_576,dangling_wire_577,dangling_wire_578,dangling_wire_579,dangling_wire_580,dangling_wire_581,dangling_wire_582,leds_c_0,dangling_wire_583,dangling_wire_584,dangling_wire_585}),
            .RADDR({N__20150,N__15977,N__14171,N__14356,N__18725,N__19901,N__21596,N__20534,N__20018,N__14452,N__14263}),
            .WADDR({N__20149,N__15976,N__14170,N__14360,N__18724,N__19900,N__21595,N__20533,N__20017,N__14453,N__14264}),
            .MASK({dangling_wire_586,dangling_wire_587,dangling_wire_588,dangling_wire_589,dangling_wire_590,dangling_wire_591,dangling_wire_592,dangling_wire_593,dangling_wire_594,dangling_wire_595,dangling_wire_596,dangling_wire_597,dangling_wire_598,dangling_wire_599,dangling_wire_600,dangling_wire_601}),
            .WDATA({dangling_wire_602,dangling_wire_603,dangling_wire_604,dangling_wire_605,N__20858,dangling_wire_606,dangling_wire_607,dangling_wire_608,dangling_wire_609,dangling_wire_610,dangling_wire_611,dangling_wire_612,N__20576,dangling_wire_613,dangling_wire_614,dangling_wire_615}),
            .RCLKE(),
            .RCLK(N__34518),
            .RE(N__37287),
            .WCLKE(N__21426),
            .WCLK(N__34519),
            .WE(N__37283));
    defparam \b2v_inst2.mem_mem_0_5_physical .WRITE_MODE=3;
    defparam \b2v_inst2.mem_mem_0_5_physical .READ_MODE=3;
    SB_RAM40_4K \b2v_inst2.mem_mem_0_5_physical  (
            .RDATA({dangling_wire_616,dangling_wire_617,dangling_wire_618,dangling_wire_619,dangling_wire_620,dangling_wire_621,dangling_wire_622,dangling_wire_623,dangling_wire_624,dangling_wire_625,dangling_wire_626,dangling_wire_627,SYNTHESIZED_WIRE_3_10,dangling_wire_628,dangling_wire_629,dangling_wire_630}),
            .RADDR({N__33418,N__33718,N__33832,N__19414,N__32725,N__33949,N__18409,N__19591,N__34999,N__35350,N__33532}),
            .WADDR({N__33415,N__33721,N__33835,N__19411,N__32728,N__33952,N__18418,N__19606,N__34996,N__35353,N__33529}),
            .MASK({dangling_wire_631,dangling_wire_632,dangling_wire_633,dangling_wire_634,dangling_wire_635,dangling_wire_636,dangling_wire_637,dangling_wire_638,dangling_wire_639,dangling_wire_640,dangling_wire_641,dangling_wire_642,dangling_wire_643,dangling_wire_644,dangling_wire_645,dangling_wire_646}),
            .WDATA({dangling_wire_647,dangling_wire_648,dangling_wire_649,dangling_wire_650,dangling_wire_651,dangling_wire_652,dangling_wire_653,dangling_wire_654,dangling_wire_655,dangling_wire_656,dangling_wire_657,dangling_wire_658,N__33632,dangling_wire_659,dangling_wire_660,dangling_wire_661}),
            .RCLKE(),
            .RCLK(N__34371),
            .RE(N__37013),
            .WCLKE(N__21427),
            .WCLK(N__34372),
            .WE(N__36938));
    defparam \b2v_inst7.mem_mem_0_5_physical .WRITE_MODE=3;
    defparam \b2v_inst7.mem_mem_0_5_physical .READ_MODE=3;
    SB_RAM40_4K \b2v_inst7.mem_mem_0_5_physical  (
            .RDATA({dangling_wire_662,dangling_wire_663,dangling_wire_664,dangling_wire_665,leds_c_11,dangling_wire_666,dangling_wire_667,dangling_wire_668,dangling_wire_669,dangling_wire_670,dangling_wire_671,dangling_wire_672,leds_c_10,dangling_wire_673,dangling_wire_674,dangling_wire_675}),
            .RADDR({N__20092,N__15919,N__14113,N__14296,N__18667,N__19843,N__21538,N__20476,N__19960,N__14392,N__14203}),
            .WADDR({N__20089,N__15916,N__14110,N__14305,N__18664,N__19840,N__21535,N__20473,N__19957,N__14395,N__14206}),
            .MASK({dangling_wire_676,dangling_wire_677,dangling_wire_678,dangling_wire_679,dangling_wire_680,dangling_wire_681,dangling_wire_682,dangling_wire_683,dangling_wire_684,dangling_wire_685,dangling_wire_686,dangling_wire_687,dangling_wire_688,dangling_wire_689,dangling_wire_690,dangling_wire_691}),
            .WDATA({dangling_wire_692,dangling_wire_693,dangling_wire_694,dangling_wire_695,N__25082,dangling_wire_696,dangling_wire_697,dangling_wire_698,dangling_wire_699,dangling_wire_700,dangling_wire_701,dangling_wire_702,N__24926,dangling_wire_703,dangling_wire_704,dangling_wire_705}),
            .RCLKE(),
            .RCLK(N__34526),
            .RE(N__37227),
            .WCLKE(N__21449),
            .WCLK(N__34527),
            .WE(N__37284));
    PRE_IO_GBUF clk_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__39654),
            .GLOBALBUFFEROUTPUT(clk_c_g));
    IO_PAD clk_ibuf_gb_io_iopad (
            .OE(N__39656),
            .DIN(N__39655),
            .DOUT(N__39654),
            .PACKAGEPIN(clk));
    defparam clk_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam clk_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO clk_ibuf_gb_io_preio (
            .PADOEN(N__39656),
            .PADOUT(N__39655),
            .PADIN(N__39654),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD leds_obuf_9_iopad (
            .OE(N__39645),
            .DIN(N__39644),
            .DOUT(N__39643),
            .PACKAGEPIN(leds[9]));
    defparam leds_obuf_9_preio.NEG_TRIGGER=1'b0;
    defparam leds_obuf_9_preio.PIN_TYPE=6'b011001;
    PRE_IO leds_obuf_9_preio (
            .PADOEN(N__39645),
            .PADOUT(N__39644),
            .PADIN(N__39643),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__26261),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD swit_ibuf_0_iopad (
            .OE(N__39636),
            .DIN(N__39635),
            .DOUT(N__39634),
            .PACKAGEPIN(swit[0]));
    defparam swit_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam swit_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO swit_ibuf_0_preio (
            .PADOEN(N__39636),
            .PADOUT(N__39635),
            .PADIN(N__39634),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(swit_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD leds_obuf_3_iopad (
            .OE(N__39627),
            .DIN(N__39626),
            .DOUT(N__39625),
            .PACKAGEPIN(leds[3]));
    defparam leds_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam leds_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO leds_obuf_3_preio (
            .PADOEN(N__39627),
            .PADOUT(N__39626),
            .PADIN(N__39625),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__23653),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD swit_ibuf_6_iopad (
            .OE(N__39618),
            .DIN(N__39617),
            .DOUT(N__39616),
            .PACKAGEPIN(swit[6]));
    defparam swit_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam swit_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO swit_ibuf_6_preio (
            .PADOEN(N__39618),
            .PADOUT(N__39617),
            .PADIN(N__39616),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(swit_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD leds_obuf_5_iopad (
            .OE(N__39609),
            .DIN(N__39608),
            .DOUT(N__39607),
            .PACKAGEPIN(leds[5]));
    defparam leds_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam leds_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO leds_obuf_5_preio (
            .PADOEN(N__39609),
            .PADOUT(N__39608),
            .PADIN(N__39607),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__17156),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD swit_ibuf_8_iopad (
            .OE(N__39600),
            .DIN(N__39599),
            .DOUT(N__39598),
            .PACKAGEPIN(swit[8]));
    defparam swit_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam swit_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO swit_ibuf_8_preio (
            .PADOEN(N__39600),
            .PADOUT(N__39599),
            .PADIN(N__39598),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(swit_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD swit_ibuf_3_iopad (
            .OE(N__39591),
            .DIN(N__39590),
            .DOUT(N__39589),
            .PACKAGEPIN(swit[3]));
    defparam swit_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam swit_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO swit_ibuf_3_preio (
            .PADOEN(N__39591),
            .PADOUT(N__39590),
            .PADIN(N__39589),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(swit_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD leds_obuf_0_iopad (
            .OE(N__39582),
            .DIN(N__39581),
            .DOUT(N__39580),
            .PACKAGEPIN(leds[0]));
    defparam leds_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam leds_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO leds_obuf_0_preio (
            .PADOEN(N__39582),
            .PADOUT(N__39581),
            .PADIN(N__39580),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__23404),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD leds_obuf_11_iopad (
            .OE(N__39573),
            .DIN(N__39572),
            .DOUT(N__39571),
            .PACKAGEPIN(leds[11]));
    defparam leds_obuf_11_preio.NEG_TRIGGER=1'b0;
    defparam leds_obuf_11_preio.PIN_TYPE=6'b011001;
    PRE_IO leds_obuf_11_preio (
            .PADOEN(N__39573),
            .PADOUT(N__39572),
            .PADIN(N__39571),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__17795),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD swit_ibuf_4_iopad (
            .OE(N__39564),
            .DIN(N__39563),
            .DOUT(N__39562),
            .PACKAGEPIN(swit[4]));
    defparam swit_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam swit_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO swit_ibuf_4_preio (
            .PADOEN(N__39564),
            .PADOUT(N__39563),
            .PADIN(N__39562),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(swit_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD leds_obuf_7_iopad (
            .OE(N__39555),
            .DIN(N__39554),
            .DOUT(N__39553),
            .PACKAGEPIN(leds[7]));
    defparam leds_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam leds_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO leds_obuf_7_preio (
            .PADOEN(N__39555),
            .PADOUT(N__39554),
            .PADIN(N__39553),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__17764),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD swit_ibuf_10_iopad (
            .OE(N__39546),
            .DIN(N__39545),
            .DOUT(N__39544),
            .PACKAGEPIN(swit[10]));
    defparam swit_ibuf_10_preio.NEG_TRIGGER=1'b0;
    defparam swit_ibuf_10_preio.PIN_TYPE=6'b000001;
    PRE_IO swit_ibuf_10_preio (
            .PADOEN(N__39546),
            .PADOUT(N__39545),
            .PADIN(N__39544),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(swit_c_10),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD uart_rx_i_ibuf_iopad (
            .OE(N__39537),
            .DIN(N__39536),
            .DOUT(N__39535),
            .PACKAGEPIN(uart_rx_i));
    defparam uart_rx_i_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam uart_rx_i_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO uart_rx_i_ibuf_preio (
            .PADOEN(N__39537),
            .PADOUT(N__39536),
            .PADIN(N__39535),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(uart_rx_i_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD leds_obuf_8_iopad (
            .OE(N__39528),
            .DIN(N__39527),
            .DOUT(N__39526),
            .PACKAGEPIN(leds[8]));
    defparam leds_obuf_8_preio.NEG_TRIGGER=1'b0;
    defparam leds_obuf_8_preio.PIN_TYPE=6'b011001;
    PRE_IO leds_obuf_8_preio (
            .PADOEN(N__39528),
            .PADOUT(N__39527),
            .PADIN(N__39526),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__24977),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD reset_ibuf_iopad (
            .OE(N__39519),
            .DIN(N__39518),
            .DOUT(N__39517),
            .PACKAGEPIN(reset));
    defparam reset_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam reset_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO reset_ibuf_preio (
            .PADOEN(N__39519),
            .PADOUT(N__39518),
            .PADIN(N__39517),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(reset_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD swit_ibuf_1_iopad (
            .OE(N__39510),
            .DIN(N__39509),
            .DOUT(N__39508),
            .PACKAGEPIN(swit[1]));
    defparam swit_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam swit_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO swit_ibuf_1_preio (
            .PADOEN(N__39510),
            .PADOUT(N__39509),
            .PADIN(N__39508),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(swit_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD leds_obuf_2_iopad (
            .OE(N__39501),
            .DIN(N__39500),
            .DOUT(N__39499),
            .PACKAGEPIN(leds[2]));
    defparam leds_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam leds_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO leds_obuf_2_preio (
            .PADOEN(N__39501),
            .PADOUT(N__39500),
            .PADIN(N__39499),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__23674),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD leds_obuf_13_iopad (
            .OE(N__39492),
            .DIN(N__39491),
            .DOUT(N__39490),
            .PACKAGEPIN(leds[13]));
    defparam leds_obuf_13_preio.NEG_TRIGGER=1'b0;
    defparam leds_obuf_13_preio.PIN_TYPE=6'b011001;
    PRE_IO leds_obuf_13_preio (
            .PADOEN(N__39492),
            .PADOUT(N__39491),
            .PADIN(N__39490),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__23332),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD swit_ibuf_2_iopad (
            .OE(N__39483),
            .DIN(N__39482),
            .DOUT(N__39481),
            .PACKAGEPIN(swit[2]));
    defparam swit_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam swit_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO swit_ibuf_2_preio (
            .PADOEN(N__39483),
            .PADOUT(N__39482),
            .PADIN(N__39481),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(swit_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD leds_obuf_1_iopad (
            .OE(N__39474),
            .DIN(N__39473),
            .DOUT(N__39472),
            .PACKAGEPIN(leds[1]));
    defparam leds_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam leds_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO leds_obuf_1_preio (
            .PADOEN(N__39474),
            .PADOUT(N__39473),
            .PADIN(N__39472),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__23372),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD leds_obuf_10_iopad (
            .OE(N__39465),
            .DIN(N__39464),
            .DOUT(N__39463),
            .PACKAGEPIN(leds[10]));
    defparam leds_obuf_10_preio.NEG_TRIGGER=1'b0;
    defparam leds_obuf_10_preio.PIN_TYPE=6'b011001;
    PRE_IO leds_obuf_10_preio (
            .PADOEN(N__39465),
            .PADOUT(N__39464),
            .PADIN(N__39463),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__17825),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD swit_ibuf_7_iopad (
            .OE(N__39456),
            .DIN(N__39455),
            .DOUT(N__39454),
            .PACKAGEPIN(swit[7]));
    defparam swit_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam swit_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO swit_ibuf_7_preio (
            .PADOEN(N__39456),
            .PADOUT(N__39455),
            .PADIN(N__39454),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(swit_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD leds_obuf_4_iopad (
            .OE(N__39447),
            .DIN(N__39446),
            .DOUT(N__39445),
            .PACKAGEPIN(leds[4]));
    defparam leds_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam leds_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO leds_obuf_4_preio (
            .PADOEN(N__39447),
            .PADOUT(N__39446),
            .PADIN(N__39445),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__17192),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD swit_ibuf_9_iopad (
            .OE(N__39438),
            .DIN(N__39437),
            .DOUT(N__39436),
            .PACKAGEPIN(swit[9]));
    defparam swit_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam swit_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO swit_ibuf_9_preio (
            .PADOEN(N__39438),
            .PADOUT(N__39437),
            .PADIN(N__39436),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(swit_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD uart_tx_o_obuf_iopad (
            .OE(N__39429),
            .DIN(N__39428),
            .DOUT(N__39427),
            .PACKAGEPIN(uart_tx_o));
    defparam uart_tx_o_obuf_preio.NEG_TRIGGER=1'b0;
    defparam uart_tx_o_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO uart_tx_o_obuf_preio (
            .PADOEN(N__39429),
            .PADOUT(N__39428),
            .PADIN(N__39427),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__26099),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD leds_obuf_12_iopad (
            .OE(N__39420),
            .DIN(N__39419),
            .DOUT(N__39418),
            .PACKAGEPIN(leds[12]));
    defparam leds_obuf_12_preio.NEG_TRIGGER=1'b0;
    defparam leds_obuf_12_preio.PIN_TYPE=6'b011001;
    PRE_IO leds_obuf_12_preio (
            .PADOEN(N__39420),
            .PADOUT(N__39419),
            .PADIN(N__39418),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__18875),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD swit_ibuf_5_iopad (
            .OE(N__39411),
            .DIN(N__39410),
            .DOUT(N__39409),
            .PACKAGEPIN(swit[5]));
    defparam swit_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam swit_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO swit_ibuf_5_preio (
            .PADOEN(N__39411),
            .PADOUT(N__39410),
            .PADIN(N__39409),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(swit_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD leds_obuf_6_iopad (
            .OE(N__39402),
            .DIN(N__39401),
            .DOUT(N__39400),
            .PACKAGEPIN(leds[6]));
    defparam leds_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam leds_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO leds_obuf_6_preio (
            .PADOEN(N__39402),
            .PADOUT(N__39401),
            .PADIN(N__39400),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__20432),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    CascadeMux I__9791 (
            .O(N__39383),
            .I(N__39380));
    InMux I__9790 (
            .O(N__39380),
            .I(N__39377));
    LocalMux I__9789 (
            .O(N__39377),
            .I(N__39373));
    InMux I__9788 (
            .O(N__39376),
            .I(N__39370));
    Span4Mux_v I__9787 (
            .O(N__39373),
            .I(N__39366));
    LocalMux I__9786 (
            .O(N__39370),
            .I(N__39363));
    InMux I__9785 (
            .O(N__39369),
            .I(N__39360));
    Span4Mux_h I__9784 (
            .O(N__39366),
            .I(N__39356));
    Span4Mux_h I__9783 (
            .O(N__39363),
            .I(N__39351));
    LocalMux I__9782 (
            .O(N__39360),
            .I(N__39351));
    InMux I__9781 (
            .O(N__39359),
            .I(N__39346));
    Span4Mux_h I__9780 (
            .O(N__39356),
            .I(N__39343));
    Span4Mux_v I__9779 (
            .O(N__39351),
            .I(N__39340));
    InMux I__9778 (
            .O(N__39350),
            .I(N__39337));
    InMux I__9777 (
            .O(N__39349),
            .I(N__39334));
    LocalMux I__9776 (
            .O(N__39346),
            .I(\b2v_inst.dir_energiaZ0Z_0 ));
    Odrv4 I__9775 (
            .O(N__39343),
            .I(\b2v_inst.dir_energiaZ0Z_0 ));
    Odrv4 I__9774 (
            .O(N__39340),
            .I(\b2v_inst.dir_energiaZ0Z_0 ));
    LocalMux I__9773 (
            .O(N__39337),
            .I(\b2v_inst.dir_energiaZ0Z_0 ));
    LocalMux I__9772 (
            .O(N__39334),
            .I(\b2v_inst.dir_energiaZ0Z_0 ));
    InMux I__9771 (
            .O(N__39323),
            .I(N__39319));
    InMux I__9770 (
            .O(N__39322),
            .I(N__39313));
    LocalMux I__9769 (
            .O(N__39319),
            .I(N__39310));
    InMux I__9768 (
            .O(N__39318),
            .I(N__39307));
    InMux I__9767 (
            .O(N__39317),
            .I(N__39300));
    CascadeMux I__9766 (
            .O(N__39316),
            .I(N__39297));
    LocalMux I__9765 (
            .O(N__39313),
            .I(N__39294));
    Span4Mux_v I__9764 (
            .O(N__39310),
            .I(N__39289));
    LocalMux I__9763 (
            .O(N__39307),
            .I(N__39289));
    InMux I__9762 (
            .O(N__39306),
            .I(N__39286));
    InMux I__9761 (
            .O(N__39305),
            .I(N__39283));
    InMux I__9760 (
            .O(N__39304),
            .I(N__39280));
    InMux I__9759 (
            .O(N__39303),
            .I(N__39277));
    LocalMux I__9758 (
            .O(N__39300),
            .I(N__39274));
    InMux I__9757 (
            .O(N__39297),
            .I(N__39270));
    Span4Mux_v I__9756 (
            .O(N__39294),
            .I(N__39267));
    Span4Mux_v I__9755 (
            .O(N__39289),
            .I(N__39264));
    LocalMux I__9754 (
            .O(N__39286),
            .I(N__39261));
    LocalMux I__9753 (
            .O(N__39283),
            .I(N__39258));
    LocalMux I__9752 (
            .O(N__39280),
            .I(N__39255));
    LocalMux I__9751 (
            .O(N__39277),
            .I(N__39252));
    Span4Mux_h I__9750 (
            .O(N__39274),
            .I(N__39249));
    InMux I__9749 (
            .O(N__39273),
            .I(N__39246));
    LocalMux I__9748 (
            .O(N__39270),
            .I(N__39243));
    Span4Mux_h I__9747 (
            .O(N__39267),
            .I(N__39237));
    Span4Mux_h I__9746 (
            .O(N__39264),
            .I(N__39237));
    Span4Mux_v I__9745 (
            .O(N__39261),
            .I(N__39228));
    Span4Mux_v I__9744 (
            .O(N__39258),
            .I(N__39228));
    Span4Mux_h I__9743 (
            .O(N__39255),
            .I(N__39228));
    Span4Mux_v I__9742 (
            .O(N__39252),
            .I(N__39228));
    Sp12to4 I__9741 (
            .O(N__39249),
            .I(N__39223));
    LocalMux I__9740 (
            .O(N__39246),
            .I(N__39220));
    Span4Mux_h I__9739 (
            .O(N__39243),
            .I(N__39217));
    InMux I__9738 (
            .O(N__39242),
            .I(N__39214));
    Span4Mux_v I__9737 (
            .O(N__39237),
            .I(N__39209));
    Span4Mux_h I__9736 (
            .O(N__39228),
            .I(N__39209));
    InMux I__9735 (
            .O(N__39227),
            .I(N__39204));
    InMux I__9734 (
            .O(N__39226),
            .I(N__39204));
    Span12Mux_v I__9733 (
            .O(N__39223),
            .I(N__39199));
    Span12Mux_h I__9732 (
            .O(N__39220),
            .I(N__39199));
    Odrv4 I__9731 (
            .O(N__39217),
            .I(\b2v_inst.indiceZ0Z_0 ));
    LocalMux I__9730 (
            .O(N__39214),
            .I(\b2v_inst.indiceZ0Z_0 ));
    Odrv4 I__9729 (
            .O(N__39209),
            .I(\b2v_inst.indiceZ0Z_0 ));
    LocalMux I__9728 (
            .O(N__39204),
            .I(\b2v_inst.indiceZ0Z_0 ));
    Odrv12 I__9727 (
            .O(N__39199),
            .I(\b2v_inst.indiceZ0Z_0 ));
    CascadeMux I__9726 (
            .O(N__39188),
            .I(N__39184));
    CascadeMux I__9725 (
            .O(N__39187),
            .I(N__39181));
    CascadeBuf I__9724 (
            .O(N__39184),
            .I(N__39178));
    CascadeBuf I__9723 (
            .O(N__39181),
            .I(N__39175));
    CascadeMux I__9722 (
            .O(N__39178),
            .I(N__39172));
    CascadeMux I__9721 (
            .O(N__39175),
            .I(N__39169));
    CascadeBuf I__9720 (
            .O(N__39172),
            .I(N__39166));
    CascadeBuf I__9719 (
            .O(N__39169),
            .I(N__39163));
    CascadeMux I__9718 (
            .O(N__39166),
            .I(N__39160));
    CascadeMux I__9717 (
            .O(N__39163),
            .I(N__39157));
    InMux I__9716 (
            .O(N__39160),
            .I(N__39154));
    InMux I__9715 (
            .O(N__39157),
            .I(N__39151));
    LocalMux I__9714 (
            .O(N__39154),
            .I(N_360_i));
    LocalMux I__9713 (
            .O(N__39151),
            .I(N_360_i));
    InMux I__9712 (
            .O(N__39146),
            .I(N__39143));
    LocalMux I__9711 (
            .O(N__39143),
            .I(N__39140));
    Span4Mux_h I__9710 (
            .O(N__39140),
            .I(N__39135));
    InMux I__9709 (
            .O(N__39139),
            .I(N__39132));
    InMux I__9708 (
            .O(N__39138),
            .I(N__39129));
    Span4Mux_h I__9707 (
            .O(N__39135),
            .I(N__39124));
    LocalMux I__9706 (
            .O(N__39132),
            .I(N__39124));
    LocalMux I__9705 (
            .O(N__39129),
            .I(N__39119));
    Span4Mux_h I__9704 (
            .O(N__39124),
            .I(N__39116));
    InMux I__9703 (
            .O(N__39123),
            .I(N__39113));
    InMux I__9702 (
            .O(N__39122),
            .I(N__39110));
    Odrv4 I__9701 (
            .O(N__39119),
            .I(\b2v_inst.dir_energiaZ0Z_8 ));
    Odrv4 I__9700 (
            .O(N__39116),
            .I(\b2v_inst.dir_energiaZ0Z_8 ));
    LocalMux I__9699 (
            .O(N__39113),
            .I(\b2v_inst.dir_energiaZ0Z_8 ));
    LocalMux I__9698 (
            .O(N__39110),
            .I(\b2v_inst.dir_energiaZ0Z_8 ));
    CascadeMux I__9697 (
            .O(N__39101),
            .I(N__39097));
    CascadeMux I__9696 (
            .O(N__39100),
            .I(N__39094));
    InMux I__9695 (
            .O(N__39097),
            .I(N__39091));
    InMux I__9694 (
            .O(N__39094),
            .I(N__39088));
    LocalMux I__9693 (
            .O(N__39091),
            .I(N__39085));
    LocalMux I__9692 (
            .O(N__39088),
            .I(N__39082));
    Span4Mux_v I__9691 (
            .O(N__39085),
            .I(N__39076));
    Span4Mux_v I__9690 (
            .O(N__39082),
            .I(N__39073));
    InMux I__9689 (
            .O(N__39081),
            .I(N__39070));
    InMux I__9688 (
            .O(N__39080),
            .I(N__39065));
    InMux I__9687 (
            .O(N__39079),
            .I(N__39062));
    Span4Mux_v I__9686 (
            .O(N__39076),
            .I(N__39059));
    Span4Mux_v I__9685 (
            .O(N__39073),
            .I(N__39053));
    LocalMux I__9684 (
            .O(N__39070),
            .I(N__39053));
    InMux I__9683 (
            .O(N__39069),
            .I(N__39050));
    InMux I__9682 (
            .O(N__39068),
            .I(N__39046));
    LocalMux I__9681 (
            .O(N__39065),
            .I(N__39041));
    LocalMux I__9680 (
            .O(N__39062),
            .I(N__39041));
    Span4Mux_v I__9679 (
            .O(N__39059),
            .I(N__39038));
    InMux I__9678 (
            .O(N__39058),
            .I(N__39035));
    Span4Mux_v I__9677 (
            .O(N__39053),
            .I(N__39031));
    LocalMux I__9676 (
            .O(N__39050),
            .I(N__39028));
    InMux I__9675 (
            .O(N__39049),
            .I(N__39023));
    LocalMux I__9674 (
            .O(N__39046),
            .I(N__39018));
    Span4Mux_v I__9673 (
            .O(N__39041),
            .I(N__39018));
    Span4Mux_v I__9672 (
            .O(N__39038),
            .I(N__39013));
    LocalMux I__9671 (
            .O(N__39035),
            .I(N__39013));
    InMux I__9670 (
            .O(N__39034),
            .I(N__39010));
    Span4Mux_h I__9669 (
            .O(N__39031),
            .I(N__39007));
    Span4Mux_v I__9668 (
            .O(N__39028),
            .I(N__39004));
    InMux I__9667 (
            .O(N__39027),
            .I(N__39001));
    InMux I__9666 (
            .O(N__39026),
            .I(N__38998));
    LocalMux I__9665 (
            .O(N__39023),
            .I(N__38995));
    Span4Mux_h I__9664 (
            .O(N__39018),
            .I(N__38992));
    Span4Mux_h I__9663 (
            .O(N__39013),
            .I(N__38987));
    LocalMux I__9662 (
            .O(N__39010),
            .I(N__38987));
    Span4Mux_h I__9661 (
            .O(N__39007),
            .I(N__38980));
    Span4Mux_h I__9660 (
            .O(N__39004),
            .I(N__38980));
    LocalMux I__9659 (
            .O(N__39001),
            .I(N__38980));
    LocalMux I__9658 (
            .O(N__38998),
            .I(\b2v_inst.indiceZ0Z_8 ));
    Odrv4 I__9657 (
            .O(N__38995),
            .I(\b2v_inst.indiceZ0Z_8 ));
    Odrv4 I__9656 (
            .O(N__38992),
            .I(\b2v_inst.indiceZ0Z_8 ));
    Odrv4 I__9655 (
            .O(N__38987),
            .I(\b2v_inst.indiceZ0Z_8 ));
    Odrv4 I__9654 (
            .O(N__38980),
            .I(\b2v_inst.indiceZ0Z_8 ));
    CascadeMux I__9653 (
            .O(N__38969),
            .I(N__38965));
    CascadeMux I__9652 (
            .O(N__38968),
            .I(N__38962));
    CascadeBuf I__9651 (
            .O(N__38965),
            .I(N__38959));
    CascadeBuf I__9650 (
            .O(N__38962),
            .I(N__38956));
    CascadeMux I__9649 (
            .O(N__38959),
            .I(N__38953));
    CascadeMux I__9648 (
            .O(N__38956),
            .I(N__38950));
    CascadeBuf I__9647 (
            .O(N__38953),
            .I(N__38947));
    CascadeBuf I__9646 (
            .O(N__38950),
            .I(N__38944));
    CascadeMux I__9645 (
            .O(N__38947),
            .I(N__38941));
    CascadeMux I__9644 (
            .O(N__38944),
            .I(N__38938));
    InMux I__9643 (
            .O(N__38941),
            .I(N__38935));
    InMux I__9642 (
            .O(N__38938),
            .I(N__38932));
    LocalMux I__9641 (
            .O(N__38935),
            .I(N_443_i));
    LocalMux I__9640 (
            .O(N__38932),
            .I(N_443_i));
    CascadeMux I__9639 (
            .O(N__38927),
            .I(N__38924));
    InMux I__9638 (
            .O(N__38924),
            .I(N__38921));
    LocalMux I__9637 (
            .O(N__38921),
            .I(N__38918));
    Span4Mux_v I__9636 (
            .O(N__38918),
            .I(N__38914));
    InMux I__9635 (
            .O(N__38917),
            .I(N__38911));
    Span4Mux_h I__9634 (
            .O(N__38914),
            .I(N__38906));
    LocalMux I__9633 (
            .O(N__38911),
            .I(N__38902));
    CascadeMux I__9632 (
            .O(N__38910),
            .I(N__38899));
    CascadeMux I__9631 (
            .O(N__38909),
            .I(N__38896));
    Span4Mux_h I__9630 (
            .O(N__38906),
            .I(N__38893));
    InMux I__9629 (
            .O(N__38905),
            .I(N__38890));
    Span4Mux_h I__9628 (
            .O(N__38902),
            .I(N__38887));
    InMux I__9627 (
            .O(N__38899),
            .I(N__38884));
    InMux I__9626 (
            .O(N__38896),
            .I(N__38881));
    Odrv4 I__9625 (
            .O(N__38893),
            .I(\b2v_inst.dir_energiaZ0Z_7 ));
    LocalMux I__9624 (
            .O(N__38890),
            .I(\b2v_inst.dir_energiaZ0Z_7 ));
    Odrv4 I__9623 (
            .O(N__38887),
            .I(\b2v_inst.dir_energiaZ0Z_7 ));
    LocalMux I__9622 (
            .O(N__38884),
            .I(\b2v_inst.dir_energiaZ0Z_7 ));
    LocalMux I__9621 (
            .O(N__38881),
            .I(\b2v_inst.dir_energiaZ0Z_7 ));
    InMux I__9620 (
            .O(N__38870),
            .I(N__38867));
    LocalMux I__9619 (
            .O(N__38867),
            .I(N__38863));
    InMux I__9618 (
            .O(N__38866),
            .I(N__38857));
    Span4Mux_v I__9617 (
            .O(N__38863),
            .I(N__38854));
    CascadeMux I__9616 (
            .O(N__38862),
            .I(N__38851));
    InMux I__9615 (
            .O(N__38861),
            .I(N__38848));
    CascadeMux I__9614 (
            .O(N__38860),
            .I(N__38844));
    LocalMux I__9613 (
            .O(N__38857),
            .I(N__38840));
    Sp12to4 I__9612 (
            .O(N__38854),
            .I(N__38837));
    InMux I__9611 (
            .O(N__38851),
            .I(N__38833));
    LocalMux I__9610 (
            .O(N__38848),
            .I(N__38830));
    InMux I__9609 (
            .O(N__38847),
            .I(N__38825));
    InMux I__9608 (
            .O(N__38844),
            .I(N__38822));
    InMux I__9607 (
            .O(N__38843),
            .I(N__38819));
    Span12Mux_h I__9606 (
            .O(N__38840),
            .I(N__38814));
    Span12Mux_h I__9605 (
            .O(N__38837),
            .I(N__38814));
    InMux I__9604 (
            .O(N__38836),
            .I(N__38811));
    LocalMux I__9603 (
            .O(N__38833),
            .I(N__38808));
    Span4Mux_v I__9602 (
            .O(N__38830),
            .I(N__38805));
    InMux I__9601 (
            .O(N__38829),
            .I(N__38802));
    InMux I__9600 (
            .O(N__38828),
            .I(N__38799));
    LocalMux I__9599 (
            .O(N__38825),
            .I(N__38794));
    LocalMux I__9598 (
            .O(N__38822),
            .I(N__38794));
    LocalMux I__9597 (
            .O(N__38819),
            .I(N__38790));
    Span12Mux_v I__9596 (
            .O(N__38814),
            .I(N__38785));
    LocalMux I__9595 (
            .O(N__38811),
            .I(N__38785));
    Span4Mux_v I__9594 (
            .O(N__38808),
            .I(N__38782));
    Span4Mux_h I__9593 (
            .O(N__38805),
            .I(N__38779));
    LocalMux I__9592 (
            .O(N__38802),
            .I(N__38772));
    LocalMux I__9591 (
            .O(N__38799),
            .I(N__38772));
    Span4Mux_v I__9590 (
            .O(N__38794),
            .I(N__38772));
    InMux I__9589 (
            .O(N__38793),
            .I(N__38769));
    Odrv12 I__9588 (
            .O(N__38790),
            .I(\b2v_inst.indiceZ0Z_7 ));
    Odrv12 I__9587 (
            .O(N__38785),
            .I(\b2v_inst.indiceZ0Z_7 ));
    Odrv4 I__9586 (
            .O(N__38782),
            .I(\b2v_inst.indiceZ0Z_7 ));
    Odrv4 I__9585 (
            .O(N__38779),
            .I(\b2v_inst.indiceZ0Z_7 ));
    Odrv4 I__9584 (
            .O(N__38772),
            .I(\b2v_inst.indiceZ0Z_7 ));
    LocalMux I__9583 (
            .O(N__38769),
            .I(\b2v_inst.indiceZ0Z_7 ));
    CascadeMux I__9582 (
            .O(N__38756),
            .I(N__38752));
    CascadeMux I__9581 (
            .O(N__38755),
            .I(N__38749));
    CascadeBuf I__9580 (
            .O(N__38752),
            .I(N__38746));
    CascadeBuf I__9579 (
            .O(N__38749),
            .I(N__38743));
    CascadeMux I__9578 (
            .O(N__38746),
            .I(N__38740));
    CascadeMux I__9577 (
            .O(N__38743),
            .I(N__38737));
    CascadeBuf I__9576 (
            .O(N__38740),
            .I(N__38734));
    CascadeBuf I__9575 (
            .O(N__38737),
            .I(N__38731));
    CascadeMux I__9574 (
            .O(N__38734),
            .I(N__38728));
    CascadeMux I__9573 (
            .O(N__38731),
            .I(N__38725));
    InMux I__9572 (
            .O(N__38728),
            .I(N__38722));
    InMux I__9571 (
            .O(N__38725),
            .I(N__38719));
    LocalMux I__9570 (
            .O(N__38722),
            .I(N_353_i));
    LocalMux I__9569 (
            .O(N__38719),
            .I(N_353_i));
    CascadeMux I__9568 (
            .O(N__38714),
            .I(N__38711));
    InMux I__9567 (
            .O(N__38711),
            .I(N__38708));
    LocalMux I__9566 (
            .O(N__38708),
            .I(N__38704));
    InMux I__9565 (
            .O(N__38707),
            .I(N__38701));
    Span4Mux_v I__9564 (
            .O(N__38704),
            .I(N__38698));
    LocalMux I__9563 (
            .O(N__38701),
            .I(N__38694));
    Sp12to4 I__9562 (
            .O(N__38698),
            .I(N__38689));
    InMux I__9561 (
            .O(N__38697),
            .I(N__38686));
    Span4Mux_h I__9560 (
            .O(N__38694),
            .I(N__38683));
    InMux I__9559 (
            .O(N__38693),
            .I(N__38680));
    InMux I__9558 (
            .O(N__38692),
            .I(N__38677));
    Odrv12 I__9557 (
            .O(N__38689),
            .I(\b2v_inst.dir_energiaZ0Z_1 ));
    LocalMux I__9556 (
            .O(N__38686),
            .I(\b2v_inst.dir_energiaZ0Z_1 ));
    Odrv4 I__9555 (
            .O(N__38683),
            .I(\b2v_inst.dir_energiaZ0Z_1 ));
    LocalMux I__9554 (
            .O(N__38680),
            .I(\b2v_inst.dir_energiaZ0Z_1 ));
    LocalMux I__9553 (
            .O(N__38677),
            .I(\b2v_inst.dir_energiaZ0Z_1 ));
    InMux I__9552 (
            .O(N__38666),
            .I(N__38661));
    InMux I__9551 (
            .O(N__38665),
            .I(N__38657));
    CascadeMux I__9550 (
            .O(N__38664),
            .I(N__38653));
    LocalMux I__9549 (
            .O(N__38661),
            .I(N__38650));
    InMux I__9548 (
            .O(N__38660),
            .I(N__38647));
    LocalMux I__9547 (
            .O(N__38657),
            .I(N__38643));
    InMux I__9546 (
            .O(N__38656),
            .I(N__38637));
    InMux I__9545 (
            .O(N__38653),
            .I(N__38634));
    Span4Mux_v I__9544 (
            .O(N__38650),
            .I(N__38629));
    LocalMux I__9543 (
            .O(N__38647),
            .I(N__38629));
    InMux I__9542 (
            .O(N__38646),
            .I(N__38626));
    Span4Mux_v I__9541 (
            .O(N__38643),
            .I(N__38622));
    InMux I__9540 (
            .O(N__38642),
            .I(N__38619));
    InMux I__9539 (
            .O(N__38641),
            .I(N__38616));
    InMux I__9538 (
            .O(N__38640),
            .I(N__38613));
    LocalMux I__9537 (
            .O(N__38637),
            .I(N__38610));
    LocalMux I__9536 (
            .O(N__38634),
            .I(N__38607));
    Span4Mux_v I__9535 (
            .O(N__38629),
            .I(N__38604));
    LocalMux I__9534 (
            .O(N__38626),
            .I(N__38600));
    InMux I__9533 (
            .O(N__38625),
            .I(N__38597));
    Span4Mux_v I__9532 (
            .O(N__38622),
            .I(N__38594));
    LocalMux I__9531 (
            .O(N__38619),
            .I(N__38591));
    LocalMux I__9530 (
            .O(N__38616),
            .I(N__38588));
    LocalMux I__9529 (
            .O(N__38613),
            .I(N__38584));
    Span4Mux_v I__9528 (
            .O(N__38610),
            .I(N__38579));
    Span4Mux_v I__9527 (
            .O(N__38607),
            .I(N__38579));
    Sp12to4 I__9526 (
            .O(N__38604),
            .I(N__38576));
    CascadeMux I__9525 (
            .O(N__38603),
            .I(N__38570));
    Span4Mux_v I__9524 (
            .O(N__38600),
            .I(N__38567));
    LocalMux I__9523 (
            .O(N__38597),
            .I(N__38564));
    Span4Mux_v I__9522 (
            .O(N__38594),
            .I(N__38559));
    Span4Mux_h I__9521 (
            .O(N__38591),
            .I(N__38559));
    Span4Mux_v I__9520 (
            .O(N__38588),
            .I(N__38556));
    InMux I__9519 (
            .O(N__38587),
            .I(N__38553));
    Span4Mux_v I__9518 (
            .O(N__38584),
            .I(N__38548));
    Span4Mux_h I__9517 (
            .O(N__38579),
            .I(N__38548));
    Span12Mux_h I__9516 (
            .O(N__38576),
            .I(N__38545));
    InMux I__9515 (
            .O(N__38575),
            .I(N__38540));
    InMux I__9514 (
            .O(N__38574),
            .I(N__38540));
    InMux I__9513 (
            .O(N__38573),
            .I(N__38537));
    InMux I__9512 (
            .O(N__38570),
            .I(N__38534));
    Span4Mux_h I__9511 (
            .O(N__38567),
            .I(N__38523));
    Span4Mux_v I__9510 (
            .O(N__38564),
            .I(N__38523));
    Span4Mux_v I__9509 (
            .O(N__38559),
            .I(N__38523));
    Span4Mux_h I__9508 (
            .O(N__38556),
            .I(N__38523));
    LocalMux I__9507 (
            .O(N__38553),
            .I(N__38523));
    Odrv4 I__9506 (
            .O(N__38548),
            .I(\b2v_inst.indiceZ0Z_1 ));
    Odrv12 I__9505 (
            .O(N__38545),
            .I(\b2v_inst.indiceZ0Z_1 ));
    LocalMux I__9504 (
            .O(N__38540),
            .I(\b2v_inst.indiceZ0Z_1 ));
    LocalMux I__9503 (
            .O(N__38537),
            .I(\b2v_inst.indiceZ0Z_1 ));
    LocalMux I__9502 (
            .O(N__38534),
            .I(\b2v_inst.indiceZ0Z_1 ));
    Odrv4 I__9501 (
            .O(N__38523),
            .I(\b2v_inst.indiceZ0Z_1 ));
    CascadeMux I__9500 (
            .O(N__38510),
            .I(N__38506));
    CascadeMux I__9499 (
            .O(N__38509),
            .I(N__38503));
    CascadeBuf I__9498 (
            .O(N__38506),
            .I(N__38500));
    CascadeBuf I__9497 (
            .O(N__38503),
            .I(N__38497));
    CascadeMux I__9496 (
            .O(N__38500),
            .I(N__38494));
    CascadeMux I__9495 (
            .O(N__38497),
            .I(N__38491));
    CascadeBuf I__9494 (
            .O(N__38494),
            .I(N__38488));
    CascadeBuf I__9493 (
            .O(N__38491),
            .I(N__38485));
    CascadeMux I__9492 (
            .O(N__38488),
            .I(N__38482));
    CascadeMux I__9491 (
            .O(N__38485),
            .I(N__38479));
    InMux I__9490 (
            .O(N__38482),
            .I(N__38476));
    InMux I__9489 (
            .O(N__38479),
            .I(N__38473));
    LocalMux I__9488 (
            .O(N__38476),
            .I(N_359_i));
    LocalMux I__9487 (
            .O(N__38473),
            .I(N_359_i));
    InMux I__9486 (
            .O(N__38468),
            .I(N__38447));
    InMux I__9485 (
            .O(N__38467),
            .I(N__38447));
    InMux I__9484 (
            .O(N__38466),
            .I(N__38447));
    InMux I__9483 (
            .O(N__38465),
            .I(N__38447));
    InMux I__9482 (
            .O(N__38464),
            .I(N__38447));
    InMux I__9481 (
            .O(N__38463),
            .I(N__38434));
    InMux I__9480 (
            .O(N__38462),
            .I(N__38434));
    InMux I__9479 (
            .O(N__38461),
            .I(N__38434));
    InMux I__9478 (
            .O(N__38460),
            .I(N__38434));
    InMux I__9477 (
            .O(N__38459),
            .I(N__38434));
    InMux I__9476 (
            .O(N__38458),
            .I(N__38434));
    LocalMux I__9475 (
            .O(N__38447),
            .I(\b2v_inst.N_645 ));
    LocalMux I__9474 (
            .O(N__38434),
            .I(\b2v_inst.N_645 ));
    InMux I__9473 (
            .O(N__38429),
            .I(N__38426));
    LocalMux I__9472 (
            .O(N__38426),
            .I(N__38423));
    Span4Mux_h I__9471 (
            .O(N__38423),
            .I(N__38419));
    InMux I__9470 (
            .O(N__38422),
            .I(N__38416));
    Span4Mux_h I__9469 (
            .O(N__38419),
            .I(N__38413));
    LocalMux I__9468 (
            .O(N__38416),
            .I(N__38409));
    Span4Mux_h I__9467 (
            .O(N__38413),
            .I(N__38404));
    InMux I__9466 (
            .O(N__38412),
            .I(N__38401));
    Span4Mux_h I__9465 (
            .O(N__38409),
            .I(N__38398));
    InMux I__9464 (
            .O(N__38408),
            .I(N__38395));
    InMux I__9463 (
            .O(N__38407),
            .I(N__38392));
    Odrv4 I__9462 (
            .O(N__38404),
            .I(\b2v_inst.dir_energiaZ0Z_6 ));
    LocalMux I__9461 (
            .O(N__38401),
            .I(\b2v_inst.dir_energiaZ0Z_6 ));
    Odrv4 I__9460 (
            .O(N__38398),
            .I(\b2v_inst.dir_energiaZ0Z_6 ));
    LocalMux I__9459 (
            .O(N__38395),
            .I(\b2v_inst.dir_energiaZ0Z_6 ));
    LocalMux I__9458 (
            .O(N__38392),
            .I(\b2v_inst.dir_energiaZ0Z_6 ));
    CascadeMux I__9457 (
            .O(N__38381),
            .I(N__38378));
    InMux I__9456 (
            .O(N__38378),
            .I(N__38374));
    InMux I__9455 (
            .O(N__38377),
            .I(N__38371));
    LocalMux I__9454 (
            .O(N__38374),
            .I(N__38366));
    LocalMux I__9453 (
            .O(N__38371),
            .I(N__38363));
    InMux I__9452 (
            .O(N__38370),
            .I(N__38360));
    InMux I__9451 (
            .O(N__38369),
            .I(N__38356));
    Span4Mux_h I__9450 (
            .O(N__38366),
            .I(N__38352));
    Span4Mux_v I__9449 (
            .O(N__38363),
            .I(N__38349));
    LocalMux I__9448 (
            .O(N__38360),
            .I(N__38346));
    InMux I__9447 (
            .O(N__38359),
            .I(N__38343));
    LocalMux I__9446 (
            .O(N__38356),
            .I(N__38339));
    InMux I__9445 (
            .O(N__38355),
            .I(N__38334));
    Sp12to4 I__9444 (
            .O(N__38352),
            .I(N__38331));
    Span4Mux_v I__9443 (
            .O(N__38349),
            .I(N__38328));
    Span4Mux_v I__9442 (
            .O(N__38346),
            .I(N__38323));
    LocalMux I__9441 (
            .O(N__38343),
            .I(N__38320));
    InMux I__9440 (
            .O(N__38342),
            .I(N__38317));
    Sp12to4 I__9439 (
            .O(N__38339),
            .I(N__38314));
    InMux I__9438 (
            .O(N__38338),
            .I(N__38310));
    InMux I__9437 (
            .O(N__38337),
            .I(N__38307));
    LocalMux I__9436 (
            .O(N__38334),
            .I(N__38300));
    Span12Mux_v I__9435 (
            .O(N__38331),
            .I(N__38300));
    Sp12to4 I__9434 (
            .O(N__38328),
            .I(N__38300));
    InMux I__9433 (
            .O(N__38327),
            .I(N__38297));
    InMux I__9432 (
            .O(N__38326),
            .I(N__38294));
    Span4Mux_h I__9431 (
            .O(N__38323),
            .I(N__38289));
    Span4Mux_v I__9430 (
            .O(N__38320),
            .I(N__38289));
    LocalMux I__9429 (
            .O(N__38317),
            .I(N__38284));
    Span12Mux_v I__9428 (
            .O(N__38314),
            .I(N__38284));
    InMux I__9427 (
            .O(N__38313),
            .I(N__38281));
    LocalMux I__9426 (
            .O(N__38310),
            .I(\b2v_inst.indiceZ0Z_6 ));
    LocalMux I__9425 (
            .O(N__38307),
            .I(\b2v_inst.indiceZ0Z_6 ));
    Odrv12 I__9424 (
            .O(N__38300),
            .I(\b2v_inst.indiceZ0Z_6 ));
    LocalMux I__9423 (
            .O(N__38297),
            .I(\b2v_inst.indiceZ0Z_6 ));
    LocalMux I__9422 (
            .O(N__38294),
            .I(\b2v_inst.indiceZ0Z_6 ));
    Odrv4 I__9421 (
            .O(N__38289),
            .I(\b2v_inst.indiceZ0Z_6 ));
    Odrv12 I__9420 (
            .O(N__38284),
            .I(\b2v_inst.indiceZ0Z_6 ));
    LocalMux I__9419 (
            .O(N__38281),
            .I(\b2v_inst.indiceZ0Z_6 ));
    InMux I__9418 (
            .O(N__38264),
            .I(N__38248));
    InMux I__9417 (
            .O(N__38263),
            .I(N__38248));
    InMux I__9416 (
            .O(N__38262),
            .I(N__38248));
    InMux I__9415 (
            .O(N__38261),
            .I(N__38248));
    InMux I__9414 (
            .O(N__38260),
            .I(N__38248));
    InMux I__9413 (
            .O(N__38259),
            .I(N__38239));
    LocalMux I__9412 (
            .O(N__38248),
            .I(N__38236));
    InMux I__9411 (
            .O(N__38247),
            .I(N__38231));
    InMux I__9410 (
            .O(N__38246),
            .I(N__38231));
    InMux I__9409 (
            .O(N__38245),
            .I(N__38222));
    InMux I__9408 (
            .O(N__38244),
            .I(N__38222));
    InMux I__9407 (
            .O(N__38243),
            .I(N__38222));
    InMux I__9406 (
            .O(N__38242),
            .I(N__38222));
    LocalMux I__9405 (
            .O(N__38239),
            .I(N__38219));
    Span4Mux_v I__9404 (
            .O(N__38236),
            .I(N__38212));
    LocalMux I__9403 (
            .O(N__38231),
            .I(N__38212));
    LocalMux I__9402 (
            .O(N__38222),
            .I(N__38212));
    Span4Mux_h I__9401 (
            .O(N__38219),
            .I(N__38209));
    Span4Mux_h I__9400 (
            .O(N__38212),
            .I(N__38206));
    Span4Mux_h I__9399 (
            .O(N__38209),
            .I(N__38203));
    Odrv4 I__9398 (
            .O(N__38206),
            .I(\b2v_inst.N_484 ));
    Odrv4 I__9397 (
            .O(N__38203),
            .I(\b2v_inst.N_484 ));
    CascadeMux I__9396 (
            .O(N__38198),
            .I(N__38194));
    CascadeMux I__9395 (
            .O(N__38197),
            .I(N__38191));
    CascadeBuf I__9394 (
            .O(N__38194),
            .I(N__38188));
    CascadeBuf I__9393 (
            .O(N__38191),
            .I(N__38185));
    CascadeMux I__9392 (
            .O(N__38188),
            .I(N__38182));
    CascadeMux I__9391 (
            .O(N__38185),
            .I(N__38179));
    CascadeBuf I__9390 (
            .O(N__38182),
            .I(N__38176));
    CascadeBuf I__9389 (
            .O(N__38179),
            .I(N__38173));
    CascadeMux I__9388 (
            .O(N__38176),
            .I(N__38170));
    CascadeMux I__9387 (
            .O(N__38173),
            .I(N__38167));
    InMux I__9386 (
            .O(N__38170),
            .I(N__38164));
    InMux I__9385 (
            .O(N__38167),
            .I(N__38161));
    LocalMux I__9384 (
            .O(N__38164),
            .I(N_354_i));
    LocalMux I__9383 (
            .O(N__38161),
            .I(N_354_i));
    CascadeMux I__9382 (
            .O(N__38156),
            .I(N__38152));
    InMux I__9381 (
            .O(N__38155),
            .I(N__38145));
    InMux I__9380 (
            .O(N__38152),
            .I(N__38145));
    InMux I__9379 (
            .O(N__38151),
            .I(N__38140));
    InMux I__9378 (
            .O(N__38150),
            .I(N__38140));
    LocalMux I__9377 (
            .O(N__38145),
            .I(N__38125));
    LocalMux I__9376 (
            .O(N__38140),
            .I(N__38120));
    SRMux I__9375 (
            .O(N__38139),
            .I(N__37847));
    SRMux I__9374 (
            .O(N__38138),
            .I(N__37847));
    SRMux I__9373 (
            .O(N__38137),
            .I(N__37847));
    SRMux I__9372 (
            .O(N__38136),
            .I(N__37847));
    SRMux I__9371 (
            .O(N__38135),
            .I(N__37847));
    SRMux I__9370 (
            .O(N__38134),
            .I(N__37847));
    SRMux I__9369 (
            .O(N__38133),
            .I(N__37847));
    SRMux I__9368 (
            .O(N__38132),
            .I(N__37847));
    SRMux I__9367 (
            .O(N__38131),
            .I(N__37847));
    SRMux I__9366 (
            .O(N__38130),
            .I(N__37847));
    SRMux I__9365 (
            .O(N__38129),
            .I(N__37847));
    SRMux I__9364 (
            .O(N__38128),
            .I(N__37847));
    Glb2LocalMux I__9363 (
            .O(N__38125),
            .I(N__37847));
    SRMux I__9362 (
            .O(N__38124),
            .I(N__37847));
    SRMux I__9361 (
            .O(N__38123),
            .I(N__37847));
    Glb2LocalMux I__9360 (
            .O(N__38120),
            .I(N__37847));
    SRMux I__9359 (
            .O(N__38119),
            .I(N__37847));
    SRMux I__9358 (
            .O(N__38118),
            .I(N__37847));
    SRMux I__9357 (
            .O(N__38117),
            .I(N__37847));
    SRMux I__9356 (
            .O(N__38116),
            .I(N__37847));
    SRMux I__9355 (
            .O(N__38115),
            .I(N__37847));
    SRMux I__9354 (
            .O(N__38114),
            .I(N__37847));
    SRMux I__9353 (
            .O(N__38113),
            .I(N__37847));
    SRMux I__9352 (
            .O(N__38112),
            .I(N__37847));
    SRMux I__9351 (
            .O(N__38111),
            .I(N__37847));
    SRMux I__9350 (
            .O(N__38110),
            .I(N__37847));
    SRMux I__9349 (
            .O(N__38109),
            .I(N__37847));
    SRMux I__9348 (
            .O(N__38108),
            .I(N__37847));
    SRMux I__9347 (
            .O(N__38107),
            .I(N__37847));
    SRMux I__9346 (
            .O(N__38106),
            .I(N__37847));
    SRMux I__9345 (
            .O(N__38105),
            .I(N__37847));
    SRMux I__9344 (
            .O(N__38104),
            .I(N__37847));
    SRMux I__9343 (
            .O(N__38103),
            .I(N__37847));
    SRMux I__9342 (
            .O(N__38102),
            .I(N__37847));
    SRMux I__9341 (
            .O(N__38101),
            .I(N__37847));
    SRMux I__9340 (
            .O(N__38100),
            .I(N__37847));
    SRMux I__9339 (
            .O(N__38099),
            .I(N__37847));
    SRMux I__9338 (
            .O(N__38098),
            .I(N__37847));
    SRMux I__9337 (
            .O(N__38097),
            .I(N__37847));
    SRMux I__9336 (
            .O(N__38096),
            .I(N__37847));
    SRMux I__9335 (
            .O(N__38095),
            .I(N__37847));
    SRMux I__9334 (
            .O(N__38094),
            .I(N__37847));
    SRMux I__9333 (
            .O(N__38093),
            .I(N__37847));
    SRMux I__9332 (
            .O(N__38092),
            .I(N__37847));
    SRMux I__9331 (
            .O(N__38091),
            .I(N__37847));
    SRMux I__9330 (
            .O(N__38090),
            .I(N__37847));
    SRMux I__9329 (
            .O(N__38089),
            .I(N__37847));
    SRMux I__9328 (
            .O(N__38088),
            .I(N__37847));
    SRMux I__9327 (
            .O(N__38087),
            .I(N__37847));
    SRMux I__9326 (
            .O(N__38086),
            .I(N__37847));
    SRMux I__9325 (
            .O(N__38085),
            .I(N__37847));
    SRMux I__9324 (
            .O(N__38084),
            .I(N__37847));
    SRMux I__9323 (
            .O(N__38083),
            .I(N__37847));
    SRMux I__9322 (
            .O(N__38082),
            .I(N__37847));
    SRMux I__9321 (
            .O(N__38081),
            .I(N__37847));
    SRMux I__9320 (
            .O(N__38080),
            .I(N__37847));
    SRMux I__9319 (
            .O(N__38079),
            .I(N__37847));
    SRMux I__9318 (
            .O(N__38078),
            .I(N__37847));
    SRMux I__9317 (
            .O(N__38077),
            .I(N__37847));
    SRMux I__9316 (
            .O(N__38076),
            .I(N__37847));
    SRMux I__9315 (
            .O(N__38075),
            .I(N__37847));
    SRMux I__9314 (
            .O(N__38074),
            .I(N__37847));
    SRMux I__9313 (
            .O(N__38073),
            .I(N__37847));
    SRMux I__9312 (
            .O(N__38072),
            .I(N__37847));
    SRMux I__9311 (
            .O(N__38071),
            .I(N__37847));
    SRMux I__9310 (
            .O(N__38070),
            .I(N__37847));
    SRMux I__9309 (
            .O(N__38069),
            .I(N__37847));
    SRMux I__9308 (
            .O(N__38068),
            .I(N__37847));
    SRMux I__9307 (
            .O(N__38067),
            .I(N__37847));
    SRMux I__9306 (
            .O(N__38066),
            .I(N__37847));
    SRMux I__9305 (
            .O(N__38065),
            .I(N__37847));
    SRMux I__9304 (
            .O(N__38064),
            .I(N__37847));
    SRMux I__9303 (
            .O(N__38063),
            .I(N__37847));
    SRMux I__9302 (
            .O(N__38062),
            .I(N__37847));
    SRMux I__9301 (
            .O(N__38061),
            .I(N__37847));
    SRMux I__9300 (
            .O(N__38060),
            .I(N__37847));
    SRMux I__9299 (
            .O(N__38059),
            .I(N__37847));
    SRMux I__9298 (
            .O(N__38058),
            .I(N__37847));
    SRMux I__9297 (
            .O(N__38057),
            .I(N__37847));
    SRMux I__9296 (
            .O(N__38056),
            .I(N__37847));
    SRMux I__9295 (
            .O(N__38055),
            .I(N__37847));
    SRMux I__9294 (
            .O(N__38054),
            .I(N__37847));
    SRMux I__9293 (
            .O(N__38053),
            .I(N__37847));
    SRMux I__9292 (
            .O(N__38052),
            .I(N__37847));
    SRMux I__9291 (
            .O(N__38051),
            .I(N__37847));
    SRMux I__9290 (
            .O(N__38050),
            .I(N__37847));
    SRMux I__9289 (
            .O(N__38049),
            .I(N__37847));
    SRMux I__9288 (
            .O(N__38048),
            .I(N__37847));
    SRMux I__9287 (
            .O(N__38047),
            .I(N__37847));
    SRMux I__9286 (
            .O(N__38046),
            .I(N__37847));
    SRMux I__9285 (
            .O(N__38045),
            .I(N__37847));
    SRMux I__9284 (
            .O(N__38044),
            .I(N__37847));
    SRMux I__9283 (
            .O(N__38043),
            .I(N__37847));
    SRMux I__9282 (
            .O(N__38042),
            .I(N__37847));
    SRMux I__9281 (
            .O(N__38041),
            .I(N__37847));
    SRMux I__9280 (
            .O(N__38040),
            .I(N__37847));
    GlobalMux I__9279 (
            .O(N__37847),
            .I(N__37844));
    gio2CtrlBuf I__9278 (
            .O(N__37844),
            .I(reset_c_i_g));
    InMux I__9277 (
            .O(N__37841),
            .I(N__37837));
    CascadeMux I__9276 (
            .O(N__37840),
            .I(N__37832));
    LocalMux I__9275 (
            .O(N__37837),
            .I(N__37827));
    InMux I__9274 (
            .O(N__37836),
            .I(N__37824));
    CascadeMux I__9273 (
            .O(N__37835),
            .I(N__37820));
    InMux I__9272 (
            .O(N__37832),
            .I(N__37814));
    InMux I__9271 (
            .O(N__37831),
            .I(N__37814));
    CascadeMux I__9270 (
            .O(N__37830),
            .I(N__37810));
    Span4Mux_v I__9269 (
            .O(N__37827),
            .I(N__37802));
    LocalMux I__9268 (
            .O(N__37824),
            .I(N__37802));
    InMux I__9267 (
            .O(N__37823),
            .I(N__37799));
    InMux I__9266 (
            .O(N__37820),
            .I(N__37794));
    InMux I__9265 (
            .O(N__37819),
            .I(N__37794));
    LocalMux I__9264 (
            .O(N__37814),
            .I(N__37786));
    InMux I__9263 (
            .O(N__37813),
            .I(N__37783));
    InMux I__9262 (
            .O(N__37810),
            .I(N__37778));
    InMux I__9261 (
            .O(N__37809),
            .I(N__37778));
    InMux I__9260 (
            .O(N__37808),
            .I(N__37773));
    InMux I__9259 (
            .O(N__37807),
            .I(N__37773));
    Span4Mux_v I__9258 (
            .O(N__37802),
            .I(N__37766));
    LocalMux I__9257 (
            .O(N__37799),
            .I(N__37766));
    LocalMux I__9256 (
            .O(N__37794),
            .I(N__37766));
    InMux I__9255 (
            .O(N__37793),
            .I(N__37763));
    InMux I__9254 (
            .O(N__37792),
            .I(N__37760));
    InMux I__9253 (
            .O(N__37791),
            .I(N__37754));
    InMux I__9252 (
            .O(N__37790),
            .I(N__37754));
    InMux I__9251 (
            .O(N__37789),
            .I(N__37750));
    Span4Mux_h I__9250 (
            .O(N__37786),
            .I(N__37741));
    LocalMux I__9249 (
            .O(N__37783),
            .I(N__37741));
    LocalMux I__9248 (
            .O(N__37778),
            .I(N__37741));
    LocalMux I__9247 (
            .O(N__37773),
            .I(N__37741));
    Span4Mux_v I__9246 (
            .O(N__37766),
            .I(N__37734));
    LocalMux I__9245 (
            .O(N__37763),
            .I(N__37734));
    LocalMux I__9244 (
            .O(N__37760),
            .I(N__37734));
    CascadeMux I__9243 (
            .O(N__37759),
            .I(N__37729));
    LocalMux I__9242 (
            .O(N__37754),
            .I(N__37725));
    InMux I__9241 (
            .O(N__37753),
            .I(N__37722));
    LocalMux I__9240 (
            .O(N__37750),
            .I(N__37719));
    Span4Mux_v I__9239 (
            .O(N__37741),
            .I(N__37716));
    Span4Mux_v I__9238 (
            .O(N__37734),
            .I(N__37713));
    InMux I__9237 (
            .O(N__37733),
            .I(N__37710));
    InMux I__9236 (
            .O(N__37732),
            .I(N__37706));
    InMux I__9235 (
            .O(N__37729),
            .I(N__37701));
    InMux I__9234 (
            .O(N__37728),
            .I(N__37701));
    Span4Mux_v I__9233 (
            .O(N__37725),
            .I(N__37698));
    LocalMux I__9232 (
            .O(N__37722),
            .I(N__37695));
    Span4Mux_v I__9231 (
            .O(N__37719),
            .I(N__37692));
    Span4Mux_h I__9230 (
            .O(N__37716),
            .I(N__37685));
    Span4Mux_h I__9229 (
            .O(N__37713),
            .I(N__37685));
    LocalMux I__9228 (
            .O(N__37710),
            .I(N__37685));
    CascadeMux I__9227 (
            .O(N__37709),
            .I(N__37682));
    LocalMux I__9226 (
            .O(N__37706),
            .I(N__37673));
    LocalMux I__9225 (
            .O(N__37701),
            .I(N__37673));
    Span4Mux_h I__9224 (
            .O(N__37698),
            .I(N__37664));
    Span4Mux_v I__9223 (
            .O(N__37695),
            .I(N__37664));
    Span4Mux_h I__9222 (
            .O(N__37692),
            .I(N__37664));
    Span4Mux_h I__9221 (
            .O(N__37685),
            .I(N__37664));
    InMux I__9220 (
            .O(N__37682),
            .I(N__37661));
    InMux I__9219 (
            .O(N__37681),
            .I(N__37658));
    InMux I__9218 (
            .O(N__37680),
            .I(N__37653));
    InMux I__9217 (
            .O(N__37679),
            .I(N__37653));
    InMux I__9216 (
            .O(N__37678),
            .I(N__37650));
    Odrv12 I__9215 (
            .O(N__37673),
            .I(\b2v_inst.N_828 ));
    Odrv4 I__9214 (
            .O(N__37664),
            .I(\b2v_inst.N_828 ));
    LocalMux I__9213 (
            .O(N__37661),
            .I(\b2v_inst.N_828 ));
    LocalMux I__9212 (
            .O(N__37658),
            .I(\b2v_inst.N_828 ));
    LocalMux I__9211 (
            .O(N__37653),
            .I(\b2v_inst.N_828 ));
    LocalMux I__9210 (
            .O(N__37650),
            .I(\b2v_inst.N_828 ));
    InMux I__9209 (
            .O(N__37637),
            .I(N__37634));
    LocalMux I__9208 (
            .O(N__37634),
            .I(\b2v_inst.un16_data_ram_cantidad_o_cry_4_c_RNIDGFOZ0 ));
    CascadeMux I__9207 (
            .O(N__37631),
            .I(N__37628));
    InMux I__9206 (
            .O(N__37628),
            .I(N__37623));
    CascadeMux I__9205 (
            .O(N__37627),
            .I(N__37620));
    CascadeMux I__9204 (
            .O(N__37626),
            .I(N__37617));
    LocalMux I__9203 (
            .O(N__37623),
            .I(N__37614));
    InMux I__9202 (
            .O(N__37620),
            .I(N__37611));
    InMux I__9201 (
            .O(N__37617),
            .I(N__37608));
    Span4Mux_v I__9200 (
            .O(N__37614),
            .I(N__37605));
    LocalMux I__9199 (
            .O(N__37611),
            .I(N__37602));
    LocalMux I__9198 (
            .O(N__37608),
            .I(N__37599));
    Span4Mux_h I__9197 (
            .O(N__37605),
            .I(N__37594));
    Span4Mux_h I__9196 (
            .O(N__37602),
            .I(N__37591));
    Span4Mux_v I__9195 (
            .O(N__37599),
            .I(N__37588));
    InMux I__9194 (
            .O(N__37598),
            .I(N__37585));
    InMux I__9193 (
            .O(N__37597),
            .I(N__37582));
    Span4Mux_h I__9192 (
            .O(N__37594),
            .I(N__37573));
    Span4Mux_v I__9191 (
            .O(N__37591),
            .I(N__37573));
    Span4Mux_h I__9190 (
            .O(N__37588),
            .I(N__37573));
    LocalMux I__9189 (
            .O(N__37585),
            .I(N__37573));
    LocalMux I__9188 (
            .O(N__37582),
            .I(N__37570));
    Span4Mux_h I__9187 (
            .O(N__37573),
            .I(N__37567));
    Odrv12 I__9186 (
            .O(N__37570),
            .I(b2v_inst_data_a_escribir_5));
    Odrv4 I__9185 (
            .O(N__37567),
            .I(b2v_inst_data_a_escribir_5));
    InMux I__9184 (
            .O(N__37562),
            .I(N__37557));
    InMux I__9183 (
            .O(N__37561),
            .I(N__37554));
    CascadeMux I__9182 (
            .O(N__37560),
            .I(N__37551));
    LocalMux I__9181 (
            .O(N__37557),
            .I(N__37540));
    LocalMux I__9180 (
            .O(N__37554),
            .I(N__37537));
    InMux I__9179 (
            .O(N__37551),
            .I(N__37532));
    InMux I__9178 (
            .O(N__37550),
            .I(N__37532));
    InMux I__9177 (
            .O(N__37549),
            .I(N__37527));
    InMux I__9176 (
            .O(N__37548),
            .I(N__37524));
    InMux I__9175 (
            .O(N__37547),
            .I(N__37521));
    InMux I__9174 (
            .O(N__37546),
            .I(N__37516));
    InMux I__9173 (
            .O(N__37545),
            .I(N__37516));
    InMux I__9172 (
            .O(N__37544),
            .I(N__37511));
    InMux I__9171 (
            .O(N__37543),
            .I(N__37511));
    Span4Mux_v I__9170 (
            .O(N__37540),
            .I(N__37504));
    Span4Mux_h I__9169 (
            .O(N__37537),
            .I(N__37504));
    LocalMux I__9168 (
            .O(N__37532),
            .I(N__37499));
    InMux I__9167 (
            .O(N__37531),
            .I(N__37491));
    InMux I__9166 (
            .O(N__37530),
            .I(N__37491));
    LocalMux I__9165 (
            .O(N__37527),
            .I(N__37480));
    LocalMux I__9164 (
            .O(N__37524),
            .I(N__37480));
    LocalMux I__9163 (
            .O(N__37521),
            .I(N__37480));
    LocalMux I__9162 (
            .O(N__37516),
            .I(N__37480));
    LocalMux I__9161 (
            .O(N__37511),
            .I(N__37480));
    InMux I__9160 (
            .O(N__37510),
            .I(N__37474));
    InMux I__9159 (
            .O(N__37509),
            .I(N__37474));
    Span4Mux_h I__9158 (
            .O(N__37504),
            .I(N__37471));
    InMux I__9157 (
            .O(N__37503),
            .I(N__37468));
    InMux I__9156 (
            .O(N__37502),
            .I(N__37462));
    Span4Mux_h I__9155 (
            .O(N__37499),
            .I(N__37456));
    InMux I__9154 (
            .O(N__37498),
            .I(N__37453));
    InMux I__9153 (
            .O(N__37497),
            .I(N__37450));
    InMux I__9152 (
            .O(N__37496),
            .I(N__37446));
    LocalMux I__9151 (
            .O(N__37491),
            .I(N__37441));
    Span4Mux_v I__9150 (
            .O(N__37480),
            .I(N__37441));
    InMux I__9149 (
            .O(N__37479),
            .I(N__37438));
    LocalMux I__9148 (
            .O(N__37474),
            .I(N__37431));
    Span4Mux_h I__9147 (
            .O(N__37471),
            .I(N__37431));
    LocalMux I__9146 (
            .O(N__37468),
            .I(N__37431));
    InMux I__9145 (
            .O(N__37467),
            .I(N__37426));
    InMux I__9144 (
            .O(N__37466),
            .I(N__37426));
    InMux I__9143 (
            .O(N__37465),
            .I(N__37423));
    LocalMux I__9142 (
            .O(N__37462),
            .I(N__37420));
    InMux I__9141 (
            .O(N__37461),
            .I(N__37415));
    InMux I__9140 (
            .O(N__37460),
            .I(N__37415));
    InMux I__9139 (
            .O(N__37459),
            .I(N__37412));
    Span4Mux_v I__9138 (
            .O(N__37456),
            .I(N__37407));
    LocalMux I__9137 (
            .O(N__37453),
            .I(N__37407));
    LocalMux I__9136 (
            .O(N__37450),
            .I(N__37401));
    InMux I__9135 (
            .O(N__37449),
            .I(N__37398));
    LocalMux I__9134 (
            .O(N__37446),
            .I(N__37393));
    Span4Mux_h I__9133 (
            .O(N__37441),
            .I(N__37390));
    LocalMux I__9132 (
            .O(N__37438),
            .I(N__37385));
    Span4Mux_v I__9131 (
            .O(N__37431),
            .I(N__37385));
    LocalMux I__9130 (
            .O(N__37426),
            .I(N__37381));
    LocalMux I__9129 (
            .O(N__37423),
            .I(N__37370));
    Span4Mux_v I__9128 (
            .O(N__37420),
            .I(N__37370));
    LocalMux I__9127 (
            .O(N__37415),
            .I(N__37370));
    LocalMux I__9126 (
            .O(N__37412),
            .I(N__37370));
    Span4Mux_h I__9125 (
            .O(N__37407),
            .I(N__37370));
    InMux I__9124 (
            .O(N__37406),
            .I(N__37365));
    InMux I__9123 (
            .O(N__37405),
            .I(N__37365));
    InMux I__9122 (
            .O(N__37404),
            .I(N__37362));
    Span12Mux_h I__9121 (
            .O(N__37401),
            .I(N__37359));
    LocalMux I__9120 (
            .O(N__37398),
            .I(N__37356));
    InMux I__9119 (
            .O(N__37397),
            .I(N__37351));
    InMux I__9118 (
            .O(N__37396),
            .I(N__37351));
    Span4Mux_h I__9117 (
            .O(N__37393),
            .I(N__37348));
    Span4Mux_h I__9116 (
            .O(N__37390),
            .I(N__37343));
    Span4Mux_v I__9115 (
            .O(N__37385),
            .I(N__37343));
    InMux I__9114 (
            .O(N__37384),
            .I(N__37340));
    Span4Mux_h I__9113 (
            .O(N__37381),
            .I(N__37335));
    Span4Mux_h I__9112 (
            .O(N__37370),
            .I(N__37335));
    LocalMux I__9111 (
            .O(N__37365),
            .I(\b2v_inst.N_514 ));
    LocalMux I__9110 (
            .O(N__37362),
            .I(\b2v_inst.N_514 ));
    Odrv12 I__9109 (
            .O(N__37359),
            .I(\b2v_inst.N_514 ));
    Odrv4 I__9108 (
            .O(N__37356),
            .I(\b2v_inst.N_514 ));
    LocalMux I__9107 (
            .O(N__37351),
            .I(\b2v_inst.N_514 ));
    Odrv4 I__9106 (
            .O(N__37348),
            .I(\b2v_inst.N_514 ));
    Odrv4 I__9105 (
            .O(N__37343),
            .I(\b2v_inst.N_514 ));
    LocalMux I__9104 (
            .O(N__37340),
            .I(\b2v_inst.N_514 ));
    Odrv4 I__9103 (
            .O(N__37335),
            .I(\b2v_inst.N_514 ));
    InMux I__9102 (
            .O(N__37316),
            .I(N__37313));
    LocalMux I__9101 (
            .O(N__37313),
            .I(N__37310));
    Odrv4 I__9100 (
            .O(N__37310),
            .I(N_547_i));
    CascadeMux I__9099 (
            .O(N__37307),
            .I(N__37304));
    InMux I__9098 (
            .O(N__37304),
            .I(N__37293));
    CascadeMux I__9097 (
            .O(N__37303),
            .I(N__37289));
    InMux I__9096 (
            .O(N__37302),
            .I(N__37273));
    InMux I__9095 (
            .O(N__37301),
            .I(N__37273));
    InMux I__9094 (
            .O(N__37300),
            .I(N__37273));
    InMux I__9093 (
            .O(N__37299),
            .I(N__37273));
    InMux I__9092 (
            .O(N__37298),
            .I(N__37266));
    InMux I__9091 (
            .O(N__37297),
            .I(N__37266));
    InMux I__9090 (
            .O(N__37296),
            .I(N__37266));
    LocalMux I__9089 (
            .O(N__37293),
            .I(N__37260));
    SRMux I__9088 (
            .O(N__37292),
            .I(N__37257));
    InMux I__9087 (
            .O(N__37289),
            .I(N__37253));
    CascadeMux I__9086 (
            .O(N__37288),
            .I(N__37250));
    SRMux I__9085 (
            .O(N__37287),
            .I(N__37246));
    SRMux I__9084 (
            .O(N__37286),
            .I(N__37243));
    SRMux I__9083 (
            .O(N__37285),
            .I(N__37239));
    SRMux I__9082 (
            .O(N__37284),
            .I(N__37236));
    SRMux I__9081 (
            .O(N__37283),
            .I(N__37232));
    SRMux I__9080 (
            .O(N__37282),
            .I(N__37228));
    LocalMux I__9079 (
            .O(N__37273),
            .I(N__37221));
    LocalMux I__9078 (
            .O(N__37266),
            .I(N__37221));
    InMux I__9077 (
            .O(N__37265),
            .I(N__37218));
    InMux I__9076 (
            .O(N__37264),
            .I(N__37214));
    InMux I__9075 (
            .O(N__37263),
            .I(N__37209));
    Span4Mux_v I__9074 (
            .O(N__37260),
            .I(N__37206));
    LocalMux I__9073 (
            .O(N__37257),
            .I(N__37203));
    SRMux I__9072 (
            .O(N__37256),
            .I(N__37200));
    LocalMux I__9071 (
            .O(N__37253),
            .I(N__37195));
    InMux I__9070 (
            .O(N__37250),
            .I(N__37192));
    SRMux I__9069 (
            .O(N__37249),
            .I(N__37189));
    LocalMux I__9068 (
            .O(N__37246),
            .I(N__37184));
    LocalMux I__9067 (
            .O(N__37243),
            .I(N__37184));
    SRMux I__9066 (
            .O(N__37242),
            .I(N__37181));
    LocalMux I__9065 (
            .O(N__37239),
            .I(N__37176));
    LocalMux I__9064 (
            .O(N__37236),
            .I(N__37176));
    SRMux I__9063 (
            .O(N__37235),
            .I(N__37173));
    LocalMux I__9062 (
            .O(N__37232),
            .I(N__37170));
    SRMux I__9061 (
            .O(N__37231),
            .I(N__37167));
    LocalMux I__9060 (
            .O(N__37228),
            .I(N__37164));
    SRMux I__9059 (
            .O(N__37227),
            .I(N__37161));
    SRMux I__9058 (
            .O(N__37226),
            .I(N__37148));
    Span4Mux_h I__9057 (
            .O(N__37221),
            .I(N__37143));
    LocalMux I__9056 (
            .O(N__37218),
            .I(N__37143));
    InMux I__9055 (
            .O(N__37217),
            .I(N__37140));
    LocalMux I__9054 (
            .O(N__37214),
            .I(N__37137));
    SRMux I__9053 (
            .O(N__37213),
            .I(N__37134));
    SRMux I__9052 (
            .O(N__37212),
            .I(N__37130));
    LocalMux I__9051 (
            .O(N__37209),
            .I(N__37126));
    Span4Mux_h I__9050 (
            .O(N__37206),
            .I(N__37119));
    Span4Mux_v I__9049 (
            .O(N__37203),
            .I(N__37119));
    LocalMux I__9048 (
            .O(N__37200),
            .I(N__37119));
    SRMux I__9047 (
            .O(N__37199),
            .I(N__37116));
    SRMux I__9046 (
            .O(N__37198),
            .I(N__37113));
    Span4Mux_h I__9045 (
            .O(N__37195),
            .I(N__37107));
    LocalMux I__9044 (
            .O(N__37192),
            .I(N__37107));
    LocalMux I__9043 (
            .O(N__37189),
            .I(N__37100));
    Span4Mux_v I__9042 (
            .O(N__37184),
            .I(N__37100));
    LocalMux I__9041 (
            .O(N__37181),
            .I(N__37100));
    Span4Mux_v I__9040 (
            .O(N__37176),
            .I(N__37095));
    LocalMux I__9039 (
            .O(N__37173),
            .I(N__37095));
    Span4Mux_v I__9038 (
            .O(N__37170),
            .I(N__37090));
    LocalMux I__9037 (
            .O(N__37167),
            .I(N__37090));
    Span4Mux_v I__9036 (
            .O(N__37164),
            .I(N__37085));
    LocalMux I__9035 (
            .O(N__37161),
            .I(N__37085));
    SRMux I__9034 (
            .O(N__37160),
            .I(N__37082));
    CascadeMux I__9033 (
            .O(N__37159),
            .I(N__37079));
    CascadeMux I__9032 (
            .O(N__37158),
            .I(N__37076));
    CascadeMux I__9031 (
            .O(N__37157),
            .I(N__37073));
    CascadeMux I__9030 (
            .O(N__37156),
            .I(N__37070));
    CascadeMux I__9029 (
            .O(N__37155),
            .I(N__37067));
    CascadeMux I__9028 (
            .O(N__37154),
            .I(N__37064));
    CascadeMux I__9027 (
            .O(N__37153),
            .I(N__37060));
    CascadeMux I__9026 (
            .O(N__37152),
            .I(N__37057));
    CascadeMux I__9025 (
            .O(N__37151),
            .I(N__37053));
    LocalMux I__9024 (
            .O(N__37148),
            .I(N__37050));
    Span4Mux_v I__9023 (
            .O(N__37143),
            .I(N__37047));
    LocalMux I__9022 (
            .O(N__37140),
            .I(N__37044));
    Span4Mux_v I__9021 (
            .O(N__37137),
            .I(N__37039));
    LocalMux I__9020 (
            .O(N__37134),
            .I(N__37039));
    CascadeMux I__9019 (
            .O(N__37133),
            .I(N__37036));
    LocalMux I__9018 (
            .O(N__37130),
            .I(N__37033));
    SRMux I__9017 (
            .O(N__37129),
            .I(N__37030));
    Span4Mux_v I__9016 (
            .O(N__37126),
            .I(N__37026));
    Span4Mux_h I__9015 (
            .O(N__37119),
            .I(N__37019));
    LocalMux I__9014 (
            .O(N__37116),
            .I(N__37019));
    LocalMux I__9013 (
            .O(N__37113),
            .I(N__37019));
    SRMux I__9012 (
            .O(N__37112),
            .I(N__37016));
    Span4Mux_v I__9011 (
            .O(N__37107),
            .I(N__37009));
    Span4Mux_v I__9010 (
            .O(N__37100),
            .I(N__37004));
    Span4Mux_v I__9009 (
            .O(N__37095),
            .I(N__37004));
    Span4Mux_v I__9008 (
            .O(N__37090),
            .I(N__36997));
    Span4Mux_v I__9007 (
            .O(N__37085),
            .I(N__36997));
    LocalMux I__9006 (
            .O(N__37082),
            .I(N__36997));
    InMux I__9005 (
            .O(N__37079),
            .I(N__36991));
    InMux I__9004 (
            .O(N__37076),
            .I(N__36991));
    InMux I__9003 (
            .O(N__37073),
            .I(N__36984));
    InMux I__9002 (
            .O(N__37070),
            .I(N__36984));
    InMux I__9001 (
            .O(N__37067),
            .I(N__36984));
    InMux I__9000 (
            .O(N__37064),
            .I(N__36975));
    InMux I__8999 (
            .O(N__37063),
            .I(N__36975));
    InMux I__8998 (
            .O(N__37060),
            .I(N__36975));
    InMux I__8997 (
            .O(N__37057),
            .I(N__36975));
    InMux I__8996 (
            .O(N__37056),
            .I(N__36970));
    InMux I__8995 (
            .O(N__37053),
            .I(N__36970));
    Span4Mux_h I__8994 (
            .O(N__37050),
            .I(N__36967));
    Span4Mux_h I__8993 (
            .O(N__37047),
            .I(N__36960));
    Span4Mux_v I__8992 (
            .O(N__37044),
            .I(N__36960));
    Span4Mux_h I__8991 (
            .O(N__37039),
            .I(N__36960));
    InMux I__8990 (
            .O(N__37036),
            .I(N__36957));
    Span4Mux_v I__8989 (
            .O(N__37033),
            .I(N__36952));
    LocalMux I__8988 (
            .O(N__37030),
            .I(N__36952));
    SRMux I__8987 (
            .O(N__37029),
            .I(N__36949));
    Span4Mux_h I__8986 (
            .O(N__37026),
            .I(N__36942));
    Span4Mux_v I__8985 (
            .O(N__37019),
            .I(N__36942));
    LocalMux I__8984 (
            .O(N__37016),
            .I(N__36942));
    SRMux I__8983 (
            .O(N__37015),
            .I(N__36939));
    SRMux I__8982 (
            .O(N__37014),
            .I(N__36935));
    SRMux I__8981 (
            .O(N__37013),
            .I(N__36932));
    SRMux I__8980 (
            .O(N__37012),
            .I(N__36929));
    Span4Mux_v I__8979 (
            .O(N__37009),
            .I(N__36922));
    Span4Mux_h I__8978 (
            .O(N__37004),
            .I(N__36922));
    Span4Mux_h I__8977 (
            .O(N__36997),
            .I(N__36922));
    SRMux I__8976 (
            .O(N__36996),
            .I(N__36918));
    LocalMux I__8975 (
            .O(N__36991),
            .I(N__36915));
    LocalMux I__8974 (
            .O(N__36984),
            .I(N__36908));
    LocalMux I__8973 (
            .O(N__36975),
            .I(N__36908));
    LocalMux I__8972 (
            .O(N__36970),
            .I(N__36908));
    Span4Mux_h I__8971 (
            .O(N__36967),
            .I(N__36905));
    Span4Mux_h I__8970 (
            .O(N__36960),
            .I(N__36900));
    LocalMux I__8969 (
            .O(N__36957),
            .I(N__36900));
    Span4Mux_v I__8968 (
            .O(N__36952),
            .I(N__36891));
    LocalMux I__8967 (
            .O(N__36949),
            .I(N__36891));
    Span4Mux_h I__8966 (
            .O(N__36942),
            .I(N__36891));
    LocalMux I__8965 (
            .O(N__36939),
            .I(N__36891));
    SRMux I__8964 (
            .O(N__36938),
            .I(N__36888));
    LocalMux I__8963 (
            .O(N__36935),
            .I(N__36883));
    LocalMux I__8962 (
            .O(N__36932),
            .I(N__36883));
    LocalMux I__8961 (
            .O(N__36929),
            .I(N__36880));
    Span4Mux_h I__8960 (
            .O(N__36922),
            .I(N__36877));
    SRMux I__8959 (
            .O(N__36921),
            .I(N__36874));
    LocalMux I__8958 (
            .O(N__36918),
            .I(N__36871));
    Span12Mux_v I__8957 (
            .O(N__36915),
            .I(N__36868));
    Span12Mux_v I__8956 (
            .O(N__36908),
            .I(N__36865));
    Sp12to4 I__8955 (
            .O(N__36905),
            .I(N__36862));
    Span4Mux_v I__8954 (
            .O(N__36900),
            .I(N__36859));
    Span4Mux_v I__8953 (
            .O(N__36891),
            .I(N__36854));
    LocalMux I__8952 (
            .O(N__36888),
            .I(N__36854));
    Span4Mux_v I__8951 (
            .O(N__36883),
            .I(N__36851));
    Span4Mux_v I__8950 (
            .O(N__36880),
            .I(N__36848));
    Span4Mux_h I__8949 (
            .O(N__36877),
            .I(N__36844));
    LocalMux I__8948 (
            .O(N__36874),
            .I(N__36841));
    Span4Mux_h I__8947 (
            .O(N__36871),
            .I(N__36838));
    Span12Mux_h I__8946 (
            .O(N__36868),
            .I(N__36831));
    Span12Mux_h I__8945 (
            .O(N__36865),
            .I(N__36831));
    Span12Mux_s11_v I__8944 (
            .O(N__36862),
            .I(N__36826));
    Sp12to4 I__8943 (
            .O(N__36859),
            .I(N__36826));
    Span4Mux_v I__8942 (
            .O(N__36854),
            .I(N__36819));
    Span4Mux_v I__8941 (
            .O(N__36851),
            .I(N__36819));
    Span4Mux_h I__8940 (
            .O(N__36848),
            .I(N__36819));
    SRMux I__8939 (
            .O(N__36847),
            .I(N__36816));
    Span4Mux_h I__8938 (
            .O(N__36844),
            .I(N__36809));
    Span4Mux_h I__8937 (
            .O(N__36841),
            .I(N__36809));
    Span4Mux_v I__8936 (
            .O(N__36838),
            .I(N__36809));
    SRMux I__8935 (
            .O(N__36837),
            .I(N__36806));
    SRMux I__8934 (
            .O(N__36836),
            .I(N__36803));
    Odrv12 I__8933 (
            .O(N__36831),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__8932 (
            .O(N__36826),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__8931 (
            .O(N__36819),
            .I(CONSTANT_ONE_NET));
    LocalMux I__8930 (
            .O(N__36816),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__8929 (
            .O(N__36809),
            .I(CONSTANT_ONE_NET));
    LocalMux I__8928 (
            .O(N__36806),
            .I(CONSTANT_ONE_NET));
    LocalMux I__8927 (
            .O(N__36803),
            .I(CONSTANT_ONE_NET));
    InMux I__8926 (
            .O(N__36788),
            .I(N__36784));
    InMux I__8925 (
            .O(N__36787),
            .I(N__36781));
    LocalMux I__8924 (
            .O(N__36784),
            .I(N__36777));
    LocalMux I__8923 (
            .O(N__36781),
            .I(N__36773));
    InMux I__8922 (
            .O(N__36780),
            .I(N__36770));
    Span12Mux_h I__8921 (
            .O(N__36777),
            .I(N__36767));
    InMux I__8920 (
            .O(N__36776),
            .I(N__36764));
    Span4Mux_v I__8919 (
            .O(N__36773),
            .I(N__36759));
    LocalMux I__8918 (
            .O(N__36770),
            .I(N__36759));
    Odrv12 I__8917 (
            .O(N__36767),
            .I(\b2v_inst.dir_energiaZ0Z_10 ));
    LocalMux I__8916 (
            .O(N__36764),
            .I(\b2v_inst.dir_energiaZ0Z_10 ));
    Odrv4 I__8915 (
            .O(N__36759),
            .I(\b2v_inst.dir_energiaZ0Z_10 ));
    CascadeMux I__8914 (
            .O(N__36752),
            .I(N__36748));
    InMux I__8913 (
            .O(N__36751),
            .I(N__36742));
    InMux I__8912 (
            .O(N__36748),
            .I(N__36739));
    InMux I__8911 (
            .O(N__36747),
            .I(N__36735));
    CascadeMux I__8910 (
            .O(N__36746),
            .I(N__36732));
    InMux I__8909 (
            .O(N__36745),
            .I(N__36729));
    LocalMux I__8908 (
            .O(N__36742),
            .I(N__36723));
    LocalMux I__8907 (
            .O(N__36739),
            .I(N__36720));
    CascadeMux I__8906 (
            .O(N__36738),
            .I(N__36717));
    LocalMux I__8905 (
            .O(N__36735),
            .I(N__36714));
    InMux I__8904 (
            .O(N__36732),
            .I(N__36711));
    LocalMux I__8903 (
            .O(N__36729),
            .I(N__36707));
    InMux I__8902 (
            .O(N__36728),
            .I(N__36704));
    InMux I__8901 (
            .O(N__36727),
            .I(N__36701));
    CascadeMux I__8900 (
            .O(N__36726),
            .I(N__36698));
    Span4Mux_v I__8899 (
            .O(N__36723),
            .I(N__36692));
    Span4Mux_v I__8898 (
            .O(N__36720),
            .I(N__36692));
    InMux I__8897 (
            .O(N__36717),
            .I(N__36689));
    Span4Mux_v I__8896 (
            .O(N__36714),
            .I(N__36684));
    LocalMux I__8895 (
            .O(N__36711),
            .I(N__36684));
    InMux I__8894 (
            .O(N__36710),
            .I(N__36681));
    Span4Mux_v I__8893 (
            .O(N__36707),
            .I(N__36674));
    LocalMux I__8892 (
            .O(N__36704),
            .I(N__36674));
    LocalMux I__8891 (
            .O(N__36701),
            .I(N__36674));
    InMux I__8890 (
            .O(N__36698),
            .I(N__36671));
    InMux I__8889 (
            .O(N__36697),
            .I(N__36668));
    Sp12to4 I__8888 (
            .O(N__36692),
            .I(N__36665));
    LocalMux I__8887 (
            .O(N__36689),
            .I(N__36662));
    Sp12to4 I__8886 (
            .O(N__36684),
            .I(N__36657));
    LocalMux I__8885 (
            .O(N__36681),
            .I(N__36657));
    Span4Mux_h I__8884 (
            .O(N__36674),
            .I(N__36652));
    LocalMux I__8883 (
            .O(N__36671),
            .I(N__36652));
    LocalMux I__8882 (
            .O(N__36668),
            .I(N__36649));
    Span12Mux_h I__8881 (
            .O(N__36665),
            .I(N__36644));
    Sp12to4 I__8880 (
            .O(N__36662),
            .I(N__36644));
    Span12Mux_v I__8879 (
            .O(N__36657),
            .I(N__36641));
    Span4Mux_h I__8878 (
            .O(N__36652),
            .I(N__36638));
    Odrv4 I__8877 (
            .O(N__36649),
            .I(\b2v_inst.indiceZ0Z_10 ));
    Odrv12 I__8876 (
            .O(N__36644),
            .I(\b2v_inst.indiceZ0Z_10 ));
    Odrv12 I__8875 (
            .O(N__36641),
            .I(\b2v_inst.indiceZ0Z_10 ));
    Odrv4 I__8874 (
            .O(N__36638),
            .I(\b2v_inst.indiceZ0Z_10 ));
    CascadeMux I__8873 (
            .O(N__36629),
            .I(N__36626));
    CascadeBuf I__8872 (
            .O(N__36626),
            .I(N__36622));
    CascadeMux I__8871 (
            .O(N__36625),
            .I(N__36619));
    CascadeMux I__8870 (
            .O(N__36622),
            .I(N__36616));
    CascadeBuf I__8869 (
            .O(N__36619),
            .I(N__36613));
    CascadeBuf I__8868 (
            .O(N__36616),
            .I(N__36610));
    CascadeMux I__8867 (
            .O(N__36613),
            .I(N__36607));
    CascadeMux I__8866 (
            .O(N__36610),
            .I(N__36604));
    CascadeBuf I__8865 (
            .O(N__36607),
            .I(N__36601));
    InMux I__8864 (
            .O(N__36604),
            .I(N__36598));
    CascadeMux I__8863 (
            .O(N__36601),
            .I(N__36595));
    LocalMux I__8862 (
            .O(N__36598),
            .I(N__36592));
    InMux I__8861 (
            .O(N__36595),
            .I(N__36589));
    Span4Mux_h I__8860 (
            .O(N__36592),
            .I(N__36586));
    LocalMux I__8859 (
            .O(N__36589),
            .I(N_445_i));
    Odrv4 I__8858 (
            .O(N__36586),
            .I(N_445_i));
    InMux I__8857 (
            .O(N__36581),
            .I(N__36577));
    InMux I__8856 (
            .O(N__36580),
            .I(N__36574));
    LocalMux I__8855 (
            .O(N__36577),
            .I(N__36566));
    LocalMux I__8854 (
            .O(N__36574),
            .I(N__36562));
    InMux I__8853 (
            .O(N__36573),
            .I(N__36559));
    InMux I__8852 (
            .O(N__36572),
            .I(N__36556));
    InMux I__8851 (
            .O(N__36571),
            .I(N__36553));
    InMux I__8850 (
            .O(N__36570),
            .I(N__36550));
    InMux I__8849 (
            .O(N__36569),
            .I(N__36547));
    Sp12to4 I__8848 (
            .O(N__36566),
            .I(N__36544));
    InMux I__8847 (
            .O(N__36565),
            .I(N__36541));
    Span4Mux_v I__8846 (
            .O(N__36562),
            .I(N__36536));
    LocalMux I__8845 (
            .O(N__36559),
            .I(N__36536));
    LocalMux I__8844 (
            .O(N__36556),
            .I(N__36531));
    LocalMux I__8843 (
            .O(N__36553),
            .I(N__36531));
    LocalMux I__8842 (
            .O(N__36550),
            .I(N__36528));
    LocalMux I__8841 (
            .O(N__36547),
            .I(N__36524));
    Span12Mux_v I__8840 (
            .O(N__36544),
            .I(N__36520));
    LocalMux I__8839 (
            .O(N__36541),
            .I(N__36513));
    Span4Mux_v I__8838 (
            .O(N__36536),
            .I(N__36513));
    Span4Mux_h I__8837 (
            .O(N__36531),
            .I(N__36513));
    Span4Mux_h I__8836 (
            .O(N__36528),
            .I(N__36509));
    InMux I__8835 (
            .O(N__36527),
            .I(N__36506));
    Span4Mux_v I__8834 (
            .O(N__36524),
            .I(N__36503));
    InMux I__8833 (
            .O(N__36523),
            .I(N__36500));
    Span12Mux_h I__8832 (
            .O(N__36520),
            .I(N__36496));
    Span4Mux_h I__8831 (
            .O(N__36513),
            .I(N__36493));
    InMux I__8830 (
            .O(N__36512),
            .I(N__36490));
    Span4Mux_v I__8829 (
            .O(N__36509),
            .I(N__36481));
    LocalMux I__8828 (
            .O(N__36506),
            .I(N__36481));
    Span4Mux_h I__8827 (
            .O(N__36503),
            .I(N__36481));
    LocalMux I__8826 (
            .O(N__36500),
            .I(N__36481));
    InMux I__8825 (
            .O(N__36499),
            .I(N__36478));
    Odrv12 I__8824 (
            .O(N__36496),
            .I(\b2v_inst.indiceZ0Z_3 ));
    Odrv4 I__8823 (
            .O(N__36493),
            .I(\b2v_inst.indiceZ0Z_3 ));
    LocalMux I__8822 (
            .O(N__36490),
            .I(\b2v_inst.indiceZ0Z_3 ));
    Odrv4 I__8821 (
            .O(N__36481),
            .I(\b2v_inst.indiceZ0Z_3 ));
    LocalMux I__8820 (
            .O(N__36478),
            .I(\b2v_inst.indiceZ0Z_3 ));
    CascadeMux I__8819 (
            .O(N__36467),
            .I(N__36464));
    InMux I__8818 (
            .O(N__36464),
            .I(N__36460));
    InMux I__8817 (
            .O(N__36463),
            .I(N__36457));
    LocalMux I__8816 (
            .O(N__36460),
            .I(N__36454));
    LocalMux I__8815 (
            .O(N__36457),
            .I(N__36450));
    Span12Mux_v I__8814 (
            .O(N__36454),
            .I(N__36445));
    InMux I__8813 (
            .O(N__36453),
            .I(N__36442));
    Span4Mux_v I__8812 (
            .O(N__36450),
            .I(N__36439));
    InMux I__8811 (
            .O(N__36449),
            .I(N__36436));
    InMux I__8810 (
            .O(N__36448),
            .I(N__36433));
    Odrv12 I__8809 (
            .O(N__36445),
            .I(\b2v_inst.dir_energiaZ0Z_3 ));
    LocalMux I__8808 (
            .O(N__36442),
            .I(\b2v_inst.dir_energiaZ0Z_3 ));
    Odrv4 I__8807 (
            .O(N__36439),
            .I(\b2v_inst.dir_energiaZ0Z_3 ));
    LocalMux I__8806 (
            .O(N__36436),
            .I(\b2v_inst.dir_energiaZ0Z_3 ));
    LocalMux I__8805 (
            .O(N__36433),
            .I(\b2v_inst.dir_energiaZ0Z_3 ));
    CascadeMux I__8804 (
            .O(N__36422),
            .I(N__36418));
    CascadeMux I__8803 (
            .O(N__36421),
            .I(N__36415));
    CascadeBuf I__8802 (
            .O(N__36418),
            .I(N__36412));
    CascadeBuf I__8801 (
            .O(N__36415),
            .I(N__36409));
    CascadeMux I__8800 (
            .O(N__36412),
            .I(N__36406));
    CascadeMux I__8799 (
            .O(N__36409),
            .I(N__36403));
    CascadeBuf I__8798 (
            .O(N__36406),
            .I(N__36400));
    CascadeBuf I__8797 (
            .O(N__36403),
            .I(N__36397));
    CascadeMux I__8796 (
            .O(N__36400),
            .I(N__36394));
    CascadeMux I__8795 (
            .O(N__36397),
            .I(N__36391));
    InMux I__8794 (
            .O(N__36394),
            .I(N__36388));
    InMux I__8793 (
            .O(N__36391),
            .I(N__36385));
    LocalMux I__8792 (
            .O(N__36388),
            .I(N__36382));
    LocalMux I__8791 (
            .O(N__36385),
            .I(N_357_i));
    Odrv4 I__8790 (
            .O(N__36382),
            .I(N_357_i));
    InMux I__8789 (
            .O(N__36377),
            .I(N__36372));
    InMux I__8788 (
            .O(N__36376),
            .I(N__36369));
    CascadeMux I__8787 (
            .O(N__36375),
            .I(N__36364));
    LocalMux I__8786 (
            .O(N__36372),
            .I(N__36360));
    LocalMux I__8785 (
            .O(N__36369),
            .I(N__36354));
    InMux I__8784 (
            .O(N__36368),
            .I(N__36351));
    InMux I__8783 (
            .O(N__36367),
            .I(N__36348));
    InMux I__8782 (
            .O(N__36364),
            .I(N__36344));
    InMux I__8781 (
            .O(N__36363),
            .I(N__36341));
    Span4Mux_v I__8780 (
            .O(N__36360),
            .I(N__36338));
    InMux I__8779 (
            .O(N__36359),
            .I(N__36334));
    InMux I__8778 (
            .O(N__36358),
            .I(N__36331));
    InMux I__8777 (
            .O(N__36357),
            .I(N__36328));
    Sp12to4 I__8776 (
            .O(N__36354),
            .I(N__36325));
    LocalMux I__8775 (
            .O(N__36351),
            .I(N__36322));
    LocalMux I__8774 (
            .O(N__36348),
            .I(N__36319));
    InMux I__8773 (
            .O(N__36347),
            .I(N__36316));
    LocalMux I__8772 (
            .O(N__36344),
            .I(N__36313));
    LocalMux I__8771 (
            .O(N__36341),
            .I(N__36310));
    Span4Mux_v I__8770 (
            .O(N__36338),
            .I(N__36306));
    InMux I__8769 (
            .O(N__36337),
            .I(N__36303));
    LocalMux I__8768 (
            .O(N__36334),
            .I(N__36296));
    LocalMux I__8767 (
            .O(N__36331),
            .I(N__36296));
    LocalMux I__8766 (
            .O(N__36328),
            .I(N__36296));
    Span12Mux_v I__8765 (
            .O(N__36325),
            .I(N__36293));
    Span4Mux_v I__8764 (
            .O(N__36322),
            .I(N__36286));
    Span4Mux_v I__8763 (
            .O(N__36319),
            .I(N__36286));
    LocalMux I__8762 (
            .O(N__36316),
            .I(N__36286));
    Span4Mux_v I__8761 (
            .O(N__36313),
            .I(N__36283));
    Span4Mux_v I__8760 (
            .O(N__36310),
            .I(N__36280));
    InMux I__8759 (
            .O(N__36309),
            .I(N__36277));
    Span4Mux_v I__8758 (
            .O(N__36306),
            .I(N__36270));
    LocalMux I__8757 (
            .O(N__36303),
            .I(N__36270));
    Span4Mux_v I__8756 (
            .O(N__36296),
            .I(N__36270));
    Odrv12 I__8755 (
            .O(N__36293),
            .I(\b2v_inst.indiceZ0Z_4 ));
    Odrv4 I__8754 (
            .O(N__36286),
            .I(\b2v_inst.indiceZ0Z_4 ));
    Odrv4 I__8753 (
            .O(N__36283),
            .I(\b2v_inst.indiceZ0Z_4 ));
    Odrv4 I__8752 (
            .O(N__36280),
            .I(\b2v_inst.indiceZ0Z_4 ));
    LocalMux I__8751 (
            .O(N__36277),
            .I(\b2v_inst.indiceZ0Z_4 ));
    Odrv4 I__8750 (
            .O(N__36270),
            .I(\b2v_inst.indiceZ0Z_4 ));
    CascadeMux I__8749 (
            .O(N__36257),
            .I(N__36254));
    InMux I__8748 (
            .O(N__36254),
            .I(N__36251));
    LocalMux I__8747 (
            .O(N__36251),
            .I(N__36248));
    Span4Mux_v I__8746 (
            .O(N__36248),
            .I(N__36243));
    InMux I__8745 (
            .O(N__36247),
            .I(N__36240));
    InMux I__8744 (
            .O(N__36246),
            .I(N__36237));
    Span4Mux_h I__8743 (
            .O(N__36243),
            .I(N__36233));
    LocalMux I__8742 (
            .O(N__36240),
            .I(N__36230));
    LocalMux I__8741 (
            .O(N__36237),
            .I(N__36227));
    InMux I__8740 (
            .O(N__36236),
            .I(N__36224));
    Span4Mux_h I__8739 (
            .O(N__36233),
            .I(N__36219));
    Span4Mux_v I__8738 (
            .O(N__36230),
            .I(N__36219));
    Span4Mux_v I__8737 (
            .O(N__36227),
            .I(N__36214));
    LocalMux I__8736 (
            .O(N__36224),
            .I(N__36214));
    Odrv4 I__8735 (
            .O(N__36219),
            .I(\b2v_inst.dir_energiaZ0Z_4 ));
    Odrv4 I__8734 (
            .O(N__36214),
            .I(\b2v_inst.dir_energiaZ0Z_4 ));
    CascadeMux I__8733 (
            .O(N__36209),
            .I(N__36205));
    CascadeMux I__8732 (
            .O(N__36208),
            .I(N__36202));
    CascadeBuf I__8731 (
            .O(N__36205),
            .I(N__36199));
    CascadeBuf I__8730 (
            .O(N__36202),
            .I(N__36196));
    CascadeMux I__8729 (
            .O(N__36199),
            .I(N__36193));
    CascadeMux I__8728 (
            .O(N__36196),
            .I(N__36190));
    CascadeBuf I__8727 (
            .O(N__36193),
            .I(N__36187));
    CascadeBuf I__8726 (
            .O(N__36190),
            .I(N__36184));
    CascadeMux I__8725 (
            .O(N__36187),
            .I(N__36181));
    CascadeMux I__8724 (
            .O(N__36184),
            .I(N__36178));
    InMux I__8723 (
            .O(N__36181),
            .I(N__36175));
    InMux I__8722 (
            .O(N__36178),
            .I(N__36172));
    LocalMux I__8721 (
            .O(N__36175),
            .I(N__36169));
    LocalMux I__8720 (
            .O(N__36172),
            .I(N_356_i));
    Odrv4 I__8719 (
            .O(N__36169),
            .I(N_356_i));
    CascadeMux I__8718 (
            .O(N__36164),
            .I(N__36161));
    InMux I__8717 (
            .O(N__36161),
            .I(N__36158));
    LocalMux I__8716 (
            .O(N__36158),
            .I(N__36155));
    Span4Mux_v I__8715 (
            .O(N__36155),
            .I(N__36151));
    InMux I__8714 (
            .O(N__36154),
            .I(N__36148));
    Span4Mux_h I__8713 (
            .O(N__36151),
            .I(N__36143));
    LocalMux I__8712 (
            .O(N__36148),
            .I(N__36140));
    InMux I__8711 (
            .O(N__36147),
            .I(N__36137));
    InMux I__8710 (
            .O(N__36146),
            .I(N__36134));
    Span4Mux_h I__8709 (
            .O(N__36143),
            .I(N__36127));
    Span4Mux_v I__8708 (
            .O(N__36140),
            .I(N__36127));
    LocalMux I__8707 (
            .O(N__36137),
            .I(N__36127));
    LocalMux I__8706 (
            .O(N__36134),
            .I(\b2v_inst.dir_energiaZ0Z_2 ));
    Odrv4 I__8705 (
            .O(N__36127),
            .I(\b2v_inst.dir_energiaZ0Z_2 ));
    InMux I__8704 (
            .O(N__36122),
            .I(N__36118));
    InMux I__8703 (
            .O(N__36121),
            .I(N__36115));
    LocalMux I__8702 (
            .O(N__36118),
            .I(N__36110));
    LocalMux I__8701 (
            .O(N__36115),
            .I(N__36107));
    InMux I__8700 (
            .O(N__36114),
            .I(N__36104));
    CascadeMux I__8699 (
            .O(N__36113),
            .I(N__36100));
    Span4Mux_h I__8698 (
            .O(N__36110),
            .I(N__36097));
    Span4Mux_h I__8697 (
            .O(N__36107),
            .I(N__36093));
    LocalMux I__8696 (
            .O(N__36104),
            .I(N__36089));
    InMux I__8695 (
            .O(N__36103),
            .I(N__36086));
    InMux I__8694 (
            .O(N__36100),
            .I(N__36083));
    Span4Mux_h I__8693 (
            .O(N__36097),
            .I(N__36080));
    InMux I__8692 (
            .O(N__36096),
            .I(N__36077));
    Span4Mux_h I__8691 (
            .O(N__36093),
            .I(N__36073));
    InMux I__8690 (
            .O(N__36092),
            .I(N__36070));
    Span4Mux_v I__8689 (
            .O(N__36089),
            .I(N__36067));
    LocalMux I__8688 (
            .O(N__36086),
            .I(N__36064));
    LocalMux I__8687 (
            .O(N__36083),
            .I(N__36057));
    Span4Mux_v I__8686 (
            .O(N__36080),
            .I(N__36057));
    LocalMux I__8685 (
            .O(N__36077),
            .I(N__36057));
    CascadeMux I__8684 (
            .O(N__36076),
            .I(N__36054));
    Sp12to4 I__8683 (
            .O(N__36073),
            .I(N__36051));
    LocalMux I__8682 (
            .O(N__36070),
            .I(N__36045));
    Span4Mux_h I__8681 (
            .O(N__36067),
            .I(N__36045));
    Span4Mux_h I__8680 (
            .O(N__36064),
            .I(N__36040));
    Span4Mux_v I__8679 (
            .O(N__36057),
            .I(N__36037));
    InMux I__8678 (
            .O(N__36054),
            .I(N__36034));
    Span12Mux_v I__8677 (
            .O(N__36051),
            .I(N__36031));
    InMux I__8676 (
            .O(N__36050),
            .I(N__36028));
    Span4Mux_v I__8675 (
            .O(N__36045),
            .I(N__36025));
    InMux I__8674 (
            .O(N__36044),
            .I(N__36022));
    InMux I__8673 (
            .O(N__36043),
            .I(N__36019));
    Span4Mux_v I__8672 (
            .O(N__36040),
            .I(N__36012));
    Span4Mux_h I__8671 (
            .O(N__36037),
            .I(N__36012));
    LocalMux I__8670 (
            .O(N__36034),
            .I(N__36012));
    Odrv12 I__8669 (
            .O(N__36031),
            .I(\b2v_inst.indiceZ0Z_2 ));
    LocalMux I__8668 (
            .O(N__36028),
            .I(\b2v_inst.indiceZ0Z_2 ));
    Odrv4 I__8667 (
            .O(N__36025),
            .I(\b2v_inst.indiceZ0Z_2 ));
    LocalMux I__8666 (
            .O(N__36022),
            .I(\b2v_inst.indiceZ0Z_2 ));
    LocalMux I__8665 (
            .O(N__36019),
            .I(\b2v_inst.indiceZ0Z_2 ));
    Odrv4 I__8664 (
            .O(N__36012),
            .I(\b2v_inst.indiceZ0Z_2 ));
    CascadeMux I__8663 (
            .O(N__35999),
            .I(N__35995));
    CascadeMux I__8662 (
            .O(N__35998),
            .I(N__35992));
    CascadeBuf I__8661 (
            .O(N__35995),
            .I(N__35989));
    CascadeBuf I__8660 (
            .O(N__35992),
            .I(N__35986));
    CascadeMux I__8659 (
            .O(N__35989),
            .I(N__35983));
    CascadeMux I__8658 (
            .O(N__35986),
            .I(N__35980));
    CascadeBuf I__8657 (
            .O(N__35983),
            .I(N__35977));
    CascadeBuf I__8656 (
            .O(N__35980),
            .I(N__35974));
    CascadeMux I__8655 (
            .O(N__35977),
            .I(N__35971));
    CascadeMux I__8654 (
            .O(N__35974),
            .I(N__35968));
    InMux I__8653 (
            .O(N__35971),
            .I(N__35965));
    InMux I__8652 (
            .O(N__35968),
            .I(N__35962));
    LocalMux I__8651 (
            .O(N__35965),
            .I(N__35959));
    LocalMux I__8650 (
            .O(N__35962),
            .I(N_358_i));
    Odrv4 I__8649 (
            .O(N__35959),
            .I(N_358_i));
    CascadeMux I__8648 (
            .O(N__35954),
            .I(N__35949));
    InMux I__8647 (
            .O(N__35953),
            .I(N__35946));
    CascadeMux I__8646 (
            .O(N__35952),
            .I(N__35943));
    InMux I__8645 (
            .O(N__35949),
            .I(N__35940));
    LocalMux I__8644 (
            .O(N__35946),
            .I(N__35934));
    InMux I__8643 (
            .O(N__35943),
            .I(N__35930));
    LocalMux I__8642 (
            .O(N__35940),
            .I(N__35927));
    InMux I__8641 (
            .O(N__35939),
            .I(N__35924));
    InMux I__8640 (
            .O(N__35938),
            .I(N__35921));
    InMux I__8639 (
            .O(N__35937),
            .I(N__35916));
    Span4Mux_v I__8638 (
            .O(N__35934),
            .I(N__35912));
    InMux I__8637 (
            .O(N__35933),
            .I(N__35907));
    LocalMux I__8636 (
            .O(N__35930),
            .I(N__35904));
    Span4Mux_h I__8635 (
            .O(N__35927),
            .I(N__35897));
    LocalMux I__8634 (
            .O(N__35924),
            .I(N__35897));
    LocalMux I__8633 (
            .O(N__35921),
            .I(N__35897));
    InMux I__8632 (
            .O(N__35920),
            .I(N__35892));
    InMux I__8631 (
            .O(N__35919),
            .I(N__35892));
    LocalMux I__8630 (
            .O(N__35916),
            .I(N__35889));
    InMux I__8629 (
            .O(N__35915),
            .I(N__35886));
    Span4Mux_h I__8628 (
            .O(N__35912),
            .I(N__35883));
    InMux I__8627 (
            .O(N__35911),
            .I(N__35880));
    InMux I__8626 (
            .O(N__35910),
            .I(N__35877));
    LocalMux I__8625 (
            .O(N__35907),
            .I(N__35874));
    Span4Mux_h I__8624 (
            .O(N__35904),
            .I(N__35871));
    Span4Mux_v I__8623 (
            .O(N__35897),
            .I(N__35866));
    LocalMux I__8622 (
            .O(N__35892),
            .I(N__35866));
    Span4Mux_v I__8621 (
            .O(N__35889),
            .I(N__35863));
    LocalMux I__8620 (
            .O(N__35886),
            .I(N__35860));
    Span4Mux_h I__8619 (
            .O(N__35883),
            .I(N__35857));
    LocalMux I__8618 (
            .O(N__35880),
            .I(N__35854));
    LocalMux I__8617 (
            .O(N__35877),
            .I(N__35847));
    Span12Mux_h I__8616 (
            .O(N__35874),
            .I(N__35847));
    Sp12to4 I__8615 (
            .O(N__35871),
            .I(N__35847));
    Span4Mux_h I__8614 (
            .O(N__35866),
            .I(N__35844));
    Odrv4 I__8613 (
            .O(N__35863),
            .I(\b2v_inst.indiceZ0Z_9 ));
    Odrv12 I__8612 (
            .O(N__35860),
            .I(\b2v_inst.indiceZ0Z_9 ));
    Odrv4 I__8611 (
            .O(N__35857),
            .I(\b2v_inst.indiceZ0Z_9 ));
    Odrv4 I__8610 (
            .O(N__35854),
            .I(\b2v_inst.indiceZ0Z_9 ));
    Odrv12 I__8609 (
            .O(N__35847),
            .I(\b2v_inst.indiceZ0Z_9 ));
    Odrv4 I__8608 (
            .O(N__35844),
            .I(\b2v_inst.indiceZ0Z_9 ));
    CascadeMux I__8607 (
            .O(N__35831),
            .I(N__35828));
    InMux I__8606 (
            .O(N__35828),
            .I(N__35824));
    CascadeMux I__8605 (
            .O(N__35827),
            .I(N__35820));
    LocalMux I__8604 (
            .O(N__35824),
            .I(N__35816));
    InMux I__8603 (
            .O(N__35823),
            .I(N__35813));
    InMux I__8602 (
            .O(N__35820),
            .I(N__35809));
    InMux I__8601 (
            .O(N__35819),
            .I(N__35806));
    Span4Mux_v I__8600 (
            .O(N__35816),
            .I(N__35803));
    LocalMux I__8599 (
            .O(N__35813),
            .I(N__35800));
    CascadeMux I__8598 (
            .O(N__35812),
            .I(N__35797));
    LocalMux I__8597 (
            .O(N__35809),
            .I(N__35792));
    LocalMux I__8596 (
            .O(N__35806),
            .I(N__35792));
    Sp12to4 I__8595 (
            .O(N__35803),
            .I(N__35789));
    Span4Mux_h I__8594 (
            .O(N__35800),
            .I(N__35786));
    InMux I__8593 (
            .O(N__35797),
            .I(N__35783));
    Span4Mux_h I__8592 (
            .O(N__35792),
            .I(N__35780));
    Odrv12 I__8591 (
            .O(N__35789),
            .I(\b2v_inst.dir_energiaZ0Z_9 ));
    Odrv4 I__8590 (
            .O(N__35786),
            .I(\b2v_inst.dir_energiaZ0Z_9 ));
    LocalMux I__8589 (
            .O(N__35783),
            .I(\b2v_inst.dir_energiaZ0Z_9 ));
    Odrv4 I__8588 (
            .O(N__35780),
            .I(\b2v_inst.dir_energiaZ0Z_9 ));
    CascadeMux I__8587 (
            .O(N__35771),
            .I(N__35767));
    CascadeMux I__8586 (
            .O(N__35770),
            .I(N__35764));
    CascadeBuf I__8585 (
            .O(N__35767),
            .I(N__35761));
    CascadeBuf I__8584 (
            .O(N__35764),
            .I(N__35758));
    CascadeMux I__8583 (
            .O(N__35761),
            .I(N__35755));
    CascadeMux I__8582 (
            .O(N__35758),
            .I(N__35752));
    CascadeBuf I__8581 (
            .O(N__35755),
            .I(N__35749));
    CascadeBuf I__8580 (
            .O(N__35752),
            .I(N__35746));
    CascadeMux I__8579 (
            .O(N__35749),
            .I(N__35743));
    CascadeMux I__8578 (
            .O(N__35746),
            .I(N__35740));
    InMux I__8577 (
            .O(N__35743),
            .I(N__35737));
    InMux I__8576 (
            .O(N__35740),
            .I(N__35734));
    LocalMux I__8575 (
            .O(N__35737),
            .I(N__35731));
    LocalMux I__8574 (
            .O(N__35734),
            .I(N_444_i));
    Odrv4 I__8573 (
            .O(N__35731),
            .I(N_444_i));
    InMux I__8572 (
            .O(N__35726),
            .I(N__35723));
    LocalMux I__8571 (
            .O(N__35723),
            .I(N__35719));
    InMux I__8570 (
            .O(N__35722),
            .I(N__35716));
    Span4Mux_h I__8569 (
            .O(N__35719),
            .I(N__35712));
    LocalMux I__8568 (
            .O(N__35716),
            .I(N__35707));
    CascadeMux I__8567 (
            .O(N__35715),
            .I(N__35702));
    Span4Mux_h I__8566 (
            .O(N__35712),
            .I(N__35697));
    InMux I__8565 (
            .O(N__35711),
            .I(N__35694));
    InMux I__8564 (
            .O(N__35710),
            .I(N__35691));
    Span4Mux_v I__8563 (
            .O(N__35707),
            .I(N__35687));
    InMux I__8562 (
            .O(N__35706),
            .I(N__35684));
    InMux I__8561 (
            .O(N__35705),
            .I(N__35679));
    InMux I__8560 (
            .O(N__35702),
            .I(N__35676));
    InMux I__8559 (
            .O(N__35701),
            .I(N__35673));
    InMux I__8558 (
            .O(N__35700),
            .I(N__35670));
    Span4Mux_v I__8557 (
            .O(N__35697),
            .I(N__35664));
    LocalMux I__8556 (
            .O(N__35694),
            .I(N__35664));
    LocalMux I__8555 (
            .O(N__35691),
            .I(N__35661));
    InMux I__8554 (
            .O(N__35690),
            .I(N__35658));
    Sp12to4 I__8553 (
            .O(N__35687),
            .I(N__35655));
    LocalMux I__8552 (
            .O(N__35684),
            .I(N__35652));
    InMux I__8551 (
            .O(N__35683),
            .I(N__35649));
    InMux I__8550 (
            .O(N__35682),
            .I(N__35646));
    LocalMux I__8549 (
            .O(N__35679),
            .I(N__35641));
    LocalMux I__8548 (
            .O(N__35676),
            .I(N__35641));
    LocalMux I__8547 (
            .O(N__35673),
            .I(N__35636));
    LocalMux I__8546 (
            .O(N__35670),
            .I(N__35636));
    InMux I__8545 (
            .O(N__35669),
            .I(N__35633));
    Span4Mux_h I__8544 (
            .O(N__35664),
            .I(N__35626));
    Span4Mux_h I__8543 (
            .O(N__35661),
            .I(N__35626));
    LocalMux I__8542 (
            .O(N__35658),
            .I(N__35626));
    Span12Mux_h I__8541 (
            .O(N__35655),
            .I(N__35621));
    Sp12to4 I__8540 (
            .O(N__35652),
            .I(N__35621));
    LocalMux I__8539 (
            .O(N__35649),
            .I(N__35618));
    LocalMux I__8538 (
            .O(N__35646),
            .I(N__35615));
    Span4Mux_v I__8537 (
            .O(N__35641),
            .I(N__35608));
    Span4Mux_h I__8536 (
            .O(N__35636),
            .I(N__35608));
    LocalMux I__8535 (
            .O(N__35633),
            .I(N__35608));
    Span4Mux_h I__8534 (
            .O(N__35626),
            .I(N__35605));
    Odrv12 I__8533 (
            .O(N__35621),
            .I(\b2v_inst.indiceZ0Z_5 ));
    Odrv4 I__8532 (
            .O(N__35618),
            .I(\b2v_inst.indiceZ0Z_5 ));
    Odrv4 I__8531 (
            .O(N__35615),
            .I(\b2v_inst.indiceZ0Z_5 ));
    Odrv4 I__8530 (
            .O(N__35608),
            .I(\b2v_inst.indiceZ0Z_5 ));
    Odrv4 I__8529 (
            .O(N__35605),
            .I(\b2v_inst.indiceZ0Z_5 ));
    CascadeMux I__8528 (
            .O(N__35594),
            .I(N__35591));
    InMux I__8527 (
            .O(N__35591),
            .I(N__35588));
    LocalMux I__8526 (
            .O(N__35588),
            .I(N__35585));
    Span4Mux_h I__8525 (
            .O(N__35585),
            .I(N__35581));
    InMux I__8524 (
            .O(N__35584),
            .I(N__35578));
    Span4Mux_h I__8523 (
            .O(N__35581),
            .I(N__35572));
    LocalMux I__8522 (
            .O(N__35578),
            .I(N__35572));
    InMux I__8521 (
            .O(N__35577),
            .I(N__35567));
    Span4Mux_h I__8520 (
            .O(N__35572),
            .I(N__35564));
    InMux I__8519 (
            .O(N__35571),
            .I(N__35561));
    InMux I__8518 (
            .O(N__35570),
            .I(N__35558));
    LocalMux I__8517 (
            .O(N__35567),
            .I(\b2v_inst.dir_energiaZ0Z_5 ));
    Odrv4 I__8516 (
            .O(N__35564),
            .I(\b2v_inst.dir_energiaZ0Z_5 ));
    LocalMux I__8515 (
            .O(N__35561),
            .I(\b2v_inst.dir_energiaZ0Z_5 ));
    LocalMux I__8514 (
            .O(N__35558),
            .I(\b2v_inst.dir_energiaZ0Z_5 ));
    CascadeMux I__8513 (
            .O(N__35549),
            .I(N__35545));
    CascadeMux I__8512 (
            .O(N__35548),
            .I(N__35542));
    CascadeBuf I__8511 (
            .O(N__35545),
            .I(N__35539));
    CascadeBuf I__8510 (
            .O(N__35542),
            .I(N__35536));
    CascadeMux I__8509 (
            .O(N__35539),
            .I(N__35533));
    CascadeMux I__8508 (
            .O(N__35536),
            .I(N__35530));
    CascadeBuf I__8507 (
            .O(N__35533),
            .I(N__35527));
    CascadeBuf I__8506 (
            .O(N__35530),
            .I(N__35524));
    CascadeMux I__8505 (
            .O(N__35527),
            .I(N__35521));
    CascadeMux I__8504 (
            .O(N__35524),
            .I(N__35518));
    InMux I__8503 (
            .O(N__35521),
            .I(N__35515));
    InMux I__8502 (
            .O(N__35518),
            .I(N__35512));
    LocalMux I__8501 (
            .O(N__35515),
            .I(N__35509));
    LocalMux I__8500 (
            .O(N__35512),
            .I(N_355_i));
    Odrv4 I__8499 (
            .O(N__35509),
            .I(N_355_i));
    InMux I__8498 (
            .O(N__35504),
            .I(N__35501));
    LocalMux I__8497 (
            .O(N__35501),
            .I(N__35497));
    InMux I__8496 (
            .O(N__35500),
            .I(N__35494));
    Span4Mux_h I__8495 (
            .O(N__35497),
            .I(N__35488));
    LocalMux I__8494 (
            .O(N__35494),
            .I(N__35488));
    InMux I__8493 (
            .O(N__35493),
            .I(N__35485));
    Span4Mux_v I__8492 (
            .O(N__35488),
            .I(N__35479));
    LocalMux I__8491 (
            .O(N__35485),
            .I(N__35479));
    InMux I__8490 (
            .O(N__35484),
            .I(N__35476));
    Span4Mux_h I__8489 (
            .O(N__35479),
            .I(N__35473));
    LocalMux I__8488 (
            .O(N__35476),
            .I(N__35470));
    Span4Mux_h I__8487 (
            .O(N__35473),
            .I(N__35467));
    Odrv12 I__8486 (
            .O(N__35470),
            .I(b2v_inst_data_a_escribir_7));
    Odrv4 I__8485 (
            .O(N__35467),
            .I(b2v_inst_data_a_escribir_7));
    InMux I__8484 (
            .O(N__35462),
            .I(N__35459));
    LocalMux I__8483 (
            .O(N__35459),
            .I(N__35456));
    Span4Mux_v I__8482 (
            .O(N__35456),
            .I(N__35453));
    Odrv4 I__8481 (
            .O(N__35453),
            .I(N_113_i));
    InMux I__8480 (
            .O(N__35450),
            .I(N__35447));
    LocalMux I__8479 (
            .O(N__35447),
            .I(N__35444));
    Span4Mux_h I__8478 (
            .O(N__35444),
            .I(N__35441));
    Span4Mux_v I__8477 (
            .O(N__35441),
            .I(N__35438));
    Span4Mux_h I__8476 (
            .O(N__35438),
            .I(N__35435));
    Odrv4 I__8475 (
            .O(N__35435),
            .I(\b2v_inst.addr_ram_iv_i_0_0_1 ));
    CascadeMux I__8474 (
            .O(N__35432),
            .I(N__35429));
    InMux I__8473 (
            .O(N__35429),
            .I(N__35426));
    LocalMux I__8472 (
            .O(N__35426),
            .I(N__35423));
    Span4Mux_h I__8471 (
            .O(N__35423),
            .I(N__35420));
    Span4Mux_h I__8470 (
            .O(N__35420),
            .I(N__35417));
    Span4Mux_v I__8469 (
            .O(N__35417),
            .I(N__35414));
    Odrv4 I__8468 (
            .O(N__35414),
            .I(\b2v_inst.addr_ram_iv_i_0_1_1 ));
    CascadeMux I__8467 (
            .O(N__35411),
            .I(N__35407));
    CascadeMux I__8466 (
            .O(N__35410),
            .I(N__35404));
    CascadeBuf I__8465 (
            .O(N__35407),
            .I(N__35401));
    CascadeBuf I__8464 (
            .O(N__35404),
            .I(N__35398));
    CascadeMux I__8463 (
            .O(N__35401),
            .I(N__35395));
    CascadeMux I__8462 (
            .O(N__35398),
            .I(N__35392));
    CascadeBuf I__8461 (
            .O(N__35395),
            .I(N__35389));
    CascadeBuf I__8460 (
            .O(N__35392),
            .I(N__35386));
    CascadeMux I__8459 (
            .O(N__35389),
            .I(N__35383));
    CascadeMux I__8458 (
            .O(N__35386),
            .I(N__35380));
    CascadeBuf I__8457 (
            .O(N__35383),
            .I(N__35377));
    CascadeBuf I__8456 (
            .O(N__35380),
            .I(N__35374));
    CascadeMux I__8455 (
            .O(N__35377),
            .I(N__35371));
    CascadeMux I__8454 (
            .O(N__35374),
            .I(N__35368));
    CascadeBuf I__8453 (
            .O(N__35371),
            .I(N__35365));
    CascadeBuf I__8452 (
            .O(N__35368),
            .I(N__35362));
    CascadeMux I__8451 (
            .O(N__35365),
            .I(N__35359));
    CascadeMux I__8450 (
            .O(N__35362),
            .I(N__35356));
    CascadeBuf I__8449 (
            .O(N__35359),
            .I(N__35353));
    CascadeBuf I__8448 (
            .O(N__35356),
            .I(N__35350));
    CascadeMux I__8447 (
            .O(N__35353),
            .I(N__35347));
    CascadeMux I__8446 (
            .O(N__35350),
            .I(N__35344));
    InMux I__8445 (
            .O(N__35347),
            .I(N__35341));
    InMux I__8444 (
            .O(N__35344),
            .I(N__35338));
    LocalMux I__8443 (
            .O(N__35341),
            .I(N__35335));
    LocalMux I__8442 (
            .O(N__35338),
            .I(indice_RNI8K233_1));
    Odrv4 I__8441 (
            .O(N__35335),
            .I(indice_RNI8K233_1));
    CascadeMux I__8440 (
            .O(N__35330),
            .I(N__35327));
    InMux I__8439 (
            .O(N__35327),
            .I(N__35323));
    InMux I__8438 (
            .O(N__35326),
            .I(N__35319));
    LocalMux I__8437 (
            .O(N__35323),
            .I(N__35316));
    CascadeMux I__8436 (
            .O(N__35322),
            .I(N__35312));
    LocalMux I__8435 (
            .O(N__35319),
            .I(N__35309));
    Span4Mux_v I__8434 (
            .O(N__35316),
            .I(N__35306));
    InMux I__8433 (
            .O(N__35315),
            .I(N__35303));
    InMux I__8432 (
            .O(N__35312),
            .I(N__35300));
    Span4Mux_h I__8431 (
            .O(N__35309),
            .I(N__35297));
    Span4Mux_h I__8430 (
            .O(N__35306),
            .I(N__35294));
    LocalMux I__8429 (
            .O(N__35303),
            .I(N__35291));
    LocalMux I__8428 (
            .O(N__35300),
            .I(N__35288));
    Span4Mux_h I__8427 (
            .O(N__35297),
            .I(N__35285));
    Span4Mux_h I__8426 (
            .O(N__35294),
            .I(N__35280));
    Span4Mux_h I__8425 (
            .O(N__35291),
            .I(N__35280));
    Span12Mux_v I__8424 (
            .O(N__35288),
            .I(N__35277));
    Odrv4 I__8423 (
            .O(N__35285),
            .I(b2v_inst_data_a_escribir_6));
    Odrv4 I__8422 (
            .O(N__35280),
            .I(b2v_inst_data_a_escribir_6));
    Odrv12 I__8421 (
            .O(N__35277),
            .I(b2v_inst_data_a_escribir_6));
    InMux I__8420 (
            .O(N__35270),
            .I(N__35267));
    LocalMux I__8419 (
            .O(N__35267),
            .I(N__35264));
    Span4Mux_v I__8418 (
            .O(N__35264),
            .I(N__35261));
    Odrv4 I__8417 (
            .O(N__35261),
            .I(N_114_i));
    InMux I__8416 (
            .O(N__35258),
            .I(N__35255));
    LocalMux I__8415 (
            .O(N__35255),
            .I(N__35252));
    Span4Mux_v I__8414 (
            .O(N__35252),
            .I(N__35249));
    Span4Mux_h I__8413 (
            .O(N__35249),
            .I(N__35246));
    Odrv4 I__8412 (
            .O(N__35246),
            .I(\b2v_inst.addr_ram_iv_i_0_2 ));
    InMux I__8411 (
            .O(N__35243),
            .I(N__35228));
    InMux I__8410 (
            .O(N__35242),
            .I(N__35228));
    InMux I__8409 (
            .O(N__35241),
            .I(N__35228));
    InMux I__8408 (
            .O(N__35240),
            .I(N__35228));
    InMux I__8407 (
            .O(N__35239),
            .I(N__35223));
    InMux I__8406 (
            .O(N__35238),
            .I(N__35223));
    InMux I__8405 (
            .O(N__35237),
            .I(N__35220));
    LocalMux I__8404 (
            .O(N__35228),
            .I(N__35210));
    LocalMux I__8403 (
            .O(N__35223),
            .I(N__35210));
    LocalMux I__8402 (
            .O(N__35220),
            .I(N__35204));
    InMux I__8401 (
            .O(N__35219),
            .I(N__35197));
    InMux I__8400 (
            .O(N__35218),
            .I(N__35197));
    InMux I__8399 (
            .O(N__35217),
            .I(N__35197));
    InMux I__8398 (
            .O(N__35216),
            .I(N__35193));
    InMux I__8397 (
            .O(N__35215),
            .I(N__35190));
    Span4Mux_v I__8396 (
            .O(N__35210),
            .I(N__35182));
    InMux I__8395 (
            .O(N__35209),
            .I(N__35179));
    InMux I__8394 (
            .O(N__35208),
            .I(N__35176));
    InMux I__8393 (
            .O(N__35207),
            .I(N__35173));
    Span4Mux_v I__8392 (
            .O(N__35204),
            .I(N__35167));
    LocalMux I__8391 (
            .O(N__35197),
            .I(N__35167));
    InMux I__8390 (
            .O(N__35196),
            .I(N__35163));
    LocalMux I__8389 (
            .O(N__35193),
            .I(N__35160));
    LocalMux I__8388 (
            .O(N__35190),
            .I(N__35157));
    InMux I__8387 (
            .O(N__35189),
            .I(N__35148));
    InMux I__8386 (
            .O(N__35188),
            .I(N__35148));
    InMux I__8385 (
            .O(N__35187),
            .I(N__35148));
    InMux I__8384 (
            .O(N__35186),
            .I(N__35148));
    InMux I__8383 (
            .O(N__35185),
            .I(N__35145));
    Sp12to4 I__8382 (
            .O(N__35182),
            .I(N__35140));
    LocalMux I__8381 (
            .O(N__35179),
            .I(N__35140));
    LocalMux I__8380 (
            .O(N__35176),
            .I(N__35137));
    LocalMux I__8379 (
            .O(N__35173),
            .I(N__35134));
    InMux I__8378 (
            .O(N__35172),
            .I(N__35131));
    Span4Mux_v I__8377 (
            .O(N__35167),
            .I(N__35128));
    InMux I__8376 (
            .O(N__35166),
            .I(N__35125));
    LocalMux I__8375 (
            .O(N__35163),
            .I(N__35122));
    Span4Mux_v I__8374 (
            .O(N__35160),
            .I(N__35119));
    Span4Mux_v I__8373 (
            .O(N__35157),
            .I(N__35116));
    LocalMux I__8372 (
            .O(N__35148),
            .I(N__35113));
    LocalMux I__8371 (
            .O(N__35145),
            .I(N__35108));
    Span12Mux_h I__8370 (
            .O(N__35140),
            .I(N__35108));
    Span12Mux_h I__8369 (
            .O(N__35137),
            .I(N__35105));
    Span4Mux_v I__8368 (
            .O(N__35134),
            .I(N__35100));
    LocalMux I__8367 (
            .O(N__35131),
            .I(N__35100));
    Span4Mux_h I__8366 (
            .O(N__35128),
            .I(N__35095));
    LocalMux I__8365 (
            .O(N__35125),
            .I(N__35095));
    Span12Mux_h I__8364 (
            .O(N__35122),
            .I(N__35092));
    Odrv4 I__8363 (
            .O(N__35119),
            .I(\b2v_inst.N_480 ));
    Odrv4 I__8362 (
            .O(N__35116),
            .I(\b2v_inst.N_480 ));
    Odrv4 I__8361 (
            .O(N__35113),
            .I(\b2v_inst.N_480 ));
    Odrv12 I__8360 (
            .O(N__35108),
            .I(\b2v_inst.N_480 ));
    Odrv12 I__8359 (
            .O(N__35105),
            .I(\b2v_inst.N_480 ));
    Odrv4 I__8358 (
            .O(N__35100),
            .I(\b2v_inst.N_480 ));
    Odrv4 I__8357 (
            .O(N__35095),
            .I(\b2v_inst.N_480 ));
    Odrv12 I__8356 (
            .O(N__35092),
            .I(\b2v_inst.N_480 ));
    CascadeMux I__8355 (
            .O(N__35075),
            .I(N__35072));
    InMux I__8354 (
            .O(N__35072),
            .I(N__35069));
    LocalMux I__8353 (
            .O(N__35069),
            .I(N__35066));
    Span4Mux_v I__8352 (
            .O(N__35066),
            .I(N__35063));
    Span4Mux_h I__8351 (
            .O(N__35063),
            .I(N__35060));
    Odrv4 I__8350 (
            .O(N__35060),
            .I(\b2v_inst.addr_ram_iv_i_1_2 ));
    CascadeMux I__8349 (
            .O(N__35057),
            .I(N__35053));
    CascadeMux I__8348 (
            .O(N__35056),
            .I(N__35050));
    CascadeBuf I__8347 (
            .O(N__35053),
            .I(N__35047));
    CascadeBuf I__8346 (
            .O(N__35050),
            .I(N__35044));
    CascadeMux I__8345 (
            .O(N__35047),
            .I(N__35041));
    CascadeMux I__8344 (
            .O(N__35044),
            .I(N__35038));
    CascadeBuf I__8343 (
            .O(N__35041),
            .I(N__35035));
    CascadeBuf I__8342 (
            .O(N__35038),
            .I(N__35032));
    CascadeMux I__8341 (
            .O(N__35035),
            .I(N__35029));
    CascadeMux I__8340 (
            .O(N__35032),
            .I(N__35026));
    CascadeBuf I__8339 (
            .O(N__35029),
            .I(N__35023));
    CascadeBuf I__8338 (
            .O(N__35026),
            .I(N__35020));
    CascadeMux I__8337 (
            .O(N__35023),
            .I(N__35017));
    CascadeMux I__8336 (
            .O(N__35020),
            .I(N__35014));
    CascadeBuf I__8335 (
            .O(N__35017),
            .I(N__35011));
    CascadeBuf I__8334 (
            .O(N__35014),
            .I(N__35008));
    CascadeMux I__8333 (
            .O(N__35011),
            .I(N__35005));
    CascadeMux I__8332 (
            .O(N__35008),
            .I(N__35002));
    CascadeBuf I__8331 (
            .O(N__35005),
            .I(N__34999));
    CascadeBuf I__8330 (
            .O(N__35002),
            .I(N__34996));
    CascadeMux I__8329 (
            .O(N__34999),
            .I(N__34993));
    CascadeMux I__8328 (
            .O(N__34996),
            .I(N__34990));
    InMux I__8327 (
            .O(N__34993),
            .I(N__34987));
    InMux I__8326 (
            .O(N__34990),
            .I(N__34984));
    LocalMux I__8325 (
            .O(N__34987),
            .I(N__34979));
    LocalMux I__8324 (
            .O(N__34984),
            .I(N__34979));
    Odrv4 I__8323 (
            .O(N__34979),
            .I(indice_RNIDP233_2));
    InMux I__8322 (
            .O(N__34976),
            .I(N__34970));
    InMux I__8321 (
            .O(N__34975),
            .I(N__34967));
    InMux I__8320 (
            .O(N__34974),
            .I(N__34963));
    InMux I__8319 (
            .O(N__34973),
            .I(N__34960));
    LocalMux I__8318 (
            .O(N__34970),
            .I(N__34957));
    LocalMux I__8317 (
            .O(N__34967),
            .I(N__34954));
    CascadeMux I__8316 (
            .O(N__34966),
            .I(N__34951));
    LocalMux I__8315 (
            .O(N__34963),
            .I(N__34948));
    LocalMux I__8314 (
            .O(N__34960),
            .I(N__34945));
    Span4Mux_h I__8313 (
            .O(N__34957),
            .I(N__34942));
    Span4Mux_v I__8312 (
            .O(N__34954),
            .I(N__34939));
    InMux I__8311 (
            .O(N__34951),
            .I(N__34936));
    Span4Mux_v I__8310 (
            .O(N__34948),
            .I(N__34931));
    Span4Mux_v I__8309 (
            .O(N__34945),
            .I(N__34931));
    Span4Mux_v I__8308 (
            .O(N__34942),
            .I(N__34928));
    Sp12to4 I__8307 (
            .O(N__34939),
            .I(N__34921));
    LocalMux I__8306 (
            .O(N__34936),
            .I(N__34921));
    Sp12to4 I__8305 (
            .O(N__34931),
            .I(N__34921));
    Odrv4 I__8304 (
            .O(N__34928),
            .I(b2v_inst_data_a_escribir_0));
    Odrv12 I__8303 (
            .O(N__34921),
            .I(b2v_inst_data_a_escribir_0));
    InMux I__8302 (
            .O(N__34916),
            .I(N__34913));
    LocalMux I__8301 (
            .O(N__34913),
            .I(N_557_i));
    InMux I__8300 (
            .O(N__34910),
            .I(N__34904));
    CascadeMux I__8299 (
            .O(N__34909),
            .I(N__34900));
    InMux I__8298 (
            .O(N__34908),
            .I(N__34897));
    InMux I__8297 (
            .O(N__34907),
            .I(N__34894));
    LocalMux I__8296 (
            .O(N__34904),
            .I(N__34891));
    InMux I__8295 (
            .O(N__34903),
            .I(N__34888));
    InMux I__8294 (
            .O(N__34900),
            .I(N__34885));
    LocalMux I__8293 (
            .O(N__34897),
            .I(b2v_inst_cantidad_temp_0));
    LocalMux I__8292 (
            .O(N__34894),
            .I(b2v_inst_cantidad_temp_0));
    Odrv12 I__8291 (
            .O(N__34891),
            .I(b2v_inst_cantidad_temp_0));
    LocalMux I__8290 (
            .O(N__34888),
            .I(b2v_inst_cantidad_temp_0));
    LocalMux I__8289 (
            .O(N__34885),
            .I(b2v_inst_cantidad_temp_0));
    InMux I__8288 (
            .O(N__34874),
            .I(N__34871));
    LocalMux I__8287 (
            .O(N__34871),
            .I(N__34867));
    InMux I__8286 (
            .O(N__34870),
            .I(N__34862));
    Span4Mux_h I__8285 (
            .O(N__34867),
            .I(N__34859));
    InMux I__8284 (
            .O(N__34866),
            .I(N__34856));
    InMux I__8283 (
            .O(N__34865),
            .I(N__34853));
    LocalMux I__8282 (
            .O(N__34862),
            .I(b2v_inst_cantidad_temp_1));
    Odrv4 I__8281 (
            .O(N__34859),
            .I(b2v_inst_cantidad_temp_1));
    LocalMux I__8280 (
            .O(N__34856),
            .I(b2v_inst_cantidad_temp_1));
    LocalMux I__8279 (
            .O(N__34853),
            .I(b2v_inst_cantidad_temp_1));
    CascadeMux I__8278 (
            .O(N__34844),
            .I(N__34841));
    InMux I__8277 (
            .O(N__34841),
            .I(N__34835));
    InMux I__8276 (
            .O(N__34840),
            .I(N__34832));
    CascadeMux I__8275 (
            .O(N__34839),
            .I(N__34829));
    InMux I__8274 (
            .O(N__34838),
            .I(N__34826));
    LocalMux I__8273 (
            .O(N__34835),
            .I(N__34822));
    LocalMux I__8272 (
            .O(N__34832),
            .I(N__34819));
    InMux I__8271 (
            .O(N__34829),
            .I(N__34816));
    LocalMux I__8270 (
            .O(N__34826),
            .I(N__34813));
    InMux I__8269 (
            .O(N__34825),
            .I(N__34810));
    Span4Mux_h I__8268 (
            .O(N__34822),
            .I(N__34807));
    Span4Mux_v I__8267 (
            .O(N__34819),
            .I(N__34804));
    LocalMux I__8266 (
            .O(N__34816),
            .I(N__34801));
    Span4Mux_v I__8265 (
            .O(N__34813),
            .I(N__34798));
    LocalMux I__8264 (
            .O(N__34810),
            .I(N__34795));
    Span4Mux_v I__8263 (
            .O(N__34807),
            .I(N__34792));
    Span4Mux_h I__8262 (
            .O(N__34804),
            .I(N__34787));
    Span4Mux_h I__8261 (
            .O(N__34801),
            .I(N__34787));
    Span4Mux_h I__8260 (
            .O(N__34798),
            .I(N__34782));
    Span4Mux_h I__8259 (
            .O(N__34795),
            .I(N__34782));
    Odrv4 I__8258 (
            .O(N__34792),
            .I(b2v_inst_data_a_escribir_1));
    Odrv4 I__8257 (
            .O(N__34787),
            .I(b2v_inst_data_a_escribir_1));
    Odrv4 I__8256 (
            .O(N__34782),
            .I(b2v_inst_data_a_escribir_1));
    CascadeMux I__8255 (
            .O(N__34775),
            .I(\b2v_inst.cantidad_temp_RNILL3KZ0Z_1_cascade_ ));
    InMux I__8254 (
            .O(N__34772),
            .I(N__34769));
    LocalMux I__8253 (
            .O(N__34769),
            .I(N_555_i));
    InMux I__8252 (
            .O(N__34766),
            .I(N__34758));
    InMux I__8251 (
            .O(N__34765),
            .I(N__34755));
    InMux I__8250 (
            .O(N__34764),
            .I(N__34752));
    InMux I__8249 (
            .O(N__34763),
            .I(N__34747));
    InMux I__8248 (
            .O(N__34762),
            .I(N__34747));
    InMux I__8247 (
            .O(N__34761),
            .I(N__34742));
    LocalMux I__8246 (
            .O(N__34758),
            .I(N__34738));
    LocalMux I__8245 (
            .O(N__34755),
            .I(N__34731));
    LocalMux I__8244 (
            .O(N__34752),
            .I(N__34731));
    LocalMux I__8243 (
            .O(N__34747),
            .I(N__34731));
    CascadeMux I__8242 (
            .O(N__34746),
            .I(N__34728));
    InMux I__8241 (
            .O(N__34745),
            .I(N__34722));
    LocalMux I__8240 (
            .O(N__34742),
            .I(N__34719));
    InMux I__8239 (
            .O(N__34741),
            .I(N__34716));
    Span4Mux_v I__8238 (
            .O(N__34738),
            .I(N__34713));
    Span4Mux_v I__8237 (
            .O(N__34731),
            .I(N__34710));
    InMux I__8236 (
            .O(N__34728),
            .I(N__34707));
    CascadeMux I__8235 (
            .O(N__34727),
            .I(N__34703));
    InMux I__8234 (
            .O(N__34726),
            .I(N__34698));
    InMux I__8233 (
            .O(N__34725),
            .I(N__34698));
    LocalMux I__8232 (
            .O(N__34722),
            .I(N__34695));
    Span4Mux_h I__8231 (
            .O(N__34719),
            .I(N__34691));
    LocalMux I__8230 (
            .O(N__34716),
            .I(N__34688));
    Sp12to4 I__8229 (
            .O(N__34713),
            .I(N__34681));
    Sp12to4 I__8228 (
            .O(N__34710),
            .I(N__34681));
    LocalMux I__8227 (
            .O(N__34707),
            .I(N__34681));
    InMux I__8226 (
            .O(N__34706),
            .I(N__34676));
    InMux I__8225 (
            .O(N__34703),
            .I(N__34676));
    LocalMux I__8224 (
            .O(N__34698),
            .I(N__34673));
    Span4Mux_h I__8223 (
            .O(N__34695),
            .I(N__34670));
    InMux I__8222 (
            .O(N__34694),
            .I(N__34667));
    Odrv4 I__8221 (
            .O(N__34691),
            .I(\b2v_inst.stateZ0Z_18 ));
    Odrv12 I__8220 (
            .O(N__34688),
            .I(\b2v_inst.stateZ0Z_18 ));
    Odrv12 I__8219 (
            .O(N__34681),
            .I(\b2v_inst.stateZ0Z_18 ));
    LocalMux I__8218 (
            .O(N__34676),
            .I(\b2v_inst.stateZ0Z_18 ));
    Odrv4 I__8217 (
            .O(N__34673),
            .I(\b2v_inst.stateZ0Z_18 ));
    Odrv4 I__8216 (
            .O(N__34670),
            .I(\b2v_inst.stateZ0Z_18 ));
    LocalMux I__8215 (
            .O(N__34667),
            .I(\b2v_inst.stateZ0Z_18 ));
    CascadeMux I__8214 (
            .O(N__34652),
            .I(N__34649));
    InMux I__8213 (
            .O(N__34649),
            .I(N__34646));
    LocalMux I__8212 (
            .O(N__34646),
            .I(SYNTHESIZED_WIRE_1_3));
    InMux I__8211 (
            .O(N__34643),
            .I(N__34639));
    InMux I__8210 (
            .O(N__34642),
            .I(N__34636));
    LocalMux I__8209 (
            .O(N__34639),
            .I(N__34633));
    LocalMux I__8208 (
            .O(N__34636),
            .I(N__34630));
    Span4Mux_v I__8207 (
            .O(N__34633),
            .I(N__34620));
    Span4Mux_v I__8206 (
            .O(N__34630),
            .I(N__34617));
    InMux I__8205 (
            .O(N__34629),
            .I(N__34610));
    InMux I__8204 (
            .O(N__34628),
            .I(N__34610));
    InMux I__8203 (
            .O(N__34627),
            .I(N__34610));
    InMux I__8202 (
            .O(N__34626),
            .I(N__34607));
    InMux I__8201 (
            .O(N__34625),
            .I(N__34604));
    InMux I__8200 (
            .O(N__34624),
            .I(N__34599));
    InMux I__8199 (
            .O(N__34623),
            .I(N__34599));
    Sp12to4 I__8198 (
            .O(N__34620),
            .I(N__34592));
    Sp12to4 I__8197 (
            .O(N__34617),
            .I(N__34592));
    LocalMux I__8196 (
            .O(N__34610),
            .I(N__34592));
    LocalMux I__8195 (
            .O(N__34607),
            .I(N__34589));
    LocalMux I__8194 (
            .O(N__34604),
            .I(N__34583));
    LocalMux I__8193 (
            .O(N__34599),
            .I(N__34583));
    Span12Mux_h I__8192 (
            .O(N__34592),
            .I(N__34579));
    Span4Mux_h I__8191 (
            .O(N__34589),
            .I(N__34576));
    InMux I__8190 (
            .O(N__34588),
            .I(N__34573));
    Span4Mux_h I__8189 (
            .O(N__34583),
            .I(N__34570));
    InMux I__8188 (
            .O(N__34582),
            .I(N__34567));
    Odrv12 I__8187 (
            .O(N__34579),
            .I(\b2v_inst.stateZ0Z_9 ));
    Odrv4 I__8186 (
            .O(N__34576),
            .I(\b2v_inst.stateZ0Z_9 ));
    LocalMux I__8185 (
            .O(N__34573),
            .I(\b2v_inst.stateZ0Z_9 ));
    Odrv4 I__8184 (
            .O(N__34570),
            .I(\b2v_inst.stateZ0Z_9 ));
    LocalMux I__8183 (
            .O(N__34567),
            .I(\b2v_inst.stateZ0Z_9 ));
    InMux I__8182 (
            .O(N__34556),
            .I(N__34553));
    LocalMux I__8181 (
            .O(N__34553),
            .I(N__34550));
    Span4Mux_h I__8180 (
            .O(N__34550),
            .I(N__34546));
    InMux I__8179 (
            .O(N__34549),
            .I(N__34542));
    Span4Mux_h I__8178 (
            .O(N__34546),
            .I(N__34539));
    InMux I__8177 (
            .O(N__34545),
            .I(N__34536));
    LocalMux I__8176 (
            .O(N__34542),
            .I(b2v_inst_cantidad_temp_3));
    Odrv4 I__8175 (
            .O(N__34539),
            .I(b2v_inst_cantidad_temp_3));
    LocalMux I__8174 (
            .O(N__34536),
            .I(b2v_inst_cantidad_temp_3));
    ClkMux I__8173 (
            .O(N__34529),
            .I(N__34052));
    ClkMux I__8172 (
            .O(N__34528),
            .I(N__34052));
    ClkMux I__8171 (
            .O(N__34527),
            .I(N__34052));
    ClkMux I__8170 (
            .O(N__34526),
            .I(N__34052));
    ClkMux I__8169 (
            .O(N__34525),
            .I(N__34052));
    ClkMux I__8168 (
            .O(N__34524),
            .I(N__34052));
    ClkMux I__8167 (
            .O(N__34523),
            .I(N__34052));
    ClkMux I__8166 (
            .O(N__34522),
            .I(N__34052));
    ClkMux I__8165 (
            .O(N__34521),
            .I(N__34052));
    ClkMux I__8164 (
            .O(N__34520),
            .I(N__34052));
    ClkMux I__8163 (
            .O(N__34519),
            .I(N__34052));
    ClkMux I__8162 (
            .O(N__34518),
            .I(N__34052));
    ClkMux I__8161 (
            .O(N__34517),
            .I(N__34052));
    ClkMux I__8160 (
            .O(N__34516),
            .I(N__34052));
    ClkMux I__8159 (
            .O(N__34515),
            .I(N__34052));
    ClkMux I__8158 (
            .O(N__34514),
            .I(N__34052));
    ClkMux I__8157 (
            .O(N__34513),
            .I(N__34052));
    ClkMux I__8156 (
            .O(N__34512),
            .I(N__34052));
    ClkMux I__8155 (
            .O(N__34511),
            .I(N__34052));
    ClkMux I__8154 (
            .O(N__34510),
            .I(N__34052));
    ClkMux I__8153 (
            .O(N__34509),
            .I(N__34052));
    ClkMux I__8152 (
            .O(N__34508),
            .I(N__34052));
    ClkMux I__8151 (
            .O(N__34507),
            .I(N__34052));
    ClkMux I__8150 (
            .O(N__34506),
            .I(N__34052));
    ClkMux I__8149 (
            .O(N__34505),
            .I(N__34052));
    ClkMux I__8148 (
            .O(N__34504),
            .I(N__34052));
    ClkMux I__8147 (
            .O(N__34503),
            .I(N__34052));
    ClkMux I__8146 (
            .O(N__34502),
            .I(N__34052));
    ClkMux I__8145 (
            .O(N__34501),
            .I(N__34052));
    ClkMux I__8144 (
            .O(N__34500),
            .I(N__34052));
    ClkMux I__8143 (
            .O(N__34499),
            .I(N__34052));
    ClkMux I__8142 (
            .O(N__34498),
            .I(N__34052));
    ClkMux I__8141 (
            .O(N__34497),
            .I(N__34052));
    ClkMux I__8140 (
            .O(N__34496),
            .I(N__34052));
    ClkMux I__8139 (
            .O(N__34495),
            .I(N__34052));
    ClkMux I__8138 (
            .O(N__34494),
            .I(N__34052));
    ClkMux I__8137 (
            .O(N__34493),
            .I(N__34052));
    ClkMux I__8136 (
            .O(N__34492),
            .I(N__34052));
    ClkMux I__8135 (
            .O(N__34491),
            .I(N__34052));
    ClkMux I__8134 (
            .O(N__34490),
            .I(N__34052));
    ClkMux I__8133 (
            .O(N__34489),
            .I(N__34052));
    ClkMux I__8132 (
            .O(N__34488),
            .I(N__34052));
    ClkMux I__8131 (
            .O(N__34487),
            .I(N__34052));
    ClkMux I__8130 (
            .O(N__34486),
            .I(N__34052));
    ClkMux I__8129 (
            .O(N__34485),
            .I(N__34052));
    ClkMux I__8128 (
            .O(N__34484),
            .I(N__34052));
    ClkMux I__8127 (
            .O(N__34483),
            .I(N__34052));
    ClkMux I__8126 (
            .O(N__34482),
            .I(N__34052));
    ClkMux I__8125 (
            .O(N__34481),
            .I(N__34052));
    ClkMux I__8124 (
            .O(N__34480),
            .I(N__34052));
    ClkMux I__8123 (
            .O(N__34479),
            .I(N__34052));
    ClkMux I__8122 (
            .O(N__34478),
            .I(N__34052));
    ClkMux I__8121 (
            .O(N__34477),
            .I(N__34052));
    ClkMux I__8120 (
            .O(N__34476),
            .I(N__34052));
    ClkMux I__8119 (
            .O(N__34475),
            .I(N__34052));
    ClkMux I__8118 (
            .O(N__34474),
            .I(N__34052));
    ClkMux I__8117 (
            .O(N__34473),
            .I(N__34052));
    ClkMux I__8116 (
            .O(N__34472),
            .I(N__34052));
    ClkMux I__8115 (
            .O(N__34471),
            .I(N__34052));
    ClkMux I__8114 (
            .O(N__34470),
            .I(N__34052));
    ClkMux I__8113 (
            .O(N__34469),
            .I(N__34052));
    ClkMux I__8112 (
            .O(N__34468),
            .I(N__34052));
    ClkMux I__8111 (
            .O(N__34467),
            .I(N__34052));
    ClkMux I__8110 (
            .O(N__34466),
            .I(N__34052));
    ClkMux I__8109 (
            .O(N__34465),
            .I(N__34052));
    ClkMux I__8108 (
            .O(N__34464),
            .I(N__34052));
    ClkMux I__8107 (
            .O(N__34463),
            .I(N__34052));
    ClkMux I__8106 (
            .O(N__34462),
            .I(N__34052));
    ClkMux I__8105 (
            .O(N__34461),
            .I(N__34052));
    ClkMux I__8104 (
            .O(N__34460),
            .I(N__34052));
    ClkMux I__8103 (
            .O(N__34459),
            .I(N__34052));
    ClkMux I__8102 (
            .O(N__34458),
            .I(N__34052));
    ClkMux I__8101 (
            .O(N__34457),
            .I(N__34052));
    ClkMux I__8100 (
            .O(N__34456),
            .I(N__34052));
    ClkMux I__8099 (
            .O(N__34455),
            .I(N__34052));
    ClkMux I__8098 (
            .O(N__34454),
            .I(N__34052));
    ClkMux I__8097 (
            .O(N__34453),
            .I(N__34052));
    ClkMux I__8096 (
            .O(N__34452),
            .I(N__34052));
    ClkMux I__8095 (
            .O(N__34451),
            .I(N__34052));
    ClkMux I__8094 (
            .O(N__34450),
            .I(N__34052));
    ClkMux I__8093 (
            .O(N__34449),
            .I(N__34052));
    ClkMux I__8092 (
            .O(N__34448),
            .I(N__34052));
    ClkMux I__8091 (
            .O(N__34447),
            .I(N__34052));
    ClkMux I__8090 (
            .O(N__34446),
            .I(N__34052));
    ClkMux I__8089 (
            .O(N__34445),
            .I(N__34052));
    ClkMux I__8088 (
            .O(N__34444),
            .I(N__34052));
    ClkMux I__8087 (
            .O(N__34443),
            .I(N__34052));
    ClkMux I__8086 (
            .O(N__34442),
            .I(N__34052));
    ClkMux I__8085 (
            .O(N__34441),
            .I(N__34052));
    ClkMux I__8084 (
            .O(N__34440),
            .I(N__34052));
    ClkMux I__8083 (
            .O(N__34439),
            .I(N__34052));
    ClkMux I__8082 (
            .O(N__34438),
            .I(N__34052));
    ClkMux I__8081 (
            .O(N__34437),
            .I(N__34052));
    ClkMux I__8080 (
            .O(N__34436),
            .I(N__34052));
    ClkMux I__8079 (
            .O(N__34435),
            .I(N__34052));
    ClkMux I__8078 (
            .O(N__34434),
            .I(N__34052));
    ClkMux I__8077 (
            .O(N__34433),
            .I(N__34052));
    ClkMux I__8076 (
            .O(N__34432),
            .I(N__34052));
    ClkMux I__8075 (
            .O(N__34431),
            .I(N__34052));
    ClkMux I__8074 (
            .O(N__34430),
            .I(N__34052));
    ClkMux I__8073 (
            .O(N__34429),
            .I(N__34052));
    ClkMux I__8072 (
            .O(N__34428),
            .I(N__34052));
    ClkMux I__8071 (
            .O(N__34427),
            .I(N__34052));
    ClkMux I__8070 (
            .O(N__34426),
            .I(N__34052));
    ClkMux I__8069 (
            .O(N__34425),
            .I(N__34052));
    ClkMux I__8068 (
            .O(N__34424),
            .I(N__34052));
    ClkMux I__8067 (
            .O(N__34423),
            .I(N__34052));
    ClkMux I__8066 (
            .O(N__34422),
            .I(N__34052));
    ClkMux I__8065 (
            .O(N__34421),
            .I(N__34052));
    ClkMux I__8064 (
            .O(N__34420),
            .I(N__34052));
    ClkMux I__8063 (
            .O(N__34419),
            .I(N__34052));
    ClkMux I__8062 (
            .O(N__34418),
            .I(N__34052));
    ClkMux I__8061 (
            .O(N__34417),
            .I(N__34052));
    ClkMux I__8060 (
            .O(N__34416),
            .I(N__34052));
    ClkMux I__8059 (
            .O(N__34415),
            .I(N__34052));
    ClkMux I__8058 (
            .O(N__34414),
            .I(N__34052));
    ClkMux I__8057 (
            .O(N__34413),
            .I(N__34052));
    ClkMux I__8056 (
            .O(N__34412),
            .I(N__34052));
    ClkMux I__8055 (
            .O(N__34411),
            .I(N__34052));
    ClkMux I__8054 (
            .O(N__34410),
            .I(N__34052));
    ClkMux I__8053 (
            .O(N__34409),
            .I(N__34052));
    ClkMux I__8052 (
            .O(N__34408),
            .I(N__34052));
    ClkMux I__8051 (
            .O(N__34407),
            .I(N__34052));
    ClkMux I__8050 (
            .O(N__34406),
            .I(N__34052));
    ClkMux I__8049 (
            .O(N__34405),
            .I(N__34052));
    ClkMux I__8048 (
            .O(N__34404),
            .I(N__34052));
    ClkMux I__8047 (
            .O(N__34403),
            .I(N__34052));
    ClkMux I__8046 (
            .O(N__34402),
            .I(N__34052));
    ClkMux I__8045 (
            .O(N__34401),
            .I(N__34052));
    ClkMux I__8044 (
            .O(N__34400),
            .I(N__34052));
    ClkMux I__8043 (
            .O(N__34399),
            .I(N__34052));
    ClkMux I__8042 (
            .O(N__34398),
            .I(N__34052));
    ClkMux I__8041 (
            .O(N__34397),
            .I(N__34052));
    ClkMux I__8040 (
            .O(N__34396),
            .I(N__34052));
    ClkMux I__8039 (
            .O(N__34395),
            .I(N__34052));
    ClkMux I__8038 (
            .O(N__34394),
            .I(N__34052));
    ClkMux I__8037 (
            .O(N__34393),
            .I(N__34052));
    ClkMux I__8036 (
            .O(N__34392),
            .I(N__34052));
    ClkMux I__8035 (
            .O(N__34391),
            .I(N__34052));
    ClkMux I__8034 (
            .O(N__34390),
            .I(N__34052));
    ClkMux I__8033 (
            .O(N__34389),
            .I(N__34052));
    ClkMux I__8032 (
            .O(N__34388),
            .I(N__34052));
    ClkMux I__8031 (
            .O(N__34387),
            .I(N__34052));
    ClkMux I__8030 (
            .O(N__34386),
            .I(N__34052));
    ClkMux I__8029 (
            .O(N__34385),
            .I(N__34052));
    ClkMux I__8028 (
            .O(N__34384),
            .I(N__34052));
    ClkMux I__8027 (
            .O(N__34383),
            .I(N__34052));
    ClkMux I__8026 (
            .O(N__34382),
            .I(N__34052));
    ClkMux I__8025 (
            .O(N__34381),
            .I(N__34052));
    ClkMux I__8024 (
            .O(N__34380),
            .I(N__34052));
    ClkMux I__8023 (
            .O(N__34379),
            .I(N__34052));
    ClkMux I__8022 (
            .O(N__34378),
            .I(N__34052));
    ClkMux I__8021 (
            .O(N__34377),
            .I(N__34052));
    ClkMux I__8020 (
            .O(N__34376),
            .I(N__34052));
    ClkMux I__8019 (
            .O(N__34375),
            .I(N__34052));
    ClkMux I__8018 (
            .O(N__34374),
            .I(N__34052));
    ClkMux I__8017 (
            .O(N__34373),
            .I(N__34052));
    ClkMux I__8016 (
            .O(N__34372),
            .I(N__34052));
    ClkMux I__8015 (
            .O(N__34371),
            .I(N__34052));
    GlobalMux I__8014 (
            .O(N__34052),
            .I(N__34049));
    gio2CtrlBuf I__8013 (
            .O(N__34049),
            .I(clk_c_g));
    InMux I__8012 (
            .O(N__34046),
            .I(N__34043));
    LocalMux I__8011 (
            .O(N__34043),
            .I(N__34040));
    Span4Mux_h I__8010 (
            .O(N__34040),
            .I(N__34037));
    Span4Mux_h I__8009 (
            .O(N__34037),
            .I(N__34034));
    Odrv4 I__8008 (
            .O(N__34034),
            .I(\b2v_inst.addr_ram_iv_i_0_5 ));
    CascadeMux I__8007 (
            .O(N__34031),
            .I(N__34028));
    InMux I__8006 (
            .O(N__34028),
            .I(N__34025));
    LocalMux I__8005 (
            .O(N__34025),
            .I(N__34022));
    Span4Mux_v I__8004 (
            .O(N__34022),
            .I(N__34019));
    Span4Mux_h I__8003 (
            .O(N__34019),
            .I(N__34016));
    Span4Mux_h I__8002 (
            .O(N__34016),
            .I(N__34013));
    Odrv4 I__8001 (
            .O(N__34013),
            .I(\b2v_inst.addr_ram_iv_i_1_5 ));
    CascadeMux I__8000 (
            .O(N__34010),
            .I(N__34006));
    CascadeMux I__7999 (
            .O(N__34009),
            .I(N__34003));
    CascadeBuf I__7998 (
            .O(N__34006),
            .I(N__34000));
    CascadeBuf I__7997 (
            .O(N__34003),
            .I(N__33997));
    CascadeMux I__7996 (
            .O(N__34000),
            .I(N__33994));
    CascadeMux I__7995 (
            .O(N__33997),
            .I(N__33991));
    CascadeBuf I__7994 (
            .O(N__33994),
            .I(N__33988));
    CascadeBuf I__7993 (
            .O(N__33991),
            .I(N__33985));
    CascadeMux I__7992 (
            .O(N__33988),
            .I(N__33982));
    CascadeMux I__7991 (
            .O(N__33985),
            .I(N__33979));
    CascadeBuf I__7990 (
            .O(N__33982),
            .I(N__33976));
    CascadeBuf I__7989 (
            .O(N__33979),
            .I(N__33973));
    CascadeMux I__7988 (
            .O(N__33976),
            .I(N__33970));
    CascadeMux I__7987 (
            .O(N__33973),
            .I(N__33967));
    CascadeBuf I__7986 (
            .O(N__33970),
            .I(N__33964));
    CascadeBuf I__7985 (
            .O(N__33967),
            .I(N__33961));
    CascadeMux I__7984 (
            .O(N__33964),
            .I(N__33958));
    CascadeMux I__7983 (
            .O(N__33961),
            .I(N__33955));
    CascadeBuf I__7982 (
            .O(N__33958),
            .I(N__33952));
    CascadeBuf I__7981 (
            .O(N__33955),
            .I(N__33949));
    CascadeMux I__7980 (
            .O(N__33952),
            .I(N__33946));
    CascadeMux I__7979 (
            .O(N__33949),
            .I(N__33943));
    InMux I__7978 (
            .O(N__33946),
            .I(N__33940));
    InMux I__7977 (
            .O(N__33943),
            .I(N__33937));
    LocalMux I__7976 (
            .O(N__33940),
            .I(N__33934));
    LocalMux I__7975 (
            .O(N__33937),
            .I(indice_RNIS8333_5));
    Odrv4 I__7974 (
            .O(N__33934),
            .I(indice_RNIS8333_5));
    InMux I__7973 (
            .O(N__33929),
            .I(N__33926));
    LocalMux I__7972 (
            .O(N__33926),
            .I(N__33923));
    Span4Mux_h I__7971 (
            .O(N__33923),
            .I(N__33920));
    Span4Mux_h I__7970 (
            .O(N__33920),
            .I(N__33917));
    Span4Mux_h I__7969 (
            .O(N__33917),
            .I(N__33914));
    Odrv4 I__7968 (
            .O(N__33914),
            .I(\b2v_inst.addr_ram_iv_i_0_8 ));
    CascadeMux I__7967 (
            .O(N__33911),
            .I(N__33908));
    InMux I__7966 (
            .O(N__33908),
            .I(N__33905));
    LocalMux I__7965 (
            .O(N__33905),
            .I(N__33902));
    Span4Mux_v I__7964 (
            .O(N__33902),
            .I(N__33899));
    Sp12to4 I__7963 (
            .O(N__33899),
            .I(N__33896));
    Odrv12 I__7962 (
            .O(N__33896),
            .I(\b2v_inst.addr_ram_iv_i_1_8 ));
    CascadeMux I__7961 (
            .O(N__33893),
            .I(N__33889));
    CascadeMux I__7960 (
            .O(N__33892),
            .I(N__33886));
    CascadeBuf I__7959 (
            .O(N__33889),
            .I(N__33883));
    CascadeBuf I__7958 (
            .O(N__33886),
            .I(N__33880));
    CascadeMux I__7957 (
            .O(N__33883),
            .I(N__33877));
    CascadeMux I__7956 (
            .O(N__33880),
            .I(N__33874));
    CascadeBuf I__7955 (
            .O(N__33877),
            .I(N__33871));
    CascadeBuf I__7954 (
            .O(N__33874),
            .I(N__33868));
    CascadeMux I__7953 (
            .O(N__33871),
            .I(N__33865));
    CascadeMux I__7952 (
            .O(N__33868),
            .I(N__33862));
    CascadeBuf I__7951 (
            .O(N__33865),
            .I(N__33859));
    CascadeBuf I__7950 (
            .O(N__33862),
            .I(N__33856));
    CascadeMux I__7949 (
            .O(N__33859),
            .I(N__33853));
    CascadeMux I__7948 (
            .O(N__33856),
            .I(N__33850));
    CascadeBuf I__7947 (
            .O(N__33853),
            .I(N__33847));
    CascadeBuf I__7946 (
            .O(N__33850),
            .I(N__33844));
    CascadeMux I__7945 (
            .O(N__33847),
            .I(N__33841));
    CascadeMux I__7944 (
            .O(N__33844),
            .I(N__33838));
    CascadeBuf I__7943 (
            .O(N__33841),
            .I(N__33835));
    CascadeBuf I__7942 (
            .O(N__33838),
            .I(N__33832));
    CascadeMux I__7941 (
            .O(N__33835),
            .I(N__33829));
    CascadeMux I__7940 (
            .O(N__33832),
            .I(N__33826));
    InMux I__7939 (
            .O(N__33829),
            .I(N__33823));
    InMux I__7938 (
            .O(N__33826),
            .I(N__33820));
    LocalMux I__7937 (
            .O(N__33823),
            .I(N__33817));
    LocalMux I__7936 (
            .O(N__33820),
            .I(indice_RNIBO333_8));
    Odrv4 I__7935 (
            .O(N__33817),
            .I(indice_RNIBO333_8));
    InMux I__7934 (
            .O(N__33812),
            .I(N__33809));
    LocalMux I__7933 (
            .O(N__33809),
            .I(N__33806));
    Span4Mux_v I__7932 (
            .O(N__33806),
            .I(N__33803));
    Span4Mux_h I__7931 (
            .O(N__33803),
            .I(N__33800));
    Odrv4 I__7930 (
            .O(N__33800),
            .I(\b2v_inst.addr_ram_iv_i_0_9 ));
    CascadeMux I__7929 (
            .O(N__33797),
            .I(N__33794));
    InMux I__7928 (
            .O(N__33794),
            .I(N__33791));
    LocalMux I__7927 (
            .O(N__33791),
            .I(N__33788));
    Span4Mux_h I__7926 (
            .O(N__33788),
            .I(N__33785));
    Span4Mux_h I__7925 (
            .O(N__33785),
            .I(N__33782));
    Odrv4 I__7924 (
            .O(N__33782),
            .I(\b2v_inst.addr_ram_iv_i_1_9 ));
    CascadeMux I__7923 (
            .O(N__33779),
            .I(N__33775));
    CascadeMux I__7922 (
            .O(N__33778),
            .I(N__33772));
    CascadeBuf I__7921 (
            .O(N__33775),
            .I(N__33769));
    CascadeBuf I__7920 (
            .O(N__33772),
            .I(N__33766));
    CascadeMux I__7919 (
            .O(N__33769),
            .I(N__33763));
    CascadeMux I__7918 (
            .O(N__33766),
            .I(N__33760));
    CascadeBuf I__7917 (
            .O(N__33763),
            .I(N__33757));
    CascadeBuf I__7916 (
            .O(N__33760),
            .I(N__33754));
    CascadeMux I__7915 (
            .O(N__33757),
            .I(N__33751));
    CascadeMux I__7914 (
            .O(N__33754),
            .I(N__33748));
    CascadeBuf I__7913 (
            .O(N__33751),
            .I(N__33745));
    CascadeBuf I__7912 (
            .O(N__33748),
            .I(N__33742));
    CascadeMux I__7911 (
            .O(N__33745),
            .I(N__33739));
    CascadeMux I__7910 (
            .O(N__33742),
            .I(N__33736));
    CascadeBuf I__7909 (
            .O(N__33739),
            .I(N__33733));
    CascadeBuf I__7908 (
            .O(N__33736),
            .I(N__33730));
    CascadeMux I__7907 (
            .O(N__33733),
            .I(N__33727));
    CascadeMux I__7906 (
            .O(N__33730),
            .I(N__33724));
    CascadeBuf I__7905 (
            .O(N__33727),
            .I(N__33721));
    CascadeBuf I__7904 (
            .O(N__33724),
            .I(N__33718));
    CascadeMux I__7903 (
            .O(N__33721),
            .I(N__33715));
    CascadeMux I__7902 (
            .O(N__33718),
            .I(N__33712));
    InMux I__7901 (
            .O(N__33715),
            .I(N__33709));
    InMux I__7900 (
            .O(N__33712),
            .I(N__33706));
    LocalMux I__7899 (
            .O(N__33709),
            .I(N__33703));
    LocalMux I__7898 (
            .O(N__33706),
            .I(indice_RNIGT333_9));
    Odrv4 I__7897 (
            .O(N__33703),
            .I(indice_RNIGT333_9));
    InMux I__7896 (
            .O(N__33698),
            .I(N__33695));
    LocalMux I__7895 (
            .O(N__33695),
            .I(N__33692));
    Span4Mux_v I__7894 (
            .O(N__33692),
            .I(N__33689));
    Odrv4 I__7893 (
            .O(N__33689),
            .I(N_115_i));
    CascadeMux I__7892 (
            .O(N__33686),
            .I(N__33683));
    InMux I__7891 (
            .O(N__33683),
            .I(N__33679));
    CascadeMux I__7890 (
            .O(N__33682),
            .I(N__33676));
    LocalMux I__7889 (
            .O(N__33679),
            .I(N__33673));
    InMux I__7888 (
            .O(N__33676),
            .I(N__33670));
    Span4Mux_v I__7887 (
            .O(N__33673),
            .I(N__33664));
    LocalMux I__7886 (
            .O(N__33670),
            .I(N__33664));
    InMux I__7885 (
            .O(N__33669),
            .I(N__33661));
    Span4Mux_h I__7884 (
            .O(N__33664),
            .I(N__33658));
    LocalMux I__7883 (
            .O(N__33661),
            .I(N__33655));
    Span4Mux_v I__7882 (
            .O(N__33658),
            .I(N__33652));
    Span4Mux_h I__7881 (
            .O(N__33655),
            .I(N__33649));
    Sp12to4 I__7880 (
            .O(N__33652),
            .I(N__33645));
    Span4Mux_h I__7879 (
            .O(N__33649),
            .I(N__33642));
    InMux I__7878 (
            .O(N__33648),
            .I(N__33639));
    Odrv12 I__7877 (
            .O(N__33645),
            .I(b2v_inst_data_a_escribir_10));
    Odrv4 I__7876 (
            .O(N__33642),
            .I(b2v_inst_data_a_escribir_10));
    LocalMux I__7875 (
            .O(N__33639),
            .I(b2v_inst_data_a_escribir_10));
    InMux I__7874 (
            .O(N__33632),
            .I(N__33629));
    LocalMux I__7873 (
            .O(N__33629),
            .I(N__33626));
    Span4Mux_v I__7872 (
            .O(N__33626),
            .I(N__33623));
    Odrv4 I__7871 (
            .O(N__33623),
            .I(N_110_i));
    InMux I__7870 (
            .O(N__33620),
            .I(N__33617));
    LocalMux I__7869 (
            .O(N__33617),
            .I(N__33614));
    Span4Mux_h I__7868 (
            .O(N__33614),
            .I(N__33611));
    Span4Mux_h I__7867 (
            .O(N__33611),
            .I(N__33608));
    Odrv4 I__7866 (
            .O(N__33608),
            .I(\b2v_inst.addr_ram_iv_i_0_0 ));
    CascadeMux I__7865 (
            .O(N__33605),
            .I(N__33602));
    InMux I__7864 (
            .O(N__33602),
            .I(N__33599));
    LocalMux I__7863 (
            .O(N__33599),
            .I(N__33596));
    Span12Mux_s9_h I__7862 (
            .O(N__33596),
            .I(N__33593));
    Odrv12 I__7861 (
            .O(N__33593),
            .I(\b2v_inst.addr_ram_iv_i_1_0 ));
    CascadeMux I__7860 (
            .O(N__33590),
            .I(N__33586));
    CascadeMux I__7859 (
            .O(N__33589),
            .I(N__33583));
    CascadeBuf I__7858 (
            .O(N__33586),
            .I(N__33580));
    CascadeBuf I__7857 (
            .O(N__33583),
            .I(N__33577));
    CascadeMux I__7856 (
            .O(N__33580),
            .I(N__33574));
    CascadeMux I__7855 (
            .O(N__33577),
            .I(N__33571));
    CascadeBuf I__7854 (
            .O(N__33574),
            .I(N__33568));
    CascadeBuf I__7853 (
            .O(N__33571),
            .I(N__33565));
    CascadeMux I__7852 (
            .O(N__33568),
            .I(N__33562));
    CascadeMux I__7851 (
            .O(N__33565),
            .I(N__33559));
    CascadeBuf I__7850 (
            .O(N__33562),
            .I(N__33556));
    CascadeBuf I__7849 (
            .O(N__33559),
            .I(N__33553));
    CascadeMux I__7848 (
            .O(N__33556),
            .I(N__33550));
    CascadeMux I__7847 (
            .O(N__33553),
            .I(N__33547));
    CascadeBuf I__7846 (
            .O(N__33550),
            .I(N__33544));
    CascadeBuf I__7845 (
            .O(N__33547),
            .I(N__33541));
    CascadeMux I__7844 (
            .O(N__33544),
            .I(N__33538));
    CascadeMux I__7843 (
            .O(N__33541),
            .I(N__33535));
    CascadeBuf I__7842 (
            .O(N__33538),
            .I(N__33532));
    CascadeBuf I__7841 (
            .O(N__33535),
            .I(N__33529));
    CascadeMux I__7840 (
            .O(N__33532),
            .I(N__33526));
    CascadeMux I__7839 (
            .O(N__33529),
            .I(N__33523));
    InMux I__7838 (
            .O(N__33526),
            .I(N__33520));
    InMux I__7837 (
            .O(N__33523),
            .I(N__33517));
    LocalMux I__7836 (
            .O(N__33520),
            .I(indice_RNI3F233_0));
    LocalMux I__7835 (
            .O(N__33517),
            .I(indice_RNI3F233_0));
    InMux I__7834 (
            .O(N__33512),
            .I(N__33509));
    LocalMux I__7833 (
            .O(N__33509),
            .I(N__33506));
    Span4Mux_v I__7832 (
            .O(N__33506),
            .I(N__33503));
    Span4Mux_h I__7831 (
            .O(N__33503),
            .I(N__33500));
    Span4Mux_h I__7830 (
            .O(N__33500),
            .I(N__33497));
    Odrv4 I__7829 (
            .O(N__33497),
            .I(\b2v_inst.addr_ram_iv_i_0_10 ));
    CascadeMux I__7828 (
            .O(N__33494),
            .I(N__33491));
    InMux I__7827 (
            .O(N__33491),
            .I(N__33488));
    LocalMux I__7826 (
            .O(N__33488),
            .I(N__33485));
    Span4Mux_h I__7825 (
            .O(N__33485),
            .I(N__33482));
    Span4Mux_h I__7824 (
            .O(N__33482),
            .I(N__33479));
    Odrv4 I__7823 (
            .O(N__33479),
            .I(\b2v_inst.addr_ram_iv_i_1_10 ));
    CascadeMux I__7822 (
            .O(N__33476),
            .I(N__33472));
    CascadeMux I__7821 (
            .O(N__33475),
            .I(N__33469));
    CascadeBuf I__7820 (
            .O(N__33472),
            .I(N__33466));
    CascadeBuf I__7819 (
            .O(N__33469),
            .I(N__33463));
    CascadeMux I__7818 (
            .O(N__33466),
            .I(N__33460));
    CascadeMux I__7817 (
            .O(N__33463),
            .I(N__33457));
    CascadeBuf I__7816 (
            .O(N__33460),
            .I(N__33454));
    CascadeBuf I__7815 (
            .O(N__33457),
            .I(N__33451));
    CascadeMux I__7814 (
            .O(N__33454),
            .I(N__33448));
    CascadeMux I__7813 (
            .O(N__33451),
            .I(N__33445));
    CascadeBuf I__7812 (
            .O(N__33448),
            .I(N__33442));
    CascadeBuf I__7811 (
            .O(N__33445),
            .I(N__33439));
    CascadeMux I__7810 (
            .O(N__33442),
            .I(N__33436));
    CascadeMux I__7809 (
            .O(N__33439),
            .I(N__33433));
    CascadeBuf I__7808 (
            .O(N__33436),
            .I(N__33430));
    CascadeBuf I__7807 (
            .O(N__33433),
            .I(N__33427));
    CascadeMux I__7806 (
            .O(N__33430),
            .I(N__33424));
    CascadeMux I__7805 (
            .O(N__33427),
            .I(N__33421));
    CascadeBuf I__7804 (
            .O(N__33424),
            .I(N__33418));
    CascadeBuf I__7803 (
            .O(N__33421),
            .I(N__33415));
    CascadeMux I__7802 (
            .O(N__33418),
            .I(N__33412));
    CascadeMux I__7801 (
            .O(N__33415),
            .I(N__33409));
    InMux I__7800 (
            .O(N__33412),
            .I(N__33406));
    InMux I__7799 (
            .O(N__33409),
            .I(N__33403));
    LocalMux I__7798 (
            .O(N__33406),
            .I(N_37));
    LocalMux I__7797 (
            .O(N__33403),
            .I(N_37));
    CascadeMux I__7796 (
            .O(N__33398),
            .I(N__33394));
    CascadeMux I__7795 (
            .O(N__33397),
            .I(N__33391));
    InMux I__7794 (
            .O(N__33394),
            .I(N__33388));
    InMux I__7793 (
            .O(N__33391),
            .I(N__33385));
    LocalMux I__7792 (
            .O(N__33388),
            .I(N__33382));
    LocalMux I__7791 (
            .O(N__33385),
            .I(N__33375));
    Sp12to4 I__7790 (
            .O(N__33382),
            .I(N__33375));
    InMux I__7789 (
            .O(N__33381),
            .I(N__33372));
    InMux I__7788 (
            .O(N__33380),
            .I(N__33369));
    Span12Mux_h I__7787 (
            .O(N__33375),
            .I(N__33366));
    LocalMux I__7786 (
            .O(N__33372),
            .I(N__33361));
    LocalMux I__7785 (
            .O(N__33369),
            .I(N__33361));
    Odrv12 I__7784 (
            .O(N__33366),
            .I(b2v_inst_data_a_escribir_8));
    Odrv12 I__7783 (
            .O(N__33361),
            .I(b2v_inst_data_a_escribir_8));
    InMux I__7782 (
            .O(N__33356),
            .I(N__33353));
    LocalMux I__7781 (
            .O(N__33353),
            .I(N__33350));
    Odrv4 I__7780 (
            .O(N__33350),
            .I(N_112_i));
    InMux I__7779 (
            .O(N__33347),
            .I(N__33344));
    LocalMux I__7778 (
            .O(N__33344),
            .I(\b2v_inst.un16_data_ram_cantidad_o_cry_3_c_RNIBDEOZ0 ));
    CascadeMux I__7777 (
            .O(N__33341),
            .I(N__33338));
    InMux I__7776 (
            .O(N__33338),
            .I(N__33333));
    InMux I__7775 (
            .O(N__33337),
            .I(N__33330));
    CascadeMux I__7774 (
            .O(N__33336),
            .I(N__33326));
    LocalMux I__7773 (
            .O(N__33333),
            .I(N__33322));
    LocalMux I__7772 (
            .O(N__33330),
            .I(N__33319));
    CascadeMux I__7771 (
            .O(N__33329),
            .I(N__33316));
    InMux I__7770 (
            .O(N__33326),
            .I(N__33313));
    InMux I__7769 (
            .O(N__33325),
            .I(N__33310));
    Span4Mux_v I__7768 (
            .O(N__33322),
            .I(N__33305));
    Span4Mux_v I__7767 (
            .O(N__33319),
            .I(N__33305));
    InMux I__7766 (
            .O(N__33316),
            .I(N__33302));
    LocalMux I__7765 (
            .O(N__33313),
            .I(N__33297));
    LocalMux I__7764 (
            .O(N__33310),
            .I(N__33297));
    Sp12to4 I__7763 (
            .O(N__33305),
            .I(N__33294));
    LocalMux I__7762 (
            .O(N__33302),
            .I(N__33291));
    Span4Mux_v I__7761 (
            .O(N__33297),
            .I(N__33288));
    Span12Mux_h I__7760 (
            .O(N__33294),
            .I(N__33285));
    Span4Mux_h I__7759 (
            .O(N__33291),
            .I(N__33280));
    Span4Mux_h I__7758 (
            .O(N__33288),
            .I(N__33280));
    Odrv12 I__7757 (
            .O(N__33285),
            .I(b2v_inst_data_a_escribir_4));
    Odrv4 I__7756 (
            .O(N__33280),
            .I(b2v_inst_data_a_escribir_4));
    InMux I__7755 (
            .O(N__33275),
            .I(N__33272));
    LocalMux I__7754 (
            .O(N__33272),
            .I(N__33269));
    Span4Mux_h I__7753 (
            .O(N__33269),
            .I(N__33266));
    Odrv4 I__7752 (
            .O(N__33266),
            .I(N_549_i));
    InMux I__7751 (
            .O(N__33263),
            .I(N__33260));
    LocalMux I__7750 (
            .O(N__33260),
            .I(\b2v_inst.un16_data_ram_cantidad_o_cry_2_c_RNI9ADOZ0 ));
    CascadeMux I__7749 (
            .O(N__33257),
            .I(N__33251));
    InMux I__7748 (
            .O(N__33256),
            .I(N__33248));
    CascadeMux I__7747 (
            .O(N__33255),
            .I(N__33245));
    InMux I__7746 (
            .O(N__33254),
            .I(N__33241));
    InMux I__7745 (
            .O(N__33251),
            .I(N__33238));
    LocalMux I__7744 (
            .O(N__33248),
            .I(N__33235));
    InMux I__7743 (
            .O(N__33245),
            .I(N__33232));
    InMux I__7742 (
            .O(N__33244),
            .I(N__33229));
    LocalMux I__7741 (
            .O(N__33241),
            .I(N__33226));
    LocalMux I__7740 (
            .O(N__33238),
            .I(N__33223));
    Span4Mux_h I__7739 (
            .O(N__33235),
            .I(N__33218));
    LocalMux I__7738 (
            .O(N__33232),
            .I(N__33218));
    LocalMux I__7737 (
            .O(N__33229),
            .I(N__33215));
    Span4Mux_v I__7736 (
            .O(N__33226),
            .I(N__33212));
    Span4Mux_v I__7735 (
            .O(N__33223),
            .I(N__33207));
    Span4Mux_h I__7734 (
            .O(N__33218),
            .I(N__33207));
    Span4Mux_h I__7733 (
            .O(N__33215),
            .I(N__33200));
    Span4Mux_h I__7732 (
            .O(N__33212),
            .I(N__33200));
    Span4Mux_h I__7731 (
            .O(N__33207),
            .I(N__33200));
    Odrv4 I__7730 (
            .O(N__33200),
            .I(b2v_inst_data_a_escribir_3));
    InMux I__7729 (
            .O(N__33197),
            .I(N__33194));
    LocalMux I__7728 (
            .O(N__33194),
            .I(N__33191));
    Odrv4 I__7727 (
            .O(N__33191),
            .I(N_551_i));
    InMux I__7726 (
            .O(N__33188),
            .I(N__33184));
    InMux I__7725 (
            .O(N__33187),
            .I(N__33181));
    LocalMux I__7724 (
            .O(N__33184),
            .I(N__33177));
    LocalMux I__7723 (
            .O(N__33181),
            .I(N__33174));
    InMux I__7722 (
            .O(N__33180),
            .I(N__33171));
    Span4Mux_v I__7721 (
            .O(N__33177),
            .I(N__33168));
    Span4Mux_h I__7720 (
            .O(N__33174),
            .I(N__33164));
    LocalMux I__7719 (
            .O(N__33171),
            .I(N__33159));
    Sp12to4 I__7718 (
            .O(N__33168),
            .I(N__33159));
    InMux I__7717 (
            .O(N__33167),
            .I(N__33156));
    Span4Mux_h I__7716 (
            .O(N__33164),
            .I(N__33153));
    Odrv12 I__7715 (
            .O(N__33159),
            .I(\b2v_inst.N_481 ));
    LocalMux I__7714 (
            .O(N__33156),
            .I(\b2v_inst.N_481 ));
    Odrv4 I__7713 (
            .O(N__33153),
            .I(\b2v_inst.N_481 ));
    InMux I__7712 (
            .O(N__33146),
            .I(N__33143));
    LocalMux I__7711 (
            .O(N__33143),
            .I(N_121_i));
    CascadeMux I__7710 (
            .O(N__33140),
            .I(N__33136));
    InMux I__7709 (
            .O(N__33139),
            .I(N__33132));
    InMux I__7708 (
            .O(N__33136),
            .I(N__33128));
    InMux I__7707 (
            .O(N__33135),
            .I(N__33125));
    LocalMux I__7706 (
            .O(N__33132),
            .I(N__33121));
    CascadeMux I__7705 (
            .O(N__33131),
            .I(N__33118));
    LocalMux I__7704 (
            .O(N__33128),
            .I(N__33115));
    LocalMux I__7703 (
            .O(N__33125),
            .I(N__33112));
    InMux I__7702 (
            .O(N__33124),
            .I(N__33109));
    Span4Mux_v I__7701 (
            .O(N__33121),
            .I(N__33106));
    InMux I__7700 (
            .O(N__33118),
            .I(N__33103));
    Span4Mux_h I__7699 (
            .O(N__33115),
            .I(N__33100));
    Span4Mux_v I__7698 (
            .O(N__33112),
            .I(N__33097));
    LocalMux I__7697 (
            .O(N__33109),
            .I(N__33094));
    Span4Mux_h I__7696 (
            .O(N__33106),
            .I(N__33089));
    LocalMux I__7695 (
            .O(N__33103),
            .I(N__33089));
    Span4Mux_v I__7694 (
            .O(N__33100),
            .I(N__33084));
    Span4Mux_h I__7693 (
            .O(N__33097),
            .I(N__33084));
    Span12Mux_v I__7692 (
            .O(N__33094),
            .I(N__33081));
    Span4Mux_h I__7691 (
            .O(N__33089),
            .I(N__33078));
    Odrv4 I__7690 (
            .O(N__33084),
            .I(b2v_inst_data_a_escribir_2));
    Odrv12 I__7689 (
            .O(N__33081),
            .I(b2v_inst_data_a_escribir_2));
    Odrv4 I__7688 (
            .O(N__33078),
            .I(b2v_inst_data_a_escribir_2));
    InMux I__7687 (
            .O(N__33071),
            .I(N__33068));
    LocalMux I__7686 (
            .O(N__33068),
            .I(N__33065));
    Odrv4 I__7685 (
            .O(N__33065),
            .I(N_118_i));
    InMux I__7684 (
            .O(N__33062),
            .I(N__33058));
    InMux I__7683 (
            .O(N__33061),
            .I(N__33055));
    LocalMux I__7682 (
            .O(N__33058),
            .I(N__33051));
    LocalMux I__7681 (
            .O(N__33055),
            .I(N__33047));
    InMux I__7680 (
            .O(N__33054),
            .I(N__33044));
    Span4Mux_h I__7679 (
            .O(N__33051),
            .I(N__33041));
    InMux I__7678 (
            .O(N__33050),
            .I(N__33038));
    Span4Mux_h I__7677 (
            .O(N__33047),
            .I(N__33035));
    LocalMux I__7676 (
            .O(N__33044),
            .I(N__33030));
    Span4Mux_h I__7675 (
            .O(N__33041),
            .I(N__33030));
    LocalMux I__7674 (
            .O(N__33038),
            .I(N__33027));
    Odrv4 I__7673 (
            .O(N__33035),
            .I(SYNTHESIZED_WIRE_3_4));
    Odrv4 I__7672 (
            .O(N__33030),
            .I(SYNTHESIZED_WIRE_3_4));
    Odrv4 I__7671 (
            .O(N__33027),
            .I(SYNTHESIZED_WIRE_3_4));
    InMux I__7670 (
            .O(N__33020),
            .I(N__33016));
    InMux I__7669 (
            .O(N__33019),
            .I(N__33011));
    LocalMux I__7668 (
            .O(N__33016),
            .I(N__33007));
    InMux I__7667 (
            .O(N__33015),
            .I(N__33004));
    InMux I__7666 (
            .O(N__33014),
            .I(N__33001));
    LocalMux I__7665 (
            .O(N__33011),
            .I(N__32998));
    CascadeMux I__7664 (
            .O(N__33010),
            .I(N__32995));
    Span4Mux_v I__7663 (
            .O(N__33007),
            .I(N__32992));
    LocalMux I__7662 (
            .O(N__33004),
            .I(N__32989));
    LocalMux I__7661 (
            .O(N__33001),
            .I(N__32986));
    Span4Mux_h I__7660 (
            .O(N__32998),
            .I(N__32983));
    InMux I__7659 (
            .O(N__32995),
            .I(N__32980));
    Span4Mux_h I__7658 (
            .O(N__32992),
            .I(N__32975));
    Span4Mux_h I__7657 (
            .O(N__32989),
            .I(N__32975));
    Odrv12 I__7656 (
            .O(N__32986),
            .I(\b2v_inst.reg_ancho_2Z0Z_4 ));
    Odrv4 I__7655 (
            .O(N__32983),
            .I(\b2v_inst.reg_ancho_2Z0Z_4 ));
    LocalMux I__7654 (
            .O(N__32980),
            .I(\b2v_inst.reg_ancho_2Z0Z_4 ));
    Odrv4 I__7653 (
            .O(N__32975),
            .I(\b2v_inst.reg_ancho_2Z0Z_4 ));
    CEMux I__7652 (
            .O(N__32966),
            .I(N__32960));
    CEMux I__7651 (
            .O(N__32965),
            .I(N__32955));
    CEMux I__7650 (
            .O(N__32964),
            .I(N__32952));
    CEMux I__7649 (
            .O(N__32963),
            .I(N__32949));
    LocalMux I__7648 (
            .O(N__32960),
            .I(N__32946));
    CEMux I__7647 (
            .O(N__32959),
            .I(N__32943));
    CEMux I__7646 (
            .O(N__32958),
            .I(N__32940));
    LocalMux I__7645 (
            .O(N__32955),
            .I(N__32937));
    LocalMux I__7644 (
            .O(N__32952),
            .I(N__32934));
    LocalMux I__7643 (
            .O(N__32949),
            .I(N__32931));
    Span4Mux_v I__7642 (
            .O(N__32946),
            .I(N__32925));
    LocalMux I__7641 (
            .O(N__32943),
            .I(N__32925));
    LocalMux I__7640 (
            .O(N__32940),
            .I(N__32922));
    Span4Mux_v I__7639 (
            .O(N__32937),
            .I(N__32919));
    Span4Mux_v I__7638 (
            .O(N__32934),
            .I(N__32914));
    Span4Mux_h I__7637 (
            .O(N__32931),
            .I(N__32914));
    CEMux I__7636 (
            .O(N__32930),
            .I(N__32911));
    Span4Mux_h I__7635 (
            .O(N__32925),
            .I(N__32900));
    Span4Mux_v I__7634 (
            .O(N__32922),
            .I(N__32900));
    Span4Mux_h I__7633 (
            .O(N__32919),
            .I(N__32900));
    Span4Mux_v I__7632 (
            .O(N__32914),
            .I(N__32900));
    LocalMux I__7631 (
            .O(N__32911),
            .I(N__32900));
    Span4Mux_h I__7630 (
            .O(N__32900),
            .I(N__32893));
    InMux I__7629 (
            .O(N__32899),
            .I(N__32890));
    InMux I__7628 (
            .O(N__32898),
            .I(N__32885));
    InMux I__7627 (
            .O(N__32897),
            .I(N__32885));
    InMux I__7626 (
            .O(N__32896),
            .I(N__32882));
    Odrv4 I__7625 (
            .O(N__32893),
            .I(\b2v_inst.stateZ0Z_23 ));
    LocalMux I__7624 (
            .O(N__32890),
            .I(\b2v_inst.stateZ0Z_23 ));
    LocalMux I__7623 (
            .O(N__32885),
            .I(\b2v_inst.stateZ0Z_23 ));
    LocalMux I__7622 (
            .O(N__32882),
            .I(\b2v_inst.stateZ0Z_23 ));
    CascadeMux I__7621 (
            .O(N__32873),
            .I(N__32869));
    CascadeMux I__7620 (
            .O(N__32872),
            .I(N__32866));
    InMux I__7619 (
            .O(N__32869),
            .I(N__32863));
    InMux I__7618 (
            .O(N__32866),
            .I(N__32860));
    LocalMux I__7617 (
            .O(N__32863),
            .I(N__32854));
    LocalMux I__7616 (
            .O(N__32860),
            .I(N__32854));
    InMux I__7615 (
            .O(N__32859),
            .I(N__32850));
    Span4Mux_h I__7614 (
            .O(N__32854),
            .I(N__32847));
    InMux I__7613 (
            .O(N__32853),
            .I(N__32844));
    LocalMux I__7612 (
            .O(N__32850),
            .I(N__32841));
    Span4Mux_h I__7611 (
            .O(N__32847),
            .I(N__32836));
    LocalMux I__7610 (
            .O(N__32844),
            .I(N__32836));
    Span4Mux_h I__7609 (
            .O(N__32841),
            .I(N__32833));
    Span4Mux_v I__7608 (
            .O(N__32836),
            .I(N__32830));
    Odrv4 I__7607 (
            .O(N__32833),
            .I(b2v_inst_data_a_escribir_9));
    Odrv4 I__7606 (
            .O(N__32830),
            .I(b2v_inst_data_a_escribir_9));
    InMux I__7605 (
            .O(N__32825),
            .I(N__32822));
    LocalMux I__7604 (
            .O(N__32822),
            .I(N_111_i));
    InMux I__7603 (
            .O(N__32819),
            .I(N__32816));
    LocalMux I__7602 (
            .O(N__32816),
            .I(N__32813));
    Span4Mux_h I__7601 (
            .O(N__32813),
            .I(N__32810));
    Span4Mux_h I__7600 (
            .O(N__32810),
            .I(N__32807));
    Span4Mux_h I__7599 (
            .O(N__32807),
            .I(N__32804));
    Odrv4 I__7598 (
            .O(N__32804),
            .I(\b2v_inst.addr_ram_iv_i_1_6 ));
    CascadeMux I__7597 (
            .O(N__32801),
            .I(N__32798));
    InMux I__7596 (
            .O(N__32798),
            .I(N__32795));
    LocalMux I__7595 (
            .O(N__32795),
            .I(N__32792));
    Span12Mux_h I__7594 (
            .O(N__32792),
            .I(N__32789));
    Odrv12 I__7593 (
            .O(N__32789),
            .I(\b2v_inst.addr_ram_iv_i_0_6 ));
    CascadeMux I__7592 (
            .O(N__32786),
            .I(N__32782));
    CascadeMux I__7591 (
            .O(N__32785),
            .I(N__32779));
    CascadeBuf I__7590 (
            .O(N__32782),
            .I(N__32776));
    CascadeBuf I__7589 (
            .O(N__32779),
            .I(N__32773));
    CascadeMux I__7588 (
            .O(N__32776),
            .I(N__32770));
    CascadeMux I__7587 (
            .O(N__32773),
            .I(N__32767));
    CascadeBuf I__7586 (
            .O(N__32770),
            .I(N__32764));
    CascadeBuf I__7585 (
            .O(N__32767),
            .I(N__32761));
    CascadeMux I__7584 (
            .O(N__32764),
            .I(N__32758));
    CascadeMux I__7583 (
            .O(N__32761),
            .I(N__32755));
    CascadeBuf I__7582 (
            .O(N__32758),
            .I(N__32752));
    CascadeBuf I__7581 (
            .O(N__32755),
            .I(N__32749));
    CascadeMux I__7580 (
            .O(N__32752),
            .I(N__32746));
    CascadeMux I__7579 (
            .O(N__32749),
            .I(N__32743));
    CascadeBuf I__7578 (
            .O(N__32746),
            .I(N__32740));
    CascadeBuf I__7577 (
            .O(N__32743),
            .I(N__32737));
    CascadeMux I__7576 (
            .O(N__32740),
            .I(N__32734));
    CascadeMux I__7575 (
            .O(N__32737),
            .I(N__32731));
    CascadeBuf I__7574 (
            .O(N__32734),
            .I(N__32728));
    CascadeBuf I__7573 (
            .O(N__32731),
            .I(N__32725));
    CascadeMux I__7572 (
            .O(N__32728),
            .I(N__32722));
    CascadeMux I__7571 (
            .O(N__32725),
            .I(N__32719));
    InMux I__7570 (
            .O(N__32722),
            .I(N__32716));
    InMux I__7569 (
            .O(N__32719),
            .I(N__32713));
    LocalMux I__7568 (
            .O(N__32716),
            .I(N__32710));
    LocalMux I__7567 (
            .O(N__32713),
            .I(N_298));
    Odrv4 I__7566 (
            .O(N__32710),
            .I(N_298));
    CascadeMux I__7565 (
            .O(N__32705),
            .I(N__32702));
    InMux I__7564 (
            .O(N__32702),
            .I(N__32699));
    LocalMux I__7563 (
            .O(N__32699),
            .I(N__32696));
    Span4Mux_h I__7562 (
            .O(N__32696),
            .I(N__32693));
    Odrv4 I__7561 (
            .O(N__32693),
            .I(SYNTHESIZED_WIRE_1_0));
    CascadeMux I__7560 (
            .O(N__32690),
            .I(N__32687));
    InMux I__7559 (
            .O(N__32687),
            .I(N__32684));
    LocalMux I__7558 (
            .O(N__32684),
            .I(N__32681));
    Odrv12 I__7557 (
            .O(N__32681),
            .I(SYNTHESIZED_WIRE_1_1));
    CascadeMux I__7556 (
            .O(N__32678),
            .I(N__32675));
    InMux I__7555 (
            .O(N__32675),
            .I(N__32672));
    LocalMux I__7554 (
            .O(N__32672),
            .I(N__32669));
    Span4Mux_h I__7553 (
            .O(N__32669),
            .I(N__32666));
    Span4Mux_v I__7552 (
            .O(N__32666),
            .I(N__32663));
    Odrv4 I__7551 (
            .O(N__32663),
            .I(SYNTHESIZED_WIRE_1_4));
    InMux I__7550 (
            .O(N__32660),
            .I(N__32657));
    LocalMux I__7549 (
            .O(N__32657),
            .I(N__32653));
    InMux I__7548 (
            .O(N__32656),
            .I(N__32649));
    Span4Mux_h I__7547 (
            .O(N__32653),
            .I(N__32646));
    InMux I__7546 (
            .O(N__32652),
            .I(N__32643));
    LocalMux I__7545 (
            .O(N__32649),
            .I(b2v_inst_cantidad_temp_2));
    Odrv4 I__7544 (
            .O(N__32646),
            .I(b2v_inst_cantidad_temp_2));
    LocalMux I__7543 (
            .O(N__32643),
            .I(b2v_inst_cantidad_temp_2));
    InMux I__7542 (
            .O(N__32636),
            .I(\b2v_inst.un16_data_ram_cantidad_o_cry_1 ));
    InMux I__7541 (
            .O(N__32633),
            .I(\b2v_inst.un16_data_ram_cantidad_o_cry_2 ));
    InMux I__7540 (
            .O(N__32630),
            .I(N__32627));
    LocalMux I__7539 (
            .O(N__32627),
            .I(N__32624));
    Span4Mux_h I__7538 (
            .O(N__32624),
            .I(N__32620));
    InMux I__7537 (
            .O(N__32623),
            .I(N__32616));
    Span4Mux_h I__7536 (
            .O(N__32620),
            .I(N__32613));
    InMux I__7535 (
            .O(N__32619),
            .I(N__32610));
    LocalMux I__7534 (
            .O(N__32616),
            .I(b2v_inst_cantidad_temp_4));
    Odrv4 I__7533 (
            .O(N__32613),
            .I(b2v_inst_cantidad_temp_4));
    LocalMux I__7532 (
            .O(N__32610),
            .I(b2v_inst_cantidad_temp_4));
    InMux I__7531 (
            .O(N__32603),
            .I(\b2v_inst.un16_data_ram_cantidad_o_cry_3 ));
    CascadeMux I__7530 (
            .O(N__32600),
            .I(N__32596));
    InMux I__7529 (
            .O(N__32599),
            .I(N__32593));
    InMux I__7528 (
            .O(N__32596),
            .I(N__32590));
    LocalMux I__7527 (
            .O(N__32593),
            .I(N__32587));
    LocalMux I__7526 (
            .O(N__32590),
            .I(N__32583));
    Span4Mux_v I__7525 (
            .O(N__32587),
            .I(N__32580));
    InMux I__7524 (
            .O(N__32586),
            .I(N__32577));
    Sp12to4 I__7523 (
            .O(N__32583),
            .I(N__32572));
    Sp12to4 I__7522 (
            .O(N__32580),
            .I(N__32572));
    LocalMux I__7521 (
            .O(N__32577),
            .I(b2v_inst_cantidad_temp_5));
    Odrv12 I__7520 (
            .O(N__32572),
            .I(b2v_inst_cantidad_temp_5));
    InMux I__7519 (
            .O(N__32567),
            .I(\b2v_inst.un16_data_ram_cantidad_o_cry_4 ));
    InMux I__7518 (
            .O(N__32564),
            .I(N__32561));
    LocalMux I__7517 (
            .O(N__32561),
            .I(\b2v_inst.un16_data_ram_cantidad_o_cry_1_c_RNI77COZ0 ));
    InMux I__7516 (
            .O(N__32558),
            .I(N__32555));
    LocalMux I__7515 (
            .O(N__32555),
            .I(N__32552));
    Span4Mux_h I__7514 (
            .O(N__32552),
            .I(N__32549));
    Odrv4 I__7513 (
            .O(N__32549),
            .I(N_553_i));
    InMux I__7512 (
            .O(N__32546),
            .I(N__32530));
    InMux I__7511 (
            .O(N__32545),
            .I(N__32530));
    InMux I__7510 (
            .O(N__32544),
            .I(N__32525));
    InMux I__7509 (
            .O(N__32543),
            .I(N__32525));
    CascadeMux I__7508 (
            .O(N__32542),
            .I(N__32522));
    InMux I__7507 (
            .O(N__32541),
            .I(N__32517));
    InMux I__7506 (
            .O(N__32540),
            .I(N__32517));
    InMux I__7505 (
            .O(N__32539),
            .I(N__32514));
    InMux I__7504 (
            .O(N__32538),
            .I(N__32511));
    InMux I__7503 (
            .O(N__32537),
            .I(N__32506));
    InMux I__7502 (
            .O(N__32536),
            .I(N__32506));
    InMux I__7501 (
            .O(N__32535),
            .I(N__32503));
    LocalMux I__7500 (
            .O(N__32530),
            .I(N__32500));
    LocalMux I__7499 (
            .O(N__32525),
            .I(N__32497));
    InMux I__7498 (
            .O(N__32522),
            .I(N__32494));
    LocalMux I__7497 (
            .O(N__32517),
            .I(N__32485));
    LocalMux I__7496 (
            .O(N__32514),
            .I(N__32485));
    LocalMux I__7495 (
            .O(N__32511),
            .I(N__32485));
    LocalMux I__7494 (
            .O(N__32506),
            .I(N__32485));
    LocalMux I__7493 (
            .O(N__32503),
            .I(N__32482));
    Span4Mux_v I__7492 (
            .O(N__32500),
            .I(N__32477));
    Span4Mux_v I__7491 (
            .O(N__32497),
            .I(N__32477));
    LocalMux I__7490 (
            .O(N__32494),
            .I(N__32474));
    Odrv12 I__7489 (
            .O(N__32485),
            .I(\b2v_inst.un2_valor_max1_THRU_CO ));
    Odrv12 I__7488 (
            .O(N__32482),
            .I(\b2v_inst.un2_valor_max1_THRU_CO ));
    Odrv4 I__7487 (
            .O(N__32477),
            .I(\b2v_inst.un2_valor_max1_THRU_CO ));
    Odrv4 I__7486 (
            .O(N__32474),
            .I(\b2v_inst.un2_valor_max1_THRU_CO ));
    InMux I__7485 (
            .O(N__32465),
            .I(N__32462));
    LocalMux I__7484 (
            .O(N__32462),
            .I(\b2v_inst.data_a_escribir_RNO_2Z0Z_3 ));
    CascadeMux I__7483 (
            .O(N__32459),
            .I(N__32455));
    CascadeMux I__7482 (
            .O(N__32458),
            .I(N__32452));
    InMux I__7481 (
            .O(N__32455),
            .I(N__32449));
    InMux I__7480 (
            .O(N__32452),
            .I(N__32445));
    LocalMux I__7479 (
            .O(N__32449),
            .I(N__32442));
    InMux I__7478 (
            .O(N__32448),
            .I(N__32439));
    LocalMux I__7477 (
            .O(N__32445),
            .I(N__32435));
    Span4Mux_h I__7476 (
            .O(N__32442),
            .I(N__32429));
    LocalMux I__7475 (
            .O(N__32439),
            .I(N__32429));
    InMux I__7474 (
            .O(N__32438),
            .I(N__32426));
    Span4Mux_v I__7473 (
            .O(N__32435),
            .I(N__32423));
    InMux I__7472 (
            .O(N__32434),
            .I(N__32420));
    Span4Mux_v I__7471 (
            .O(N__32429),
            .I(N__32417));
    LocalMux I__7470 (
            .O(N__32426),
            .I(\b2v_inst.reg_ancho_2Z0Z_3 ));
    Odrv4 I__7469 (
            .O(N__32423),
            .I(\b2v_inst.reg_ancho_2Z0Z_3 ));
    LocalMux I__7468 (
            .O(N__32420),
            .I(\b2v_inst.reg_ancho_2Z0Z_3 ));
    Odrv4 I__7467 (
            .O(N__32417),
            .I(\b2v_inst.reg_ancho_2Z0Z_3 ));
    InMux I__7466 (
            .O(N__32408),
            .I(N__32402));
    InMux I__7465 (
            .O(N__32407),
            .I(N__32399));
    InMux I__7464 (
            .O(N__32406),
            .I(N__32386));
    InMux I__7463 (
            .O(N__32405),
            .I(N__32386));
    LocalMux I__7462 (
            .O(N__32402),
            .I(N__32383));
    LocalMux I__7461 (
            .O(N__32399),
            .I(N__32380));
    InMux I__7460 (
            .O(N__32398),
            .I(N__32377));
    InMux I__7459 (
            .O(N__32397),
            .I(N__32374));
    InMux I__7458 (
            .O(N__32396),
            .I(N__32369));
    InMux I__7457 (
            .O(N__32395),
            .I(N__32369));
    InMux I__7456 (
            .O(N__32394),
            .I(N__32366));
    InMux I__7455 (
            .O(N__32393),
            .I(N__32359));
    InMux I__7454 (
            .O(N__32392),
            .I(N__32359));
    InMux I__7453 (
            .O(N__32391),
            .I(N__32359));
    LocalMux I__7452 (
            .O(N__32386),
            .I(N__32350));
    Span4Mux_v I__7451 (
            .O(N__32383),
            .I(N__32350));
    Span4Mux_h I__7450 (
            .O(N__32380),
            .I(N__32350));
    LocalMux I__7449 (
            .O(N__32377),
            .I(N__32350));
    LocalMux I__7448 (
            .O(N__32374),
            .I(N__32344));
    LocalMux I__7447 (
            .O(N__32369),
            .I(N__32344));
    LocalMux I__7446 (
            .O(N__32366),
            .I(N__32341));
    LocalMux I__7445 (
            .O(N__32359),
            .I(N__32336));
    Span4Mux_v I__7444 (
            .O(N__32350),
            .I(N__32336));
    InMux I__7443 (
            .O(N__32349),
            .I(N__32333));
    Odrv12 I__7442 (
            .O(N__32344),
            .I(\b2v_inst.un2_valor_max2_THRU_CO ));
    Odrv4 I__7441 (
            .O(N__32341),
            .I(\b2v_inst.un2_valor_max2_THRU_CO ));
    Odrv4 I__7440 (
            .O(N__32336),
            .I(\b2v_inst.un2_valor_max2_THRU_CO ));
    LocalMux I__7439 (
            .O(N__32333),
            .I(\b2v_inst.un2_valor_max2_THRU_CO ));
    CascadeMux I__7438 (
            .O(N__32324),
            .I(N__32321));
    InMux I__7437 (
            .O(N__32321),
            .I(N__32318));
    LocalMux I__7436 (
            .O(N__32318),
            .I(N__32315));
    Span4Mux_h I__7435 (
            .O(N__32315),
            .I(N__32312));
    Odrv4 I__7434 (
            .O(N__32312),
            .I(\b2v_inst.N_264 ));
    InMux I__7433 (
            .O(N__32309),
            .I(N__32306));
    LocalMux I__7432 (
            .O(N__32306),
            .I(N__32302));
    InMux I__7431 (
            .O(N__32305),
            .I(N__32298));
    Span4Mux_h I__7430 (
            .O(N__32302),
            .I(N__32295));
    InMux I__7429 (
            .O(N__32301),
            .I(N__32292));
    LocalMux I__7428 (
            .O(N__32298),
            .I(\b2v_inst.reg_ancho_3Z0Z_10 ));
    Odrv4 I__7427 (
            .O(N__32295),
            .I(\b2v_inst.reg_ancho_3Z0Z_10 ));
    LocalMux I__7426 (
            .O(N__32292),
            .I(\b2v_inst.reg_ancho_3Z0Z_10 ));
    InMux I__7425 (
            .O(N__32285),
            .I(N__32279));
    InMux I__7424 (
            .O(N__32284),
            .I(N__32276));
    InMux I__7423 (
            .O(N__32283),
            .I(N__32273));
    InMux I__7422 (
            .O(N__32282),
            .I(N__32270));
    LocalMux I__7421 (
            .O(N__32279),
            .I(N__32267));
    LocalMux I__7420 (
            .O(N__32276),
            .I(N__32264));
    LocalMux I__7419 (
            .O(N__32273),
            .I(N__32261));
    LocalMux I__7418 (
            .O(N__32270),
            .I(N__32258));
    Span4Mux_h I__7417 (
            .O(N__32267),
            .I(N__32255));
    Span4Mux_h I__7416 (
            .O(N__32264),
            .I(N__32252));
    Span4Mux_h I__7415 (
            .O(N__32261),
            .I(N__32249));
    Span4Mux_h I__7414 (
            .O(N__32258),
            .I(N__32246));
    Span4Mux_h I__7413 (
            .O(N__32255),
            .I(N__32241));
    Span4Mux_v I__7412 (
            .O(N__32252),
            .I(N__32241));
    Span4Mux_v I__7411 (
            .O(N__32249),
            .I(N__32236));
    Span4Mux_h I__7410 (
            .O(N__32246),
            .I(N__32236));
    Odrv4 I__7409 (
            .O(N__32241),
            .I(SYNTHESIZED_WIRE_3_3));
    Odrv4 I__7408 (
            .O(N__32236),
            .I(SYNTHESIZED_WIRE_3_3));
    InMux I__7407 (
            .O(N__32231),
            .I(N__32226));
    InMux I__7406 (
            .O(N__32230),
            .I(N__32223));
    InMux I__7405 (
            .O(N__32229),
            .I(N__32220));
    LocalMux I__7404 (
            .O(N__32226),
            .I(N__32215));
    LocalMux I__7403 (
            .O(N__32223),
            .I(N__32215));
    LocalMux I__7402 (
            .O(N__32220),
            .I(\b2v_inst.reg_ancho_3Z0Z_3 ));
    Odrv4 I__7401 (
            .O(N__32215),
            .I(\b2v_inst.reg_ancho_3Z0Z_3 ));
    InMux I__7400 (
            .O(N__32210),
            .I(N__32206));
    InMux I__7399 (
            .O(N__32209),
            .I(N__32201));
    LocalMux I__7398 (
            .O(N__32206),
            .I(N__32198));
    InMux I__7397 (
            .O(N__32205),
            .I(N__32195));
    InMux I__7396 (
            .O(N__32204),
            .I(N__32192));
    LocalMux I__7395 (
            .O(N__32201),
            .I(N__32189));
    Span4Mux_h I__7394 (
            .O(N__32198),
            .I(N__32186));
    LocalMux I__7393 (
            .O(N__32195),
            .I(N__32183));
    LocalMux I__7392 (
            .O(N__32192),
            .I(N__32180));
    Span4Mux_v I__7391 (
            .O(N__32189),
            .I(N__32177));
    Span4Mux_h I__7390 (
            .O(N__32186),
            .I(N__32172));
    Span4Mux_h I__7389 (
            .O(N__32183),
            .I(N__32172));
    Span4Mux_v I__7388 (
            .O(N__32180),
            .I(N__32169));
    Span4Mux_v I__7387 (
            .O(N__32177),
            .I(N__32166));
    Span4Mux_v I__7386 (
            .O(N__32172),
            .I(N__32163));
    Span4Mux_h I__7385 (
            .O(N__32169),
            .I(N__32160));
    Odrv4 I__7384 (
            .O(N__32166),
            .I(SYNTHESIZED_WIRE_3_2));
    Odrv4 I__7383 (
            .O(N__32163),
            .I(SYNTHESIZED_WIRE_3_2));
    Odrv4 I__7382 (
            .O(N__32160),
            .I(SYNTHESIZED_WIRE_3_2));
    InMux I__7381 (
            .O(N__32153),
            .I(N__32148));
    InMux I__7380 (
            .O(N__32152),
            .I(N__32145));
    InMux I__7379 (
            .O(N__32151),
            .I(N__32142));
    LocalMux I__7378 (
            .O(N__32148),
            .I(N__32139));
    LocalMux I__7377 (
            .O(N__32145),
            .I(\b2v_inst.reg_ancho_3Z0Z_2 ));
    LocalMux I__7376 (
            .O(N__32142),
            .I(\b2v_inst.reg_ancho_3Z0Z_2 ));
    Odrv4 I__7375 (
            .O(N__32139),
            .I(\b2v_inst.reg_ancho_3Z0Z_2 ));
    InMux I__7374 (
            .O(N__32132),
            .I(N__32128));
    InMux I__7373 (
            .O(N__32131),
            .I(N__32125));
    LocalMux I__7372 (
            .O(N__32128),
            .I(N__32121));
    LocalMux I__7371 (
            .O(N__32125),
            .I(N__32118));
    InMux I__7370 (
            .O(N__32124),
            .I(N__32114));
    Span4Mux_h I__7369 (
            .O(N__32121),
            .I(N__32111));
    Span4Mux_v I__7368 (
            .O(N__32118),
            .I(N__32108));
    InMux I__7367 (
            .O(N__32117),
            .I(N__32105));
    LocalMux I__7366 (
            .O(N__32114),
            .I(N__32102));
    Span4Mux_h I__7365 (
            .O(N__32111),
            .I(N__32099));
    Span4Mux_v I__7364 (
            .O(N__32108),
            .I(N__32096));
    LocalMux I__7363 (
            .O(N__32105),
            .I(N__32093));
    Odrv12 I__7362 (
            .O(N__32102),
            .I(SYNTHESIZED_WIRE_3_5));
    Odrv4 I__7361 (
            .O(N__32099),
            .I(SYNTHESIZED_WIRE_3_5));
    Odrv4 I__7360 (
            .O(N__32096),
            .I(SYNTHESIZED_WIRE_3_5));
    Odrv4 I__7359 (
            .O(N__32093),
            .I(SYNTHESIZED_WIRE_3_5));
    CascadeMux I__7358 (
            .O(N__32084),
            .I(N__32079));
    InMux I__7357 (
            .O(N__32083),
            .I(N__32076));
    InMux I__7356 (
            .O(N__32082),
            .I(N__32073));
    InMux I__7355 (
            .O(N__32079),
            .I(N__32070));
    LocalMux I__7354 (
            .O(N__32076),
            .I(N__32065));
    LocalMux I__7353 (
            .O(N__32073),
            .I(N__32065));
    LocalMux I__7352 (
            .O(N__32070),
            .I(\b2v_inst.reg_ancho_3Z0Z_5 ));
    Odrv4 I__7351 (
            .O(N__32065),
            .I(\b2v_inst.reg_ancho_3Z0Z_5 ));
    CEMux I__7350 (
            .O(N__32060),
            .I(N__32056));
    CEMux I__7349 (
            .O(N__32059),
            .I(N__32053));
    LocalMux I__7348 (
            .O(N__32056),
            .I(N__32048));
    LocalMux I__7347 (
            .O(N__32053),
            .I(N__32045));
    CEMux I__7346 (
            .O(N__32052),
            .I(N__32042));
    InMux I__7345 (
            .O(N__32051),
            .I(N__32039));
    Span4Mux_v I__7344 (
            .O(N__32048),
            .I(N__32036));
    Span4Mux_v I__7343 (
            .O(N__32045),
            .I(N__32033));
    LocalMux I__7342 (
            .O(N__32042),
            .I(N__32030));
    LocalMux I__7341 (
            .O(N__32039),
            .I(N__32027));
    Span4Mux_h I__7340 (
            .O(N__32036),
            .I(N__32021));
    Span4Mux_h I__7339 (
            .O(N__32033),
            .I(N__32016));
    Span4Mux_h I__7338 (
            .O(N__32030),
            .I(N__32016));
    Span4Mux_h I__7337 (
            .O(N__32027),
            .I(N__32013));
    InMux I__7336 (
            .O(N__32026),
            .I(N__32008));
    InMux I__7335 (
            .O(N__32025),
            .I(N__32008));
    InMux I__7334 (
            .O(N__32024),
            .I(N__32005));
    Odrv4 I__7333 (
            .O(N__32021),
            .I(\b2v_inst.stateZ0Z_21 ));
    Odrv4 I__7332 (
            .O(N__32016),
            .I(\b2v_inst.stateZ0Z_21 ));
    Odrv4 I__7331 (
            .O(N__32013),
            .I(\b2v_inst.stateZ0Z_21 ));
    LocalMux I__7330 (
            .O(N__32008),
            .I(\b2v_inst.stateZ0Z_21 ));
    LocalMux I__7329 (
            .O(N__32005),
            .I(\b2v_inst.stateZ0Z_21 ));
    InMux I__7328 (
            .O(N__31994),
            .I(N__31990));
    InMux I__7327 (
            .O(N__31993),
            .I(N__31986));
    LocalMux I__7326 (
            .O(N__31990),
            .I(N__31982));
    InMux I__7325 (
            .O(N__31989),
            .I(N__31979));
    LocalMux I__7324 (
            .O(N__31986),
            .I(N__31976));
    InMux I__7323 (
            .O(N__31985),
            .I(N__31973));
    Span4Mux_h I__7322 (
            .O(N__31982),
            .I(N__31966));
    LocalMux I__7321 (
            .O(N__31979),
            .I(N__31966));
    Span4Mux_v I__7320 (
            .O(N__31976),
            .I(N__31966));
    LocalMux I__7319 (
            .O(N__31973),
            .I(N__31963));
    Span4Mux_h I__7318 (
            .O(N__31966),
            .I(N__31958));
    Span4Mux_h I__7317 (
            .O(N__31963),
            .I(N__31958));
    Odrv4 I__7316 (
            .O(N__31958),
            .I(SYNTHESIZED_WIRE_3_9));
    InMux I__7315 (
            .O(N__31955),
            .I(N__31951));
    InMux I__7314 (
            .O(N__31954),
            .I(N__31947));
    LocalMux I__7313 (
            .O(N__31951),
            .I(N__31943));
    InMux I__7312 (
            .O(N__31950),
            .I(N__31940));
    LocalMux I__7311 (
            .O(N__31947),
            .I(N__31937));
    InMux I__7310 (
            .O(N__31946),
            .I(N__31934));
    Span4Mux_h I__7309 (
            .O(N__31943),
            .I(N__31931));
    LocalMux I__7308 (
            .O(N__31940),
            .I(N__31928));
    Odrv12 I__7307 (
            .O(N__31937),
            .I(\b2v_inst.reg_anteriorZ0Z_9 ));
    LocalMux I__7306 (
            .O(N__31934),
            .I(\b2v_inst.reg_anteriorZ0Z_9 ));
    Odrv4 I__7305 (
            .O(N__31931),
            .I(\b2v_inst.reg_anteriorZ0Z_9 ));
    Odrv4 I__7304 (
            .O(N__31928),
            .I(\b2v_inst.reg_anteriorZ0Z_9 ));
    InMux I__7303 (
            .O(N__31919),
            .I(N__31914));
    InMux I__7302 (
            .O(N__31918),
            .I(N__31909));
    InMux I__7301 (
            .O(N__31917),
            .I(N__31909));
    LocalMux I__7300 (
            .O(N__31914),
            .I(N__31889));
    LocalMux I__7299 (
            .O(N__31909),
            .I(N__31889));
    InMux I__7298 (
            .O(N__31908),
            .I(N__31876));
    InMux I__7297 (
            .O(N__31907),
            .I(N__31876));
    InMux I__7296 (
            .O(N__31906),
            .I(N__31876));
    InMux I__7295 (
            .O(N__31905),
            .I(N__31876));
    InMux I__7294 (
            .O(N__31904),
            .I(N__31876));
    InMux I__7293 (
            .O(N__31903),
            .I(N__31876));
    InMux I__7292 (
            .O(N__31902),
            .I(N__31873));
    InMux I__7291 (
            .O(N__31901),
            .I(N__31864));
    InMux I__7290 (
            .O(N__31900),
            .I(N__31864));
    InMux I__7289 (
            .O(N__31899),
            .I(N__31864));
    InMux I__7288 (
            .O(N__31898),
            .I(N__31864));
    InMux I__7287 (
            .O(N__31897),
            .I(N__31859));
    InMux I__7286 (
            .O(N__31896),
            .I(N__31859));
    InMux I__7285 (
            .O(N__31895),
            .I(N__31853));
    InMux I__7284 (
            .O(N__31894),
            .I(N__31853));
    Span4Mux_v I__7283 (
            .O(N__31889),
            .I(N__31848));
    LocalMux I__7282 (
            .O(N__31876),
            .I(N__31848));
    LocalMux I__7281 (
            .O(N__31873),
            .I(N__31843));
    LocalMux I__7280 (
            .O(N__31864),
            .I(N__31843));
    LocalMux I__7279 (
            .O(N__31859),
            .I(N__31840));
    InMux I__7278 (
            .O(N__31858),
            .I(N__31837));
    LocalMux I__7277 (
            .O(N__31853),
            .I(N__31834));
    Span4Mux_h I__7276 (
            .O(N__31848),
            .I(N__31828));
    Span4Mux_v I__7275 (
            .O(N__31843),
            .I(N__31825));
    Span4Mux_h I__7274 (
            .O(N__31840),
            .I(N__31820));
    LocalMux I__7273 (
            .O(N__31837),
            .I(N__31820));
    Span4Mux_v I__7272 (
            .O(N__31834),
            .I(N__31817));
    InMux I__7271 (
            .O(N__31833),
            .I(N__31814));
    InMux I__7270 (
            .O(N__31832),
            .I(N__31809));
    InMux I__7269 (
            .O(N__31831),
            .I(N__31809));
    Span4Mux_v I__7268 (
            .O(N__31828),
            .I(N__31802));
    Span4Mux_h I__7267 (
            .O(N__31825),
            .I(N__31802));
    Span4Mux_h I__7266 (
            .O(N__31820),
            .I(N__31802));
    Sp12to4 I__7265 (
            .O(N__31817),
            .I(N__31795));
    LocalMux I__7264 (
            .O(N__31814),
            .I(N__31795));
    LocalMux I__7263 (
            .O(N__31809),
            .I(N__31795));
    Span4Mux_h I__7262 (
            .O(N__31802),
            .I(N__31792));
    Span12Mux_h I__7261 (
            .O(N__31795),
            .I(N__31789));
    Span4Mux_h I__7260 (
            .O(N__31792),
            .I(N__31786));
    Odrv12 I__7259 (
            .O(N__31789),
            .I(\b2v_inst.ignorar_anteriorZ0 ));
    Odrv4 I__7258 (
            .O(N__31786),
            .I(\b2v_inst.ignorar_anteriorZ0 ));
    InMux I__7257 (
            .O(N__31781),
            .I(N__31777));
    InMux I__7256 (
            .O(N__31780),
            .I(N__31773));
    LocalMux I__7255 (
            .O(N__31777),
            .I(N__31769));
    InMux I__7254 (
            .O(N__31776),
            .I(N__31766));
    LocalMux I__7253 (
            .O(N__31773),
            .I(N__31763));
    InMux I__7252 (
            .O(N__31772),
            .I(N__31760));
    Span4Mux_v I__7251 (
            .O(N__31769),
            .I(N__31757));
    LocalMux I__7250 (
            .O(N__31766),
            .I(N__31754));
    Span4Mux_h I__7249 (
            .O(N__31763),
            .I(N__31751));
    LocalMux I__7248 (
            .O(N__31760),
            .I(N__31748));
    Span4Mux_h I__7247 (
            .O(N__31757),
            .I(N__31745));
    Span4Mux_h I__7246 (
            .O(N__31754),
            .I(N__31742));
    Span4Mux_v I__7245 (
            .O(N__31751),
            .I(N__31737));
    Span4Mux_h I__7244 (
            .O(N__31748),
            .I(N__31737));
    Odrv4 I__7243 (
            .O(N__31745),
            .I(SYNTHESIZED_WIRE_3_10));
    Odrv4 I__7242 (
            .O(N__31742),
            .I(SYNTHESIZED_WIRE_3_10));
    Odrv4 I__7241 (
            .O(N__31737),
            .I(SYNTHESIZED_WIRE_3_10));
    CascadeMux I__7240 (
            .O(N__31730),
            .I(N__31727));
    InMux I__7239 (
            .O(N__31727),
            .I(N__31723));
    InMux I__7238 (
            .O(N__31726),
            .I(N__31720));
    LocalMux I__7237 (
            .O(N__31723),
            .I(N__31715));
    LocalMux I__7236 (
            .O(N__31720),
            .I(N__31712));
    InMux I__7235 (
            .O(N__31719),
            .I(N__31709));
    InMux I__7234 (
            .O(N__31718),
            .I(N__31706));
    Span4Mux_v I__7233 (
            .O(N__31715),
            .I(N__31703));
    Span4Mux_h I__7232 (
            .O(N__31712),
            .I(N__31700));
    LocalMux I__7231 (
            .O(N__31709),
            .I(N__31697));
    LocalMux I__7230 (
            .O(N__31706),
            .I(\b2v_inst.reg_anteriorZ0Z_10 ));
    Odrv4 I__7229 (
            .O(N__31703),
            .I(\b2v_inst.reg_anteriorZ0Z_10 ));
    Odrv4 I__7228 (
            .O(N__31700),
            .I(\b2v_inst.reg_anteriorZ0Z_10 ));
    Odrv4 I__7227 (
            .O(N__31697),
            .I(\b2v_inst.reg_anteriorZ0Z_10 ));
    CEMux I__7226 (
            .O(N__31688),
            .I(N__31683));
    CEMux I__7225 (
            .O(N__31687),
            .I(N__31680));
    CEMux I__7224 (
            .O(N__31686),
            .I(N__31677));
    LocalMux I__7223 (
            .O(N__31683),
            .I(N__31674));
    LocalMux I__7222 (
            .O(N__31680),
            .I(N__31668));
    LocalMux I__7221 (
            .O(N__31677),
            .I(N__31663));
    Span4Mux_v I__7220 (
            .O(N__31674),
            .I(N__31660));
    CEMux I__7219 (
            .O(N__31673),
            .I(N__31657));
    CEMux I__7218 (
            .O(N__31672),
            .I(N__31654));
    CEMux I__7217 (
            .O(N__31671),
            .I(N__31651));
    Span4Mux_h I__7216 (
            .O(N__31668),
            .I(N__31648));
    CascadeMux I__7215 (
            .O(N__31667),
            .I(N__31645));
    InMux I__7214 (
            .O(N__31666),
            .I(N__31642));
    Span4Mux_v I__7213 (
            .O(N__31663),
            .I(N__31639));
    Span4Mux_v I__7212 (
            .O(N__31660),
            .I(N__31634));
    LocalMux I__7211 (
            .O(N__31657),
            .I(N__31634));
    LocalMux I__7210 (
            .O(N__31654),
            .I(N__31631));
    LocalMux I__7209 (
            .O(N__31651),
            .I(N__31626));
    Span4Mux_v I__7208 (
            .O(N__31648),
            .I(N__31626));
    InMux I__7207 (
            .O(N__31645),
            .I(N__31623));
    LocalMux I__7206 (
            .O(N__31642),
            .I(N__31619));
    Sp12to4 I__7205 (
            .O(N__31639),
            .I(N__31614));
    Sp12to4 I__7204 (
            .O(N__31634),
            .I(N__31614));
    Span4Mux_v I__7203 (
            .O(N__31631),
            .I(N__31610));
    Span4Mux_h I__7202 (
            .O(N__31626),
            .I(N__31605));
    LocalMux I__7201 (
            .O(N__31623),
            .I(N__31605));
    InMux I__7200 (
            .O(N__31622),
            .I(N__31601));
    Span4Mux_h I__7199 (
            .O(N__31619),
            .I(N__31598));
    Span12Mux_h I__7198 (
            .O(N__31614),
            .I(N__31595));
    InMux I__7197 (
            .O(N__31613),
            .I(N__31592));
    Span4Mux_h I__7196 (
            .O(N__31610),
            .I(N__31587));
    Span4Mux_v I__7195 (
            .O(N__31605),
            .I(N__31587));
    InMux I__7194 (
            .O(N__31604),
            .I(N__31584));
    LocalMux I__7193 (
            .O(N__31601),
            .I(\b2v_inst.stateZ0Z_27 ));
    Odrv4 I__7192 (
            .O(N__31598),
            .I(\b2v_inst.stateZ0Z_27 ));
    Odrv12 I__7191 (
            .O(N__31595),
            .I(\b2v_inst.stateZ0Z_27 ));
    LocalMux I__7190 (
            .O(N__31592),
            .I(\b2v_inst.stateZ0Z_27 ));
    Odrv4 I__7189 (
            .O(N__31587),
            .I(\b2v_inst.stateZ0Z_27 ));
    LocalMux I__7188 (
            .O(N__31584),
            .I(\b2v_inst.stateZ0Z_27 ));
    InMux I__7187 (
            .O(N__31571),
            .I(N__31567));
    InMux I__7186 (
            .O(N__31570),
            .I(N__31564));
    LocalMux I__7185 (
            .O(N__31567),
            .I(N__31559));
    LocalMux I__7184 (
            .O(N__31564),
            .I(N__31556));
    InMux I__7183 (
            .O(N__31563),
            .I(N__31553));
    InMux I__7182 (
            .O(N__31562),
            .I(N__31550));
    Span4Mux_h I__7181 (
            .O(N__31559),
            .I(N__31543));
    Span4Mux_v I__7180 (
            .O(N__31556),
            .I(N__31543));
    LocalMux I__7179 (
            .O(N__31553),
            .I(N__31543));
    LocalMux I__7178 (
            .O(N__31550),
            .I(N__31540));
    Span4Mux_h I__7177 (
            .O(N__31543),
            .I(N__31537));
    Span4Mux_h I__7176 (
            .O(N__31540),
            .I(N__31534));
    Odrv4 I__7175 (
            .O(N__31537),
            .I(SYNTHESIZED_WIRE_3_6));
    Odrv4 I__7174 (
            .O(N__31534),
            .I(SYNTHESIZED_WIRE_3_6));
    CascadeMux I__7173 (
            .O(N__31529),
            .I(N__31526));
    InMux I__7172 (
            .O(N__31526),
            .I(N__31522));
    InMux I__7171 (
            .O(N__31525),
            .I(N__31519));
    LocalMux I__7170 (
            .O(N__31522),
            .I(N__31515));
    LocalMux I__7169 (
            .O(N__31519),
            .I(N__31511));
    InMux I__7168 (
            .O(N__31518),
            .I(N__31508));
    Span4Mux_h I__7167 (
            .O(N__31515),
            .I(N__31505));
    InMux I__7166 (
            .O(N__31514),
            .I(N__31502));
    Span4Mux_v I__7165 (
            .O(N__31511),
            .I(N__31499));
    LocalMux I__7164 (
            .O(N__31508),
            .I(\b2v_inst.reg_anteriorZ0Z_6 ));
    Odrv4 I__7163 (
            .O(N__31505),
            .I(\b2v_inst.reg_anteriorZ0Z_6 ));
    LocalMux I__7162 (
            .O(N__31502),
            .I(\b2v_inst.reg_anteriorZ0Z_6 ));
    Odrv4 I__7161 (
            .O(N__31499),
            .I(\b2v_inst.reg_anteriorZ0Z_6 ));
    InMux I__7160 (
            .O(N__31490),
            .I(N__31484));
    InMux I__7159 (
            .O(N__31489),
            .I(N__31480));
    CascadeMux I__7158 (
            .O(N__31488),
            .I(N__31477));
    InMux I__7157 (
            .O(N__31487),
            .I(N__31474));
    LocalMux I__7156 (
            .O(N__31484),
            .I(N__31471));
    InMux I__7155 (
            .O(N__31483),
            .I(N__31468));
    LocalMux I__7154 (
            .O(N__31480),
            .I(N__31465));
    InMux I__7153 (
            .O(N__31477),
            .I(N__31462));
    LocalMux I__7152 (
            .O(N__31474),
            .I(N__31459));
    Span4Mux_h I__7151 (
            .O(N__31471),
            .I(N__31450));
    LocalMux I__7150 (
            .O(N__31468),
            .I(N__31450));
    Span4Mux_v I__7149 (
            .O(N__31465),
            .I(N__31450));
    LocalMux I__7148 (
            .O(N__31462),
            .I(N__31450));
    Span4Mux_h I__7147 (
            .O(N__31459),
            .I(N__31445));
    Span4Mux_v I__7146 (
            .O(N__31450),
            .I(N__31445));
    Odrv4 I__7145 (
            .O(N__31445),
            .I(\b2v_inst.reg_ancho_2Z0Z_10 ));
    InMux I__7144 (
            .O(N__31442),
            .I(N__31439));
    LocalMux I__7143 (
            .O(N__31439),
            .I(N__31435));
    InMux I__7142 (
            .O(N__31438),
            .I(N__31432));
    Span4Mux_v I__7141 (
            .O(N__31435),
            .I(N__31427));
    LocalMux I__7140 (
            .O(N__31432),
            .I(N__31427));
    Span4Mux_h I__7139 (
            .O(N__31427),
            .I(N__31423));
    InMux I__7138 (
            .O(N__31426),
            .I(N__31420));
    Odrv4 I__7137 (
            .O(N__31423),
            .I(\b2v_inst.reg_ancho_3Z0Z_4 ));
    LocalMux I__7136 (
            .O(N__31420),
            .I(\b2v_inst.reg_ancho_3Z0Z_4 ));
    InMux I__7135 (
            .O(N__31415),
            .I(N__31412));
    LocalMux I__7134 (
            .O(N__31412),
            .I(N__31409));
    Span4Mux_v I__7133 (
            .O(N__31409),
            .I(N__31406));
    Span4Mux_h I__7132 (
            .O(N__31406),
            .I(N__31403));
    Odrv4 I__7131 (
            .O(N__31403),
            .I(\b2v_inst.data_a_escribir11_3_and ));
    InMux I__7130 (
            .O(N__31400),
            .I(N__31397));
    LocalMux I__7129 (
            .O(N__31397),
            .I(N__31391));
    InMux I__7128 (
            .O(N__31396),
            .I(N__31388));
    InMux I__7127 (
            .O(N__31395),
            .I(N__31385));
    InMux I__7126 (
            .O(N__31394),
            .I(N__31382));
    Span4Mux_v I__7125 (
            .O(N__31391),
            .I(N__31377));
    LocalMux I__7124 (
            .O(N__31388),
            .I(N__31377));
    LocalMux I__7123 (
            .O(N__31385),
            .I(N__31374));
    LocalMux I__7122 (
            .O(N__31382),
            .I(N__31371));
    Span4Mux_v I__7121 (
            .O(N__31377),
            .I(N__31368));
    Span4Mux_v I__7120 (
            .O(N__31374),
            .I(N__31363));
    Span4Mux_h I__7119 (
            .O(N__31371),
            .I(N__31363));
    Span4Mux_h I__7118 (
            .O(N__31368),
            .I(N__31360));
    Span4Mux_v I__7117 (
            .O(N__31363),
            .I(N__31357));
    Odrv4 I__7116 (
            .O(N__31360),
            .I(SYNTHESIZED_WIRE_3_1));
    Odrv4 I__7115 (
            .O(N__31357),
            .I(SYNTHESIZED_WIRE_3_1));
    CascadeMux I__7114 (
            .O(N__31352),
            .I(N__31347));
    InMux I__7113 (
            .O(N__31351),
            .I(N__31343));
    InMux I__7112 (
            .O(N__31350),
            .I(N__31340));
    InMux I__7111 (
            .O(N__31347),
            .I(N__31337));
    InMux I__7110 (
            .O(N__31346),
            .I(N__31334));
    LocalMux I__7109 (
            .O(N__31343),
            .I(N__31331));
    LocalMux I__7108 (
            .O(N__31340),
            .I(N__31327));
    LocalMux I__7107 (
            .O(N__31337),
            .I(N__31322));
    LocalMux I__7106 (
            .O(N__31334),
            .I(N__31322));
    Span4Mux_h I__7105 (
            .O(N__31331),
            .I(N__31319));
    InMux I__7104 (
            .O(N__31330),
            .I(N__31316));
    Span4Mux_v I__7103 (
            .O(N__31327),
            .I(N__31311));
    Span4Mux_v I__7102 (
            .O(N__31322),
            .I(N__31311));
    Odrv4 I__7101 (
            .O(N__31319),
            .I(\b2v_inst.reg_ancho_2Z0Z_1 ));
    LocalMux I__7100 (
            .O(N__31316),
            .I(\b2v_inst.reg_ancho_2Z0Z_1 ));
    Odrv4 I__7099 (
            .O(N__31311),
            .I(\b2v_inst.reg_ancho_2Z0Z_1 ));
    CascadeMux I__7098 (
            .O(N__31304),
            .I(N__31301));
    InMux I__7097 (
            .O(N__31301),
            .I(N__31296));
    InMux I__7096 (
            .O(N__31300),
            .I(N__31293));
    InMux I__7095 (
            .O(N__31299),
            .I(N__31290));
    LocalMux I__7094 (
            .O(N__31296),
            .I(N__31287));
    LocalMux I__7093 (
            .O(N__31293),
            .I(N__31284));
    LocalMux I__7092 (
            .O(N__31290),
            .I(N__31279));
    Span4Mux_h I__7091 (
            .O(N__31287),
            .I(N__31276));
    Span4Mux_h I__7090 (
            .O(N__31284),
            .I(N__31273));
    InMux I__7089 (
            .O(N__31283),
            .I(N__31268));
    InMux I__7088 (
            .O(N__31282),
            .I(N__31268));
    Span4Mux_h I__7087 (
            .O(N__31279),
            .I(N__31265));
    Odrv4 I__7086 (
            .O(N__31276),
            .I(\b2v_inst.reg_ancho_2Z0Z_2 ));
    Odrv4 I__7085 (
            .O(N__31273),
            .I(\b2v_inst.reg_ancho_2Z0Z_2 ));
    LocalMux I__7084 (
            .O(N__31268),
            .I(\b2v_inst.reg_ancho_2Z0Z_2 ));
    Odrv4 I__7083 (
            .O(N__31265),
            .I(\b2v_inst.reg_ancho_2Z0Z_2 ));
    InMux I__7082 (
            .O(N__31256),
            .I(N__31252));
    InMux I__7081 (
            .O(N__31255),
            .I(N__31249));
    LocalMux I__7080 (
            .O(N__31252),
            .I(N__31246));
    LocalMux I__7079 (
            .O(N__31249),
            .I(N__31242));
    Span4Mux_v I__7078 (
            .O(N__31246),
            .I(N__31238));
    InMux I__7077 (
            .O(N__31245),
            .I(N__31235));
    Span4Mux_v I__7076 (
            .O(N__31242),
            .I(N__31232));
    InMux I__7075 (
            .O(N__31241),
            .I(N__31229));
    Span4Mux_h I__7074 (
            .O(N__31238),
            .I(N__31224));
    LocalMux I__7073 (
            .O(N__31235),
            .I(N__31224));
    Span4Mux_h I__7072 (
            .O(N__31232),
            .I(N__31220));
    LocalMux I__7071 (
            .O(N__31229),
            .I(N__31217));
    Span4Mux_h I__7070 (
            .O(N__31224),
            .I(N__31214));
    InMux I__7069 (
            .O(N__31223),
            .I(N__31211));
    Odrv4 I__7068 (
            .O(N__31220),
            .I(\b2v_inst.reg_ancho_1Z0Z_2 ));
    Odrv12 I__7067 (
            .O(N__31217),
            .I(\b2v_inst.reg_ancho_1Z0Z_2 ));
    Odrv4 I__7066 (
            .O(N__31214),
            .I(\b2v_inst.reg_ancho_1Z0Z_2 ));
    LocalMux I__7065 (
            .O(N__31211),
            .I(\b2v_inst.reg_ancho_1Z0Z_2 ));
    InMux I__7064 (
            .O(N__31202),
            .I(N__31199));
    LocalMux I__7063 (
            .O(N__31199),
            .I(N__31196));
    Span4Mux_h I__7062 (
            .O(N__31196),
            .I(N__31192));
    InMux I__7061 (
            .O(N__31195),
            .I(N__31189));
    Odrv4 I__7060 (
            .O(N__31192),
            .I(\b2v_inst.eventosZ0Z_2 ));
    LocalMux I__7059 (
            .O(N__31189),
            .I(\b2v_inst.eventosZ0Z_2 ));
    CascadeMux I__7058 (
            .O(N__31184),
            .I(\b2v_inst.data_a_escribir_RNO_2Z0Z_2_cascade_ ));
    InMux I__7057 (
            .O(N__31181),
            .I(N__31161));
    InMux I__7056 (
            .O(N__31180),
            .I(N__31158));
    InMux I__7055 (
            .O(N__31179),
            .I(N__31151));
    InMux I__7054 (
            .O(N__31178),
            .I(N__31151));
    InMux I__7053 (
            .O(N__31177),
            .I(N__31151));
    InMux I__7052 (
            .O(N__31176),
            .I(N__31148));
    InMux I__7051 (
            .O(N__31175),
            .I(N__31139));
    InMux I__7050 (
            .O(N__31174),
            .I(N__31139));
    InMux I__7049 (
            .O(N__31173),
            .I(N__31139));
    InMux I__7048 (
            .O(N__31172),
            .I(N__31139));
    InMux I__7047 (
            .O(N__31171),
            .I(N__31130));
    InMux I__7046 (
            .O(N__31170),
            .I(N__31130));
    InMux I__7045 (
            .O(N__31169),
            .I(N__31130));
    InMux I__7044 (
            .O(N__31168),
            .I(N__31130));
    InMux I__7043 (
            .O(N__31167),
            .I(N__31120));
    InMux I__7042 (
            .O(N__31166),
            .I(N__31120));
    InMux I__7041 (
            .O(N__31165),
            .I(N__31120));
    InMux I__7040 (
            .O(N__31164),
            .I(N__31120));
    LocalMux I__7039 (
            .O(N__31161),
            .I(N__31105));
    LocalMux I__7038 (
            .O(N__31158),
            .I(N__31105));
    LocalMux I__7037 (
            .O(N__31151),
            .I(N__31096));
    LocalMux I__7036 (
            .O(N__31148),
            .I(N__31096));
    LocalMux I__7035 (
            .O(N__31139),
            .I(N__31096));
    LocalMux I__7034 (
            .O(N__31130),
            .I(N__31096));
    InMux I__7033 (
            .O(N__31129),
            .I(N__31093));
    LocalMux I__7032 (
            .O(N__31120),
            .I(N__31090));
    InMux I__7031 (
            .O(N__31119),
            .I(N__31077));
    InMux I__7030 (
            .O(N__31118),
            .I(N__31077));
    InMux I__7029 (
            .O(N__31117),
            .I(N__31077));
    InMux I__7028 (
            .O(N__31116),
            .I(N__31077));
    InMux I__7027 (
            .O(N__31115),
            .I(N__31077));
    InMux I__7026 (
            .O(N__31114),
            .I(N__31077));
    InMux I__7025 (
            .O(N__31113),
            .I(N__31068));
    InMux I__7024 (
            .O(N__31112),
            .I(N__31068));
    InMux I__7023 (
            .O(N__31111),
            .I(N__31068));
    InMux I__7022 (
            .O(N__31110),
            .I(N__31068));
    Span4Mux_h I__7021 (
            .O(N__31105),
            .I(N__31061));
    Span4Mux_v I__7020 (
            .O(N__31096),
            .I(N__31061));
    LocalMux I__7019 (
            .O(N__31093),
            .I(N__31061));
    Span4Mux_h I__7018 (
            .O(N__31090),
            .I(N__31056));
    LocalMux I__7017 (
            .O(N__31077),
            .I(N__31056));
    LocalMux I__7016 (
            .O(N__31068),
            .I(\b2v_inst.data_a_escribir12_THRU_CO ));
    Odrv4 I__7015 (
            .O(N__31061),
            .I(\b2v_inst.data_a_escribir12_THRU_CO ));
    Odrv4 I__7014 (
            .O(N__31056),
            .I(\b2v_inst.data_a_escribir12_THRU_CO ));
    InMux I__7013 (
            .O(N__31049),
            .I(N__31046));
    LocalMux I__7012 (
            .O(N__31046),
            .I(\b2v_inst.un1_reg_anterior_0_i_1_2 ));
    InMux I__7011 (
            .O(N__31043),
            .I(N__31038));
    CascadeMux I__7010 (
            .O(N__31042),
            .I(N__31034));
    InMux I__7009 (
            .O(N__31041),
            .I(N__31031));
    LocalMux I__7008 (
            .O(N__31038),
            .I(N__31028));
    InMux I__7007 (
            .O(N__31037),
            .I(N__31025));
    InMux I__7006 (
            .O(N__31034),
            .I(N__31022));
    LocalMux I__7005 (
            .O(N__31031),
            .I(N__31019));
    Span4Mux_v I__7004 (
            .O(N__31028),
            .I(N__31014));
    LocalMux I__7003 (
            .O(N__31025),
            .I(N__31014));
    LocalMux I__7002 (
            .O(N__31022),
            .I(N__31011));
    Span4Mux_v I__7001 (
            .O(N__31019),
            .I(N__31007));
    Span4Mux_h I__7000 (
            .O(N__31014),
            .I(N__31002));
    Span4Mux_v I__6999 (
            .O(N__31011),
            .I(N__31002));
    InMux I__6998 (
            .O(N__31010),
            .I(N__30999));
    Odrv4 I__6997 (
            .O(N__31007),
            .I(\b2v_inst.reg_ancho_1Z0Z_3 ));
    Odrv4 I__6996 (
            .O(N__31002),
            .I(\b2v_inst.reg_ancho_1Z0Z_3 ));
    LocalMux I__6995 (
            .O(N__30999),
            .I(\b2v_inst.reg_ancho_1Z0Z_3 ));
    CascadeMux I__6994 (
            .O(N__30992),
            .I(N__30984));
    InMux I__6993 (
            .O(N__30991),
            .I(N__30972));
    InMux I__6992 (
            .O(N__30990),
            .I(N__30972));
    CascadeMux I__6991 (
            .O(N__30989),
            .I(N__30968));
    CascadeMux I__6990 (
            .O(N__30988),
            .I(N__30965));
    CascadeMux I__6989 (
            .O(N__30987),
            .I(N__30962));
    InMux I__6988 (
            .O(N__30984),
            .I(N__30958));
    CascadeMux I__6987 (
            .O(N__30983),
            .I(N__30953));
    CascadeMux I__6986 (
            .O(N__30982),
            .I(N__30950));
    CascadeMux I__6985 (
            .O(N__30981),
            .I(N__30947));
    CascadeMux I__6984 (
            .O(N__30980),
            .I(N__30942));
    CascadeMux I__6983 (
            .O(N__30979),
            .I(N__30938));
    CascadeMux I__6982 (
            .O(N__30978),
            .I(N__30935));
    InMux I__6981 (
            .O(N__30977),
            .I(N__30932));
    LocalMux I__6980 (
            .O(N__30972),
            .I(N__30928));
    InMux I__6979 (
            .O(N__30971),
            .I(N__30925));
    InMux I__6978 (
            .O(N__30968),
            .I(N__30922));
    InMux I__6977 (
            .O(N__30965),
            .I(N__30915));
    InMux I__6976 (
            .O(N__30962),
            .I(N__30915));
    InMux I__6975 (
            .O(N__30961),
            .I(N__30915));
    LocalMux I__6974 (
            .O(N__30958),
            .I(N__30912));
    InMux I__6973 (
            .O(N__30957),
            .I(N__30907));
    InMux I__6972 (
            .O(N__30956),
            .I(N__30904));
    InMux I__6971 (
            .O(N__30953),
            .I(N__30901));
    InMux I__6970 (
            .O(N__30950),
            .I(N__30894));
    InMux I__6969 (
            .O(N__30947),
            .I(N__30894));
    InMux I__6968 (
            .O(N__30946),
            .I(N__30894));
    InMux I__6967 (
            .O(N__30945),
            .I(N__30889));
    InMux I__6966 (
            .O(N__30942),
            .I(N__30889));
    InMux I__6965 (
            .O(N__30941),
            .I(N__30882));
    InMux I__6964 (
            .O(N__30938),
            .I(N__30882));
    InMux I__6963 (
            .O(N__30935),
            .I(N__30882));
    LocalMux I__6962 (
            .O(N__30932),
            .I(N__30879));
    CascadeMux I__6961 (
            .O(N__30931),
            .I(N__30876));
    Span4Mux_v I__6960 (
            .O(N__30928),
            .I(N__30869));
    LocalMux I__6959 (
            .O(N__30925),
            .I(N__30869));
    LocalMux I__6958 (
            .O(N__30922),
            .I(N__30862));
    LocalMux I__6957 (
            .O(N__30915),
            .I(N__30862));
    Span4Mux_v I__6956 (
            .O(N__30912),
            .I(N__30862));
    CascadeMux I__6955 (
            .O(N__30911),
            .I(N__30857));
    CascadeMux I__6954 (
            .O(N__30910),
            .I(N__30854));
    LocalMux I__6953 (
            .O(N__30907),
            .I(N__30849));
    LocalMux I__6952 (
            .O(N__30904),
            .I(N__30849));
    LocalMux I__6951 (
            .O(N__30901),
            .I(N__30846));
    LocalMux I__6950 (
            .O(N__30894),
            .I(N__30843));
    LocalMux I__6949 (
            .O(N__30889),
            .I(N__30840));
    LocalMux I__6948 (
            .O(N__30882),
            .I(N__30837));
    Span4Mux_v I__6947 (
            .O(N__30879),
            .I(N__30834));
    InMux I__6946 (
            .O(N__30876),
            .I(N__30831));
    InMux I__6945 (
            .O(N__30875),
            .I(N__30828));
    InMux I__6944 (
            .O(N__30874),
            .I(N__30825));
    Span4Mux_h I__6943 (
            .O(N__30869),
            .I(N__30820));
    Span4Mux_h I__6942 (
            .O(N__30862),
            .I(N__30820));
    InMux I__6941 (
            .O(N__30861),
            .I(N__30811));
    InMux I__6940 (
            .O(N__30860),
            .I(N__30811));
    InMux I__6939 (
            .O(N__30857),
            .I(N__30811));
    InMux I__6938 (
            .O(N__30854),
            .I(N__30811));
    Span4Mux_v I__6937 (
            .O(N__30849),
            .I(N__30806));
    Span4Mux_v I__6936 (
            .O(N__30846),
            .I(N__30806));
    Span4Mux_v I__6935 (
            .O(N__30843),
            .I(N__30799));
    Span4Mux_v I__6934 (
            .O(N__30840),
            .I(N__30799));
    Span4Mux_v I__6933 (
            .O(N__30837),
            .I(N__30799));
    Span4Mux_h I__6932 (
            .O(N__30834),
            .I(N__30792));
    LocalMux I__6931 (
            .O(N__30831),
            .I(N__30792));
    LocalMux I__6930 (
            .O(N__30828),
            .I(N__30792));
    LocalMux I__6929 (
            .O(N__30825),
            .I(N__30787));
    Span4Mux_h I__6928 (
            .O(N__30820),
            .I(N__30787));
    LocalMux I__6927 (
            .O(N__30811),
            .I(N__30780));
    Sp12to4 I__6926 (
            .O(N__30806),
            .I(N__30780));
    Sp12to4 I__6925 (
            .O(N__30799),
            .I(N__30780));
    Span4Mux_h I__6924 (
            .O(N__30792),
            .I(N__30777));
    Odrv4 I__6923 (
            .O(N__30787),
            .I(\b2v_inst.stateZ0Z_20 ));
    Odrv12 I__6922 (
            .O(N__30780),
            .I(\b2v_inst.stateZ0Z_20 ));
    Odrv4 I__6921 (
            .O(N__30777),
            .I(\b2v_inst.stateZ0Z_20 ));
    InMux I__6920 (
            .O(N__30770),
            .I(N__30765));
    InMux I__6919 (
            .O(N__30769),
            .I(N__30762));
    InMux I__6918 (
            .O(N__30768),
            .I(N__30758));
    LocalMux I__6917 (
            .O(N__30765),
            .I(N__30755));
    LocalMux I__6916 (
            .O(N__30762),
            .I(N__30752));
    InMux I__6915 (
            .O(N__30761),
            .I(N__30749));
    LocalMux I__6914 (
            .O(N__30758),
            .I(N__30746));
    Span4Mux_v I__6913 (
            .O(N__30755),
            .I(N__30743));
    Span4Mux_h I__6912 (
            .O(N__30752),
            .I(N__30738));
    LocalMux I__6911 (
            .O(N__30749),
            .I(N__30738));
    Span4Mux_v I__6910 (
            .O(N__30746),
            .I(N__30733));
    Span4Mux_h I__6909 (
            .O(N__30743),
            .I(N__30733));
    Odrv4 I__6908 (
            .O(N__30738),
            .I(\b2v_inst.reg_anteriorZ0Z_8 ));
    Odrv4 I__6907 (
            .O(N__30733),
            .I(\b2v_inst.reg_anteriorZ0Z_8 ));
    InMux I__6906 (
            .O(N__30728),
            .I(N__30725));
    LocalMux I__6905 (
            .O(N__30725),
            .I(N__30720));
    InMux I__6904 (
            .O(N__30724),
            .I(N__30717));
    InMux I__6903 (
            .O(N__30723),
            .I(N__30714));
    Span4Mux_v I__6902 (
            .O(N__30720),
            .I(N__30709));
    LocalMux I__6901 (
            .O(N__30717),
            .I(N__30709));
    LocalMux I__6900 (
            .O(N__30714),
            .I(\b2v_inst.reg_ancho_3Z0Z_8 ));
    Odrv4 I__6899 (
            .O(N__30709),
            .I(\b2v_inst.reg_ancho_3Z0Z_8 ));
    InMux I__6898 (
            .O(N__30704),
            .I(N__30701));
    LocalMux I__6897 (
            .O(N__30701),
            .I(\b2v_inst.N_544 ));
    InMux I__6896 (
            .O(N__30698),
            .I(N__30695));
    LocalMux I__6895 (
            .O(N__30695),
            .I(N__30692));
    Span4Mux_v I__6894 (
            .O(N__30692),
            .I(N__30687));
    InMux I__6893 (
            .O(N__30691),
            .I(N__30684));
    InMux I__6892 (
            .O(N__30690),
            .I(N__30681));
    Odrv4 I__6891 (
            .O(N__30687),
            .I(\b2v_inst.reg_ancho_3Z0Z_7 ));
    LocalMux I__6890 (
            .O(N__30684),
            .I(\b2v_inst.reg_ancho_3Z0Z_7 ));
    LocalMux I__6889 (
            .O(N__30681),
            .I(\b2v_inst.reg_ancho_3Z0Z_7 ));
    CascadeMux I__6888 (
            .O(N__30674),
            .I(N__30671));
    InMux I__6887 (
            .O(N__30671),
            .I(N__30664));
    InMux I__6886 (
            .O(N__30670),
            .I(N__30664));
    InMux I__6885 (
            .O(N__30669),
            .I(N__30661));
    LocalMux I__6884 (
            .O(N__30664),
            .I(N__30658));
    LocalMux I__6883 (
            .O(N__30661),
            .I(N__30654));
    Span4Mux_h I__6882 (
            .O(N__30658),
            .I(N__30651));
    InMux I__6881 (
            .O(N__30657),
            .I(N__30648));
    Span4Mux_h I__6880 (
            .O(N__30654),
            .I(N__30645));
    Odrv4 I__6879 (
            .O(N__30651),
            .I(\b2v_inst.reg_anteriorZ0Z_7 ));
    LocalMux I__6878 (
            .O(N__30648),
            .I(\b2v_inst.reg_anteriorZ0Z_7 ));
    Odrv4 I__6877 (
            .O(N__30645),
            .I(\b2v_inst.reg_anteriorZ0Z_7 ));
    InMux I__6876 (
            .O(N__30638),
            .I(N__30635));
    LocalMux I__6875 (
            .O(N__30635),
            .I(\b2v_inst.un1_reg_anterior_0_i_1_7 ));
    CascadeMux I__6874 (
            .O(N__30632),
            .I(\b2v_inst.data_a_escribir_RNO_0Z0Z_7_cascade_ ));
    InMux I__6873 (
            .O(N__30629),
            .I(N__30615));
    InMux I__6872 (
            .O(N__30628),
            .I(N__30615));
    InMux I__6871 (
            .O(N__30627),
            .I(N__30615));
    InMux I__6870 (
            .O(N__30626),
            .I(N__30601));
    InMux I__6869 (
            .O(N__30625),
            .I(N__30601));
    InMux I__6868 (
            .O(N__30624),
            .I(N__30594));
    InMux I__6867 (
            .O(N__30623),
            .I(N__30594));
    InMux I__6866 (
            .O(N__30622),
            .I(N__30594));
    LocalMux I__6865 (
            .O(N__30615),
            .I(N__30591));
    InMux I__6864 (
            .O(N__30614),
            .I(N__30584));
    InMux I__6863 (
            .O(N__30613),
            .I(N__30584));
    InMux I__6862 (
            .O(N__30612),
            .I(N__30584));
    InMux I__6861 (
            .O(N__30611),
            .I(N__30577));
    InMux I__6860 (
            .O(N__30610),
            .I(N__30577));
    InMux I__6859 (
            .O(N__30609),
            .I(N__30577));
    InMux I__6858 (
            .O(N__30608),
            .I(N__30570));
    InMux I__6857 (
            .O(N__30607),
            .I(N__30570));
    InMux I__6856 (
            .O(N__30606),
            .I(N__30570));
    LocalMux I__6855 (
            .O(N__30601),
            .I(\b2v_inst.N_711 ));
    LocalMux I__6854 (
            .O(N__30594),
            .I(\b2v_inst.N_711 ));
    Odrv4 I__6853 (
            .O(N__30591),
            .I(\b2v_inst.N_711 ));
    LocalMux I__6852 (
            .O(N__30584),
            .I(\b2v_inst.N_711 ));
    LocalMux I__6851 (
            .O(N__30577),
            .I(\b2v_inst.N_711 ));
    LocalMux I__6850 (
            .O(N__30570),
            .I(\b2v_inst.N_711 ));
    CEMux I__6849 (
            .O(N__30557),
            .I(N__30549));
    CEMux I__6848 (
            .O(N__30556),
            .I(N__30546));
    CEMux I__6847 (
            .O(N__30555),
            .I(N__30543));
    CEMux I__6846 (
            .O(N__30554),
            .I(N__30540));
    CEMux I__6845 (
            .O(N__30553),
            .I(N__30537));
    CEMux I__6844 (
            .O(N__30552),
            .I(N__30534));
    LocalMux I__6843 (
            .O(N__30549),
            .I(N__30531));
    LocalMux I__6842 (
            .O(N__30546),
            .I(N__30528));
    LocalMux I__6841 (
            .O(N__30543),
            .I(N__30525));
    LocalMux I__6840 (
            .O(N__30540),
            .I(N__30522));
    LocalMux I__6839 (
            .O(N__30537),
            .I(N__30517));
    LocalMux I__6838 (
            .O(N__30534),
            .I(N__30517));
    Span4Mux_h I__6837 (
            .O(N__30531),
            .I(N__30512));
    Span4Mux_h I__6836 (
            .O(N__30528),
            .I(N__30512));
    Odrv4 I__6835 (
            .O(N__30525),
            .I(\b2v_inst.un1_reset_inv_0 ));
    Odrv4 I__6834 (
            .O(N__30522),
            .I(\b2v_inst.un1_reset_inv_0 ));
    Odrv4 I__6833 (
            .O(N__30517),
            .I(\b2v_inst.un1_reset_inv_0 ));
    Odrv4 I__6832 (
            .O(N__30512),
            .I(\b2v_inst.un1_reset_inv_0 ));
    InMux I__6831 (
            .O(N__30503),
            .I(N__30500));
    LocalMux I__6830 (
            .O(N__30500),
            .I(\b2v_inst9.un1_cycle_counter_2_cry_1_THRU_CO ));
    CascadeMux I__6829 (
            .O(N__30497),
            .I(N__30494));
    InMux I__6828 (
            .O(N__30494),
            .I(N__30488));
    InMux I__6827 (
            .O(N__30493),
            .I(N__30485));
    InMux I__6826 (
            .O(N__30492),
            .I(N__30480));
    InMux I__6825 (
            .O(N__30491),
            .I(N__30480));
    LocalMux I__6824 (
            .O(N__30488),
            .I(\b2v_inst9.cycle_counterZ0Z_2 ));
    LocalMux I__6823 (
            .O(N__30485),
            .I(\b2v_inst9.cycle_counterZ0Z_2 ));
    LocalMux I__6822 (
            .O(N__30480),
            .I(\b2v_inst9.cycle_counterZ0Z_2 ));
    InMux I__6821 (
            .O(N__30473),
            .I(N__30468));
    InMux I__6820 (
            .O(N__30472),
            .I(N__30463));
    InMux I__6819 (
            .O(N__30471),
            .I(N__30460));
    LocalMux I__6818 (
            .O(N__30468),
            .I(N__30457));
    InMux I__6817 (
            .O(N__30467),
            .I(N__30452));
    InMux I__6816 (
            .O(N__30466),
            .I(N__30452));
    LocalMux I__6815 (
            .O(N__30463),
            .I(N__30449));
    LocalMux I__6814 (
            .O(N__30460),
            .I(N__30446));
    Span4Mux_h I__6813 (
            .O(N__30457),
            .I(N__30443));
    LocalMux I__6812 (
            .O(N__30452),
            .I(\b2v_inst9.cycle_counter_RNIQAGDZ0Z_3 ));
    Odrv4 I__6811 (
            .O(N__30449),
            .I(\b2v_inst9.cycle_counter_RNIQAGDZ0Z_3 ));
    Odrv4 I__6810 (
            .O(N__30446),
            .I(\b2v_inst9.cycle_counter_RNIQAGDZ0Z_3 ));
    Odrv4 I__6809 (
            .O(N__30443),
            .I(\b2v_inst9.cycle_counter_RNIQAGDZ0Z_3 ));
    CascadeMux I__6808 (
            .O(N__30434),
            .I(N__30430));
    InMux I__6807 (
            .O(N__30433),
            .I(N__30427));
    InMux I__6806 (
            .O(N__30430),
            .I(N__30423));
    LocalMux I__6805 (
            .O(N__30427),
            .I(N__30413));
    InMux I__6804 (
            .O(N__30426),
            .I(N__30408));
    LocalMux I__6803 (
            .O(N__30423),
            .I(N__30405));
    InMux I__6802 (
            .O(N__30422),
            .I(N__30402));
    InMux I__6801 (
            .O(N__30421),
            .I(N__30397));
    InMux I__6800 (
            .O(N__30420),
            .I(N__30397));
    InMux I__6799 (
            .O(N__30419),
            .I(N__30390));
    InMux I__6798 (
            .O(N__30418),
            .I(N__30390));
    InMux I__6797 (
            .O(N__30417),
            .I(N__30390));
    InMux I__6796 (
            .O(N__30416),
            .I(N__30387));
    Span4Mux_v I__6795 (
            .O(N__30413),
            .I(N__30384));
    CascadeMux I__6794 (
            .O(N__30412),
            .I(N__30380));
    CascadeMux I__6793 (
            .O(N__30411),
            .I(N__30372));
    LocalMux I__6792 (
            .O(N__30408),
            .I(N__30368));
    Span4Mux_v I__6791 (
            .O(N__30405),
            .I(N__30361));
    LocalMux I__6790 (
            .O(N__30402),
            .I(N__30361));
    LocalMux I__6789 (
            .O(N__30397),
            .I(N__30361));
    LocalMux I__6788 (
            .O(N__30390),
            .I(N__30358));
    LocalMux I__6787 (
            .O(N__30387),
            .I(N__30355));
    Span4Mux_h I__6786 (
            .O(N__30384),
            .I(N__30352));
    InMux I__6785 (
            .O(N__30383),
            .I(N__30343));
    InMux I__6784 (
            .O(N__30380),
            .I(N__30343));
    InMux I__6783 (
            .O(N__30379),
            .I(N__30343));
    InMux I__6782 (
            .O(N__30378),
            .I(N__30343));
    InMux I__6781 (
            .O(N__30377),
            .I(N__30338));
    InMux I__6780 (
            .O(N__30376),
            .I(N__30338));
    InMux I__6779 (
            .O(N__30375),
            .I(N__30335));
    InMux I__6778 (
            .O(N__30372),
            .I(N__30330));
    InMux I__6777 (
            .O(N__30371),
            .I(N__30330));
    Span4Mux_v I__6776 (
            .O(N__30368),
            .I(N__30321));
    Span4Mux_h I__6775 (
            .O(N__30361),
            .I(N__30321));
    Span4Mux_v I__6774 (
            .O(N__30358),
            .I(N__30321));
    Span4Mux_v I__6773 (
            .O(N__30355),
            .I(N__30321));
    Odrv4 I__6772 (
            .O(N__30352),
            .I(N_478));
    LocalMux I__6771 (
            .O(N__30343),
            .I(N_478));
    LocalMux I__6770 (
            .O(N__30338),
            .I(N_478));
    LocalMux I__6769 (
            .O(N__30335),
            .I(N_478));
    LocalMux I__6768 (
            .O(N__30330),
            .I(N_478));
    Odrv4 I__6767 (
            .O(N__30321),
            .I(N_478));
    CascadeMux I__6766 (
            .O(N__30308),
            .I(N__30305));
    InMux I__6765 (
            .O(N__30305),
            .I(N__30299));
    InMux I__6764 (
            .O(N__30304),
            .I(N__30294));
    InMux I__6763 (
            .O(N__30303),
            .I(N__30294));
    InMux I__6762 (
            .O(N__30302),
            .I(N__30291));
    LocalMux I__6761 (
            .O(N__30299),
            .I(N__30286));
    LocalMux I__6760 (
            .O(N__30294),
            .I(N__30286));
    LocalMux I__6759 (
            .O(N__30291),
            .I(\b2v_inst9.cycle_counterZ0Z_0 ));
    Odrv4 I__6758 (
            .O(N__30286),
            .I(\b2v_inst9.cycle_counterZ0Z_0 ));
    InMux I__6757 (
            .O(N__30281),
            .I(N__30278));
    LocalMux I__6756 (
            .O(N__30278),
            .I(N__30274));
    CascadeMux I__6755 (
            .O(N__30277),
            .I(N__30271));
    Span4Mux_h I__6754 (
            .O(N__30274),
            .I(N__30268));
    InMux I__6753 (
            .O(N__30271),
            .I(N__30265));
    Odrv4 I__6752 (
            .O(N__30268),
            .I(SYNTHESIZED_WIRE_5_3));
    LocalMux I__6751 (
            .O(N__30265),
            .I(SYNTHESIZED_WIRE_5_3));
    InMux I__6750 (
            .O(N__30260),
            .I(N__30257));
    LocalMux I__6749 (
            .O(N__30257),
            .I(N__30254));
    Span4Mux_h I__6748 (
            .O(N__30254),
            .I(N__30251));
    Odrv4 I__6747 (
            .O(N__30251),
            .I(\b2v_inst.pix_data_regZ0Z_3 ));
    CEMux I__6746 (
            .O(N__30248),
            .I(N__30245));
    LocalMux I__6745 (
            .O(N__30245),
            .I(N__30240));
    CEMux I__6744 (
            .O(N__30244),
            .I(N__30237));
    CEMux I__6743 (
            .O(N__30243),
            .I(N__30234));
    Sp12to4 I__6742 (
            .O(N__30240),
            .I(N__30227));
    LocalMux I__6741 (
            .O(N__30237),
            .I(N__30227));
    LocalMux I__6740 (
            .O(N__30234),
            .I(N__30224));
    InMux I__6739 (
            .O(N__30233),
            .I(N__30221));
    InMux I__6738 (
            .O(N__30232),
            .I(N__30218));
    Span12Mux_h I__6737 (
            .O(N__30227),
            .I(N__30214));
    Span4Mux_v I__6736 (
            .O(N__30224),
            .I(N__30211));
    LocalMux I__6735 (
            .O(N__30221),
            .I(N__30208));
    LocalMux I__6734 (
            .O(N__30218),
            .I(N__30205));
    InMux I__6733 (
            .O(N__30217),
            .I(N__30202));
    Odrv12 I__6732 (
            .O(N__30214),
            .I(\b2v_inst.stateZ0Z_24 ));
    Odrv4 I__6731 (
            .O(N__30211),
            .I(\b2v_inst.stateZ0Z_24 ));
    Odrv4 I__6730 (
            .O(N__30208),
            .I(\b2v_inst.stateZ0Z_24 ));
    Odrv4 I__6729 (
            .O(N__30205),
            .I(\b2v_inst.stateZ0Z_24 ));
    LocalMux I__6728 (
            .O(N__30202),
            .I(\b2v_inst.stateZ0Z_24 ));
    CascadeMux I__6727 (
            .O(N__30191),
            .I(N__30188));
    InMux I__6726 (
            .O(N__30188),
            .I(N__30185));
    LocalMux I__6725 (
            .O(N__30185),
            .I(N__30182));
    Span4Mux_h I__6724 (
            .O(N__30182),
            .I(N__30179));
    Odrv4 I__6723 (
            .O(N__30179),
            .I(SYNTHESIZED_WIRE_1_2));
    InMux I__6722 (
            .O(N__30176),
            .I(N__30172));
    InMux I__6721 (
            .O(N__30175),
            .I(N__30168));
    LocalMux I__6720 (
            .O(N__30172),
            .I(N__30165));
    InMux I__6719 (
            .O(N__30171),
            .I(N__30162));
    LocalMux I__6718 (
            .O(N__30168),
            .I(N__30159));
    Span4Mux_v I__6717 (
            .O(N__30165),
            .I(N__30153));
    LocalMux I__6716 (
            .O(N__30162),
            .I(N__30153));
    Span12Mux_v I__6715 (
            .O(N__30159),
            .I(N__30150));
    InMux I__6714 (
            .O(N__30158),
            .I(N__30147));
    Span4Mux_v I__6713 (
            .O(N__30153),
            .I(N__30144));
    Odrv12 I__6712 (
            .O(N__30150),
            .I(\b2v_inst.reg_anteriorZ0Z_4 ));
    LocalMux I__6711 (
            .O(N__30147),
            .I(\b2v_inst.reg_anteriorZ0Z_4 ));
    Odrv4 I__6710 (
            .O(N__30144),
            .I(\b2v_inst.reg_anteriorZ0Z_4 ));
    InMux I__6709 (
            .O(N__30137),
            .I(N__30133));
    CascadeMux I__6708 (
            .O(N__30136),
            .I(N__30129));
    LocalMux I__6707 (
            .O(N__30133),
            .I(N__30126));
    InMux I__6706 (
            .O(N__30132),
            .I(N__30123));
    InMux I__6705 (
            .O(N__30129),
            .I(N__30120));
    Span4Mux_v I__6704 (
            .O(N__30126),
            .I(N__30115));
    LocalMux I__6703 (
            .O(N__30123),
            .I(N__30115));
    LocalMux I__6702 (
            .O(N__30120),
            .I(\b2v_inst.reg_ancho_3Z0Z_9 ));
    Odrv4 I__6701 (
            .O(N__30115),
            .I(\b2v_inst.reg_ancho_3Z0Z_9 ));
    InMux I__6700 (
            .O(N__30110),
            .I(N__30106));
    InMux I__6699 (
            .O(N__30109),
            .I(N__30103));
    LocalMux I__6698 (
            .O(N__30106),
            .I(N__30100));
    LocalMux I__6697 (
            .O(N__30103),
            .I(\b2v_inst.eventosZ0Z_9 ));
    Odrv4 I__6696 (
            .O(N__30100),
            .I(\b2v_inst.eventosZ0Z_9 ));
    InMux I__6695 (
            .O(N__30095),
            .I(N__30092));
    LocalMux I__6694 (
            .O(N__30092),
            .I(\b2v_inst.N_545 ));
    CascadeMux I__6693 (
            .O(N__30089),
            .I(\b2v_inst.un1_reg_anterior_iv_0_0_0_9_cascade_ ));
    InMux I__6692 (
            .O(N__30086),
            .I(N__30083));
    LocalMux I__6691 (
            .O(N__30083),
            .I(N__30080));
    Odrv4 I__6690 (
            .O(N__30080),
            .I(\b2v_inst.N_543 ));
    CascadeMux I__6689 (
            .O(N__30077),
            .I(\b2v_inst.un1_reg_anterior_iv_0_0_1_9_cascade_ ));
    CascadeMux I__6688 (
            .O(N__30074),
            .I(N__30071));
    InMux I__6687 (
            .O(N__30071),
            .I(N__30068));
    LocalMux I__6686 (
            .O(N__30068),
            .I(N__30065));
    Span4Mux_v I__6685 (
            .O(N__30065),
            .I(N__30062));
    Odrv4 I__6684 (
            .O(N__30062),
            .I(\b2v_inst.valor_max2_6 ));
    InMux I__6683 (
            .O(N__30059),
            .I(N__30056));
    LocalMux I__6682 (
            .O(N__30056),
            .I(N__30053));
    Odrv4 I__6681 (
            .O(N__30053),
            .I(\b2v_inst.un1_reg_anterior_iv_0_1_6 ));
    InMux I__6680 (
            .O(N__30050),
            .I(N__30047));
    LocalMux I__6679 (
            .O(N__30047),
            .I(N__30044));
    Span4Mux_h I__6678 (
            .O(N__30044),
            .I(N__30041));
    Odrv4 I__6677 (
            .O(N__30041),
            .I(\b2v_inst.data_a_escribir11_10_and ));
    InMux I__6676 (
            .O(N__30038),
            .I(N__30035));
    LocalMux I__6675 (
            .O(N__30035),
            .I(N__30031));
    InMux I__6674 (
            .O(N__30034),
            .I(N__30028));
    Span4Mux_h I__6673 (
            .O(N__30031),
            .I(N__30025));
    LocalMux I__6672 (
            .O(N__30028),
            .I(\b2v_inst.eventosZ0Z_8 ));
    Odrv4 I__6671 (
            .O(N__30025),
            .I(\b2v_inst.eventosZ0Z_8 ));
    CascadeMux I__6670 (
            .O(N__30020),
            .I(\b2v_inst.un1_reg_anterior_iv_0_0_0_8_cascade_ ));
    InMux I__6669 (
            .O(N__30017),
            .I(N__30014));
    LocalMux I__6668 (
            .O(N__30014),
            .I(N__30011));
    Odrv12 I__6667 (
            .O(N__30011),
            .I(\b2v_inst.N_542 ));
    CascadeMux I__6666 (
            .O(N__30008),
            .I(\b2v_inst.un1_reg_anterior_iv_0_0_1_8_cascade_ ));
    InMux I__6665 (
            .O(N__30005),
            .I(N__30000));
    InMux I__6664 (
            .O(N__30004),
            .I(N__29997));
    InMux I__6663 (
            .O(N__30003),
            .I(N__29994));
    LocalMux I__6662 (
            .O(N__30000),
            .I(N__29989));
    LocalMux I__6661 (
            .O(N__29997),
            .I(N__29989));
    LocalMux I__6660 (
            .O(N__29994),
            .I(N__29984));
    Span4Mux_h I__6659 (
            .O(N__29989),
            .I(N__29981));
    InMux I__6658 (
            .O(N__29988),
            .I(N__29978));
    InMux I__6657 (
            .O(N__29987),
            .I(N__29975));
    Odrv4 I__6656 (
            .O(N__29984),
            .I(\b2v_inst.reg_ancho_1Z0Z_9 ));
    Odrv4 I__6655 (
            .O(N__29981),
            .I(\b2v_inst.reg_ancho_1Z0Z_9 ));
    LocalMux I__6654 (
            .O(N__29978),
            .I(\b2v_inst.reg_ancho_1Z0Z_9 ));
    LocalMux I__6653 (
            .O(N__29975),
            .I(\b2v_inst.reg_ancho_1Z0Z_9 ));
    InMux I__6652 (
            .O(N__29966),
            .I(N__29961));
    InMux I__6651 (
            .O(N__29965),
            .I(N__29956));
    InMux I__6650 (
            .O(N__29964),
            .I(N__29956));
    LocalMux I__6649 (
            .O(N__29961),
            .I(N__29953));
    LocalMux I__6648 (
            .O(N__29956),
            .I(N__29950));
    Span4Mux_v I__6647 (
            .O(N__29953),
            .I(N__29945));
    Span4Mux_h I__6646 (
            .O(N__29950),
            .I(N__29942));
    InMux I__6645 (
            .O(N__29949),
            .I(N__29939));
    InMux I__6644 (
            .O(N__29948),
            .I(N__29936));
    Odrv4 I__6643 (
            .O(N__29945),
            .I(\b2v_inst.reg_ancho_1Z0Z_8 ));
    Odrv4 I__6642 (
            .O(N__29942),
            .I(\b2v_inst.reg_ancho_1Z0Z_8 ));
    LocalMux I__6641 (
            .O(N__29939),
            .I(\b2v_inst.reg_ancho_1Z0Z_8 ));
    LocalMux I__6640 (
            .O(N__29936),
            .I(\b2v_inst.reg_ancho_1Z0Z_8 ));
    InMux I__6639 (
            .O(N__29927),
            .I(N__29922));
    CascadeMux I__6638 (
            .O(N__29926),
            .I(N__29919));
    InMux I__6637 (
            .O(N__29925),
            .I(N__29916));
    LocalMux I__6636 (
            .O(N__29922),
            .I(N__29913));
    InMux I__6635 (
            .O(N__29919),
            .I(N__29910));
    LocalMux I__6634 (
            .O(N__29916),
            .I(N__29906));
    Span4Mux_v I__6633 (
            .O(N__29913),
            .I(N__29903));
    LocalMux I__6632 (
            .O(N__29910),
            .I(N__29900));
    CascadeMux I__6631 (
            .O(N__29909),
            .I(N__29896));
    Span4Mux_v I__6630 (
            .O(N__29906),
            .I(N__29891));
    Span4Mux_h I__6629 (
            .O(N__29903),
            .I(N__29891));
    Span4Mux_h I__6628 (
            .O(N__29900),
            .I(N__29888));
    InMux I__6627 (
            .O(N__29899),
            .I(N__29885));
    InMux I__6626 (
            .O(N__29896),
            .I(N__29882));
    Odrv4 I__6625 (
            .O(N__29891),
            .I(\b2v_inst.reg_ancho_2Z0Z_8 ));
    Odrv4 I__6624 (
            .O(N__29888),
            .I(\b2v_inst.reg_ancho_2Z0Z_8 ));
    LocalMux I__6623 (
            .O(N__29885),
            .I(\b2v_inst.reg_ancho_2Z0Z_8 ));
    LocalMux I__6622 (
            .O(N__29882),
            .I(\b2v_inst.reg_ancho_2Z0Z_8 ));
    CascadeMux I__6621 (
            .O(N__29873),
            .I(N__29870));
    InMux I__6620 (
            .O(N__29870),
            .I(N__29867));
    LocalMux I__6619 (
            .O(N__29867),
            .I(N__29864));
    Span4Mux_h I__6618 (
            .O(N__29864),
            .I(N__29860));
    InMux I__6617 (
            .O(N__29863),
            .I(N__29857));
    Odrv4 I__6616 (
            .O(N__29860),
            .I(\b2v_inst.eventosZ0Z_3 ));
    LocalMux I__6615 (
            .O(N__29857),
            .I(\b2v_inst.eventosZ0Z_3 ));
    InMux I__6614 (
            .O(N__29852),
            .I(N__29849));
    LocalMux I__6613 (
            .O(N__29849),
            .I(N__29846));
    Span4Mux_h I__6612 (
            .O(N__29846),
            .I(N__29843));
    Odrv4 I__6611 (
            .O(N__29843),
            .I(\b2v_inst.un1_reg_anterior_0_i_1_3 ));
    CascadeMux I__6610 (
            .O(N__29840),
            .I(N__29834));
    InMux I__6609 (
            .O(N__29839),
            .I(N__29831));
    InMux I__6608 (
            .O(N__29838),
            .I(N__29828));
    InMux I__6607 (
            .O(N__29837),
            .I(N__29825));
    InMux I__6606 (
            .O(N__29834),
            .I(N__29822));
    LocalMux I__6605 (
            .O(N__29831),
            .I(N__29819));
    LocalMux I__6604 (
            .O(N__29828),
            .I(N__29814));
    LocalMux I__6603 (
            .O(N__29825),
            .I(N__29814));
    LocalMux I__6602 (
            .O(N__29822),
            .I(N__29811));
    Span4Mux_h I__6601 (
            .O(N__29819),
            .I(N__29806));
    Span4Mux_v I__6600 (
            .O(N__29814),
            .I(N__29806));
    Odrv4 I__6599 (
            .O(N__29811),
            .I(\b2v_inst.reg_anteriorZ0Z_2 ));
    Odrv4 I__6598 (
            .O(N__29806),
            .I(\b2v_inst.reg_anteriorZ0Z_2 ));
    InMux I__6597 (
            .O(N__29801),
            .I(N__29798));
    LocalMux I__6596 (
            .O(N__29798),
            .I(N__29795));
    Span4Mux_h I__6595 (
            .O(N__29795),
            .I(N__29792));
    Odrv4 I__6594 (
            .O(N__29792),
            .I(\b2v_inst.data_a_escribir11_6_and ));
    InMux I__6593 (
            .O(N__29789),
            .I(N__29786));
    LocalMux I__6592 (
            .O(N__29786),
            .I(N__29783));
    Span4Mux_v I__6591 (
            .O(N__29783),
            .I(N__29780));
    Sp12to4 I__6590 (
            .O(N__29780),
            .I(N__29777));
    Odrv12 I__6589 (
            .O(N__29777),
            .I(\b2v_inst.N_273 ));
    CascadeMux I__6588 (
            .O(N__29774),
            .I(N__29771));
    InMux I__6587 (
            .O(N__29771),
            .I(N__29768));
    LocalMux I__6586 (
            .O(N__29768),
            .I(\b2v_inst.un1_reg_anterior_iv_0_0_5 ));
    InMux I__6585 (
            .O(N__29765),
            .I(N__29762));
    LocalMux I__6584 (
            .O(N__29762),
            .I(N__29759));
    Span4Mux_v I__6583 (
            .O(N__29759),
            .I(N__29756));
    Odrv4 I__6582 (
            .O(N__29756),
            .I(\b2v_inst.N_267 ));
    CascadeMux I__6581 (
            .O(N__29753),
            .I(\b2v_inst.un1_reg_anterior_iv_0_1_5_cascade_ ));
    CascadeMux I__6580 (
            .O(N__29750),
            .I(N__29747));
    InMux I__6579 (
            .O(N__29747),
            .I(N__29744));
    LocalMux I__6578 (
            .O(N__29744),
            .I(\b2v_inst.data_a_escribir_RNO_0Z0Z_2 ));
    CascadeMux I__6577 (
            .O(N__29741),
            .I(N__29738));
    InMux I__6576 (
            .O(N__29738),
            .I(N__29733));
    InMux I__6575 (
            .O(N__29737),
            .I(N__29730));
    InMux I__6574 (
            .O(N__29736),
            .I(N__29727));
    LocalMux I__6573 (
            .O(N__29733),
            .I(N__29718));
    LocalMux I__6572 (
            .O(N__29730),
            .I(N__29718));
    LocalMux I__6571 (
            .O(N__29727),
            .I(N__29718));
    InMux I__6570 (
            .O(N__29726),
            .I(N__29715));
    InMux I__6569 (
            .O(N__29725),
            .I(N__29712));
    Span4Mux_v I__6568 (
            .O(N__29718),
            .I(N__29709));
    LocalMux I__6567 (
            .O(N__29715),
            .I(\b2v_inst.reg_ancho_2Z0Z_9 ));
    LocalMux I__6566 (
            .O(N__29712),
            .I(\b2v_inst.reg_ancho_2Z0Z_9 ));
    Odrv4 I__6565 (
            .O(N__29709),
            .I(\b2v_inst.reg_ancho_2Z0Z_9 ));
    InMux I__6564 (
            .O(N__29702),
            .I(N__29698));
    InMux I__6563 (
            .O(N__29701),
            .I(N__29695));
    LocalMux I__6562 (
            .O(N__29698),
            .I(N__29692));
    LocalMux I__6561 (
            .O(N__29695),
            .I(N__29688));
    Span4Mux_v I__6560 (
            .O(N__29692),
            .I(N__29685));
    InMux I__6559 (
            .O(N__29691),
            .I(N__29682));
    Odrv4 I__6558 (
            .O(N__29688),
            .I(\b2v_inst.reg_ancho_3Z0Z_1 ));
    Odrv4 I__6557 (
            .O(N__29685),
            .I(\b2v_inst.reg_ancho_3Z0Z_1 ));
    LocalMux I__6556 (
            .O(N__29682),
            .I(\b2v_inst.reg_ancho_3Z0Z_1 ));
    InMux I__6555 (
            .O(N__29675),
            .I(N__29671));
    InMux I__6554 (
            .O(N__29674),
            .I(N__29668));
    LocalMux I__6553 (
            .O(N__29671),
            .I(N__29665));
    LocalMux I__6552 (
            .O(N__29668),
            .I(N__29661));
    Span4Mux_v I__6551 (
            .O(N__29665),
            .I(N__29658));
    InMux I__6550 (
            .O(N__29664),
            .I(N__29655));
    Odrv4 I__6549 (
            .O(N__29661),
            .I(\b2v_inst.reg_ancho_3Z0Z_0 ));
    Odrv4 I__6548 (
            .O(N__29658),
            .I(\b2v_inst.reg_ancho_3Z0Z_0 ));
    LocalMux I__6547 (
            .O(N__29655),
            .I(\b2v_inst.reg_ancho_3Z0Z_0 ));
    InMux I__6546 (
            .O(N__29648),
            .I(N__29645));
    LocalMux I__6545 (
            .O(N__29645),
            .I(N__29642));
    Span4Mux_h I__6544 (
            .O(N__29642),
            .I(N__29639));
    Odrv4 I__6543 (
            .O(N__29639),
            .I(\b2v_inst.data_a_escribir11_5_and ));
    InMux I__6542 (
            .O(N__29636),
            .I(N__29630));
    InMux I__6541 (
            .O(N__29635),
            .I(N__29627));
    InMux I__6540 (
            .O(N__29634),
            .I(N__29622));
    InMux I__6539 (
            .O(N__29633),
            .I(N__29622));
    LocalMux I__6538 (
            .O(N__29630),
            .I(N__29619));
    LocalMux I__6537 (
            .O(N__29627),
            .I(N__29616));
    LocalMux I__6536 (
            .O(N__29622),
            .I(N__29612));
    Span4Mux_v I__6535 (
            .O(N__29619),
            .I(N__29609));
    Span4Mux_v I__6534 (
            .O(N__29616),
            .I(N__29606));
    InMux I__6533 (
            .O(N__29615),
            .I(N__29603));
    Span4Mux_v I__6532 (
            .O(N__29612),
            .I(N__29600));
    Odrv4 I__6531 (
            .O(N__29609),
            .I(\b2v_inst.reg_ancho_1Z0Z_4 ));
    Odrv4 I__6530 (
            .O(N__29606),
            .I(\b2v_inst.reg_ancho_1Z0Z_4 ));
    LocalMux I__6529 (
            .O(N__29603),
            .I(\b2v_inst.reg_ancho_1Z0Z_4 ));
    Odrv4 I__6528 (
            .O(N__29600),
            .I(\b2v_inst.reg_ancho_1Z0Z_4 ));
    CascadeMux I__6527 (
            .O(N__29591),
            .I(N__29586));
    CascadeMux I__6526 (
            .O(N__29590),
            .I(N__29583));
    CascadeMux I__6525 (
            .O(N__29589),
            .I(N__29580));
    InMux I__6524 (
            .O(N__29586),
            .I(N__29577));
    InMux I__6523 (
            .O(N__29583),
            .I(N__29574));
    InMux I__6522 (
            .O(N__29580),
            .I(N__29571));
    LocalMux I__6521 (
            .O(N__29577),
            .I(N__29566));
    LocalMux I__6520 (
            .O(N__29574),
            .I(N__29566));
    LocalMux I__6519 (
            .O(N__29571),
            .I(\b2v_inst.reg_ancho_3_i_4 ));
    Odrv4 I__6518 (
            .O(N__29566),
            .I(\b2v_inst.reg_ancho_3_i_4 ));
    CascadeMux I__6517 (
            .O(N__29561),
            .I(N__29556));
    InMux I__6516 (
            .O(N__29560),
            .I(N__29553));
    InMux I__6515 (
            .O(N__29559),
            .I(N__29548));
    InMux I__6514 (
            .O(N__29556),
            .I(N__29545));
    LocalMux I__6513 (
            .O(N__29553),
            .I(N__29542));
    InMux I__6512 (
            .O(N__29552),
            .I(N__29539));
    InMux I__6511 (
            .O(N__29551),
            .I(N__29536));
    LocalMux I__6510 (
            .O(N__29548),
            .I(N__29533));
    LocalMux I__6509 (
            .O(N__29545),
            .I(N__29530));
    Span12Mux_h I__6508 (
            .O(N__29542),
            .I(N__29525));
    LocalMux I__6507 (
            .O(N__29539),
            .I(N__29525));
    LocalMux I__6506 (
            .O(N__29536),
            .I(N__29522));
    Odrv4 I__6505 (
            .O(N__29533),
            .I(\b2v_inst.reg_ancho_1Z0Z_5 ));
    Odrv4 I__6504 (
            .O(N__29530),
            .I(\b2v_inst.reg_ancho_1Z0Z_5 ));
    Odrv12 I__6503 (
            .O(N__29525),
            .I(\b2v_inst.reg_ancho_1Z0Z_5 ));
    Odrv4 I__6502 (
            .O(N__29522),
            .I(\b2v_inst.reg_ancho_1Z0Z_5 ));
    CascadeMux I__6501 (
            .O(N__29513),
            .I(N__29509));
    InMux I__6500 (
            .O(N__29512),
            .I(N__29506));
    InMux I__6499 (
            .O(N__29509),
            .I(N__29502));
    LocalMux I__6498 (
            .O(N__29506),
            .I(N__29499));
    InMux I__6497 (
            .O(N__29505),
            .I(N__29496));
    LocalMux I__6496 (
            .O(N__29502),
            .I(N__29493));
    Odrv4 I__6495 (
            .O(N__29499),
            .I(\b2v_inst.reg_ancho_3_i_5 ));
    LocalMux I__6494 (
            .O(N__29496),
            .I(\b2v_inst.reg_ancho_3_i_5 ));
    Odrv4 I__6493 (
            .O(N__29493),
            .I(\b2v_inst.reg_ancho_3_i_5 ));
    InMux I__6492 (
            .O(N__29486),
            .I(N__29481));
    InMux I__6491 (
            .O(N__29485),
            .I(N__29478));
    InMux I__6490 (
            .O(N__29484),
            .I(N__29475));
    LocalMux I__6489 (
            .O(N__29481),
            .I(N__29469));
    LocalMux I__6488 (
            .O(N__29478),
            .I(N__29469));
    LocalMux I__6487 (
            .O(N__29475),
            .I(N__29466));
    InMux I__6486 (
            .O(N__29474),
            .I(N__29462));
    Span4Mux_v I__6485 (
            .O(N__29469),
            .I(N__29457));
    Span4Mux_h I__6484 (
            .O(N__29466),
            .I(N__29457));
    InMux I__6483 (
            .O(N__29465),
            .I(N__29454));
    LocalMux I__6482 (
            .O(N__29462),
            .I(N__29451));
    Odrv4 I__6481 (
            .O(N__29457),
            .I(\b2v_inst.reg_ancho_1Z0Z_6 ));
    LocalMux I__6480 (
            .O(N__29454),
            .I(\b2v_inst.reg_ancho_1Z0Z_6 ));
    Odrv12 I__6479 (
            .O(N__29451),
            .I(\b2v_inst.reg_ancho_1Z0Z_6 ));
    InMux I__6478 (
            .O(N__29444),
            .I(N__29439));
    InMux I__6477 (
            .O(N__29443),
            .I(N__29436));
    InMux I__6476 (
            .O(N__29442),
            .I(N__29433));
    LocalMux I__6475 (
            .O(N__29439),
            .I(\b2v_inst.reg_ancho_3Z0Z_6 ));
    LocalMux I__6474 (
            .O(N__29436),
            .I(\b2v_inst.reg_ancho_3Z0Z_6 ));
    LocalMux I__6473 (
            .O(N__29433),
            .I(\b2v_inst.reg_ancho_3Z0Z_6 ));
    InMux I__6472 (
            .O(N__29426),
            .I(N__29421));
    CascadeMux I__6471 (
            .O(N__29425),
            .I(N__29418));
    CascadeMux I__6470 (
            .O(N__29424),
            .I(N__29415));
    LocalMux I__6469 (
            .O(N__29421),
            .I(N__29412));
    InMux I__6468 (
            .O(N__29418),
            .I(N__29409));
    InMux I__6467 (
            .O(N__29415),
            .I(N__29406));
    Span4Mux_h I__6466 (
            .O(N__29412),
            .I(N__29401));
    LocalMux I__6465 (
            .O(N__29409),
            .I(N__29401));
    LocalMux I__6464 (
            .O(N__29406),
            .I(\b2v_inst.reg_ancho_3_i_6 ));
    Odrv4 I__6463 (
            .O(N__29401),
            .I(\b2v_inst.reg_ancho_3_i_6 ));
    InMux I__6462 (
            .O(N__29396),
            .I(N__29392));
    CascadeMux I__6461 (
            .O(N__29395),
            .I(N__29387));
    LocalMux I__6460 (
            .O(N__29392),
            .I(N__29383));
    InMux I__6459 (
            .O(N__29391),
            .I(N__29380));
    InMux I__6458 (
            .O(N__29390),
            .I(N__29375));
    InMux I__6457 (
            .O(N__29387),
            .I(N__29375));
    InMux I__6456 (
            .O(N__29386),
            .I(N__29372));
    Span4Mux_h I__6455 (
            .O(N__29383),
            .I(N__29369));
    LocalMux I__6454 (
            .O(N__29380),
            .I(N__29366));
    LocalMux I__6453 (
            .O(N__29375),
            .I(N__29363));
    LocalMux I__6452 (
            .O(N__29372),
            .I(N__29360));
    Odrv4 I__6451 (
            .O(N__29369),
            .I(\b2v_inst.reg_ancho_1Z0Z_7 ));
    Odrv4 I__6450 (
            .O(N__29366),
            .I(\b2v_inst.reg_ancho_1Z0Z_7 ));
    Odrv12 I__6449 (
            .O(N__29363),
            .I(\b2v_inst.reg_ancho_1Z0Z_7 ));
    Odrv4 I__6448 (
            .O(N__29360),
            .I(\b2v_inst.reg_ancho_1Z0Z_7 ));
    InMux I__6447 (
            .O(N__29351),
            .I(N__29346));
    CascadeMux I__6446 (
            .O(N__29350),
            .I(N__29343));
    CascadeMux I__6445 (
            .O(N__29349),
            .I(N__29340));
    LocalMux I__6444 (
            .O(N__29346),
            .I(N__29337));
    InMux I__6443 (
            .O(N__29343),
            .I(N__29334));
    InMux I__6442 (
            .O(N__29340),
            .I(N__29331));
    Span4Mux_h I__6441 (
            .O(N__29337),
            .I(N__29326));
    LocalMux I__6440 (
            .O(N__29334),
            .I(N__29326));
    LocalMux I__6439 (
            .O(N__29331),
            .I(\b2v_inst.reg_ancho_3_i_7 ));
    Odrv4 I__6438 (
            .O(N__29326),
            .I(\b2v_inst.reg_ancho_3_i_7 ));
    CascadeMux I__6437 (
            .O(N__29321),
            .I(N__29316));
    InMux I__6436 (
            .O(N__29320),
            .I(N__29313));
    CascadeMux I__6435 (
            .O(N__29319),
            .I(N__29310));
    InMux I__6434 (
            .O(N__29316),
            .I(N__29307));
    LocalMux I__6433 (
            .O(N__29313),
            .I(N__29304));
    InMux I__6432 (
            .O(N__29310),
            .I(N__29301));
    LocalMux I__6431 (
            .O(N__29307),
            .I(N__29298));
    Odrv4 I__6430 (
            .O(N__29304),
            .I(\b2v_inst.reg_ancho_3_i_8 ));
    LocalMux I__6429 (
            .O(N__29301),
            .I(\b2v_inst.reg_ancho_3_i_8 ));
    Odrv4 I__6428 (
            .O(N__29298),
            .I(\b2v_inst.reg_ancho_3_i_8 ));
    CascadeMux I__6427 (
            .O(N__29291),
            .I(N__29287));
    CascadeMux I__6426 (
            .O(N__29290),
            .I(N__29283));
    InMux I__6425 (
            .O(N__29287),
            .I(N__29280));
    CascadeMux I__6424 (
            .O(N__29286),
            .I(N__29277));
    InMux I__6423 (
            .O(N__29283),
            .I(N__29274));
    LocalMux I__6422 (
            .O(N__29280),
            .I(N__29271));
    InMux I__6421 (
            .O(N__29277),
            .I(N__29268));
    LocalMux I__6420 (
            .O(N__29274),
            .I(N__29265));
    Odrv4 I__6419 (
            .O(N__29271),
            .I(\b2v_inst.reg_ancho_3_i_9 ));
    LocalMux I__6418 (
            .O(N__29268),
            .I(\b2v_inst.reg_ancho_3_i_9 ));
    Odrv4 I__6417 (
            .O(N__29265),
            .I(\b2v_inst.reg_ancho_3_i_9 ));
    InMux I__6416 (
            .O(N__29258),
            .I(N__29253));
    InMux I__6415 (
            .O(N__29257),
            .I(N__29250));
    InMux I__6414 (
            .O(N__29256),
            .I(N__29247));
    LocalMux I__6413 (
            .O(N__29253),
            .I(N__29240));
    LocalMux I__6412 (
            .O(N__29250),
            .I(N__29240));
    LocalMux I__6411 (
            .O(N__29247),
            .I(N__29237));
    InMux I__6410 (
            .O(N__29246),
            .I(N__29234));
    InMux I__6409 (
            .O(N__29245),
            .I(N__29231));
    Span4Mux_v I__6408 (
            .O(N__29240),
            .I(N__29228));
    Span4Mux_v I__6407 (
            .O(N__29237),
            .I(N__29225));
    LocalMux I__6406 (
            .O(N__29234),
            .I(N__29220));
    LocalMux I__6405 (
            .O(N__29231),
            .I(N__29220));
    Odrv4 I__6404 (
            .O(N__29228),
            .I(\b2v_inst.reg_ancho_1Z0Z_10 ));
    Odrv4 I__6403 (
            .O(N__29225),
            .I(\b2v_inst.reg_ancho_1Z0Z_10 ));
    Odrv4 I__6402 (
            .O(N__29220),
            .I(\b2v_inst.reg_ancho_1Z0Z_10 ));
    CascadeMux I__6401 (
            .O(N__29213),
            .I(N__29209));
    CascadeMux I__6400 (
            .O(N__29212),
            .I(N__29205));
    InMux I__6399 (
            .O(N__29209),
            .I(N__29202));
    CascadeMux I__6398 (
            .O(N__29208),
            .I(N__29199));
    InMux I__6397 (
            .O(N__29205),
            .I(N__29196));
    LocalMux I__6396 (
            .O(N__29202),
            .I(N__29193));
    InMux I__6395 (
            .O(N__29199),
            .I(N__29190));
    LocalMux I__6394 (
            .O(N__29196),
            .I(N__29187));
    Odrv4 I__6393 (
            .O(N__29193),
            .I(\b2v_inst.reg_ancho_3_i_10 ));
    LocalMux I__6392 (
            .O(N__29190),
            .I(\b2v_inst.reg_ancho_3_i_10 ));
    Odrv4 I__6391 (
            .O(N__29187),
            .I(\b2v_inst.reg_ancho_3_i_10 ));
    InMux I__6390 (
            .O(N__29180),
            .I(\b2v_inst.valor_max_final40 ));
    InMux I__6389 (
            .O(N__29177),
            .I(N__29174));
    LocalMux I__6388 (
            .O(N__29174),
            .I(N__29171));
    Span4Mux_v I__6387 (
            .O(N__29171),
            .I(N__29168));
    Odrv4 I__6386 (
            .O(N__29168),
            .I(\b2v_inst.valor_max_final40_THRU_CO ));
    InMux I__6385 (
            .O(N__29165),
            .I(\b2v_inst.un2_valor_max2 ));
    InMux I__6384 (
            .O(N__29162),
            .I(N__29159));
    LocalMux I__6383 (
            .O(N__29159),
            .I(N__29154));
    InMux I__6382 (
            .O(N__29158),
            .I(N__29150));
    InMux I__6381 (
            .O(N__29157),
            .I(N__29147));
    Span4Mux_v I__6380 (
            .O(N__29154),
            .I(N__29144));
    InMux I__6379 (
            .O(N__29153),
            .I(N__29141));
    LocalMux I__6378 (
            .O(N__29150),
            .I(N__29138));
    LocalMux I__6377 (
            .O(N__29147),
            .I(N__29135));
    Span4Mux_h I__6376 (
            .O(N__29144),
            .I(N__29130));
    LocalMux I__6375 (
            .O(N__29141),
            .I(N__29130));
    Span4Mux_v I__6374 (
            .O(N__29138),
            .I(N__29127));
    Odrv4 I__6373 (
            .O(N__29135),
            .I(\b2v_inst.reg_anteriorZ0Z_3 ));
    Odrv4 I__6372 (
            .O(N__29130),
            .I(\b2v_inst.reg_anteriorZ0Z_3 ));
    Odrv4 I__6371 (
            .O(N__29127),
            .I(\b2v_inst.reg_anteriorZ0Z_3 ));
    CascadeMux I__6370 (
            .O(N__29120),
            .I(N__29117));
    InMux I__6369 (
            .O(N__29117),
            .I(N__29114));
    LocalMux I__6368 (
            .O(N__29114),
            .I(N__29111));
    Span4Mux_v I__6367 (
            .O(N__29111),
            .I(N__29108));
    Odrv4 I__6366 (
            .O(N__29108),
            .I(\b2v_inst.data_a_escribir_RNO_0Z0Z_3 ));
    InMux I__6365 (
            .O(N__29105),
            .I(N__29102));
    LocalMux I__6364 (
            .O(N__29102),
            .I(N__29098));
    InMux I__6363 (
            .O(N__29101),
            .I(N__29094));
    Span4Mux_h I__6362 (
            .O(N__29098),
            .I(N__29091));
    InMux I__6361 (
            .O(N__29097),
            .I(N__29087));
    LocalMux I__6360 (
            .O(N__29094),
            .I(N__29084));
    Span4Mux_v I__6359 (
            .O(N__29091),
            .I(N__29081));
    InMux I__6358 (
            .O(N__29090),
            .I(N__29078));
    LocalMux I__6357 (
            .O(N__29087),
            .I(N__29073));
    Span4Mux_v I__6356 (
            .O(N__29084),
            .I(N__29073));
    Odrv4 I__6355 (
            .O(N__29081),
            .I(\b2v_inst.reg_anteriorZ0Z_5 ));
    LocalMux I__6354 (
            .O(N__29078),
            .I(\b2v_inst.reg_anteriorZ0Z_5 ));
    Odrv4 I__6353 (
            .O(N__29073),
            .I(\b2v_inst.reg_anteriorZ0Z_5 ));
    InMux I__6352 (
            .O(N__29066),
            .I(N__29062));
    InMux I__6351 (
            .O(N__29065),
            .I(N__29057));
    LocalMux I__6350 (
            .O(N__29062),
            .I(N__29054));
    InMux I__6349 (
            .O(N__29061),
            .I(N__29049));
    InMux I__6348 (
            .O(N__29060),
            .I(N__29049));
    LocalMux I__6347 (
            .O(N__29057),
            .I(N__29046));
    Span4Mux_v I__6346 (
            .O(N__29054),
            .I(N__29042));
    LocalMux I__6345 (
            .O(N__29049),
            .I(N__29039));
    Span4Mux_v I__6344 (
            .O(N__29046),
            .I(N__29036));
    InMux I__6343 (
            .O(N__29045),
            .I(N__29033));
    Odrv4 I__6342 (
            .O(N__29042),
            .I(\b2v_inst.reg_ancho_1Z0Z_0 ));
    Odrv12 I__6341 (
            .O(N__29039),
            .I(\b2v_inst.reg_ancho_1Z0Z_0 ));
    Odrv4 I__6340 (
            .O(N__29036),
            .I(\b2v_inst.reg_ancho_1Z0Z_0 ));
    LocalMux I__6339 (
            .O(N__29033),
            .I(\b2v_inst.reg_ancho_1Z0Z_0 ));
    CascadeMux I__6338 (
            .O(N__29024),
            .I(N__29019));
    InMux I__6337 (
            .O(N__29023),
            .I(N__29016));
    CascadeMux I__6336 (
            .O(N__29022),
            .I(N__29013));
    InMux I__6335 (
            .O(N__29019),
            .I(N__29010));
    LocalMux I__6334 (
            .O(N__29016),
            .I(N__29007));
    InMux I__6333 (
            .O(N__29013),
            .I(N__29004));
    LocalMux I__6332 (
            .O(N__29010),
            .I(N__29001));
    Odrv4 I__6331 (
            .O(N__29007),
            .I(\b2v_inst.reg_ancho_3_i_0 ));
    LocalMux I__6330 (
            .O(N__29004),
            .I(\b2v_inst.reg_ancho_3_i_0 ));
    Odrv4 I__6329 (
            .O(N__29001),
            .I(\b2v_inst.reg_ancho_3_i_0 ));
    InMux I__6328 (
            .O(N__28994),
            .I(N__28991));
    LocalMux I__6327 (
            .O(N__28991),
            .I(N__28987));
    InMux I__6326 (
            .O(N__28990),
            .I(N__28984));
    Span4Mux_v I__6325 (
            .O(N__28987),
            .I(N__28977));
    LocalMux I__6324 (
            .O(N__28984),
            .I(N__28977));
    InMux I__6323 (
            .O(N__28983),
            .I(N__28972));
    InMux I__6322 (
            .O(N__28982),
            .I(N__28972));
    Span4Mux_v I__6321 (
            .O(N__28977),
            .I(N__28968));
    LocalMux I__6320 (
            .O(N__28972),
            .I(N__28965));
    InMux I__6319 (
            .O(N__28971),
            .I(N__28962));
    Span4Mux_h I__6318 (
            .O(N__28968),
            .I(N__28959));
    Odrv12 I__6317 (
            .O(N__28965),
            .I(\b2v_inst.reg_ancho_1Z0Z_1 ));
    LocalMux I__6316 (
            .O(N__28962),
            .I(\b2v_inst.reg_ancho_1Z0Z_1 ));
    Odrv4 I__6315 (
            .O(N__28959),
            .I(\b2v_inst.reg_ancho_1Z0Z_1 ));
    CascadeMux I__6314 (
            .O(N__28952),
            .I(N__28948));
    CascadeMux I__6313 (
            .O(N__28951),
            .I(N__28945));
    InMux I__6312 (
            .O(N__28948),
            .I(N__28941));
    InMux I__6311 (
            .O(N__28945),
            .I(N__28938));
    CascadeMux I__6310 (
            .O(N__28944),
            .I(N__28935));
    LocalMux I__6309 (
            .O(N__28941),
            .I(N__28932));
    LocalMux I__6308 (
            .O(N__28938),
            .I(N__28929));
    InMux I__6307 (
            .O(N__28935),
            .I(N__28926));
    Span4Mux_h I__6306 (
            .O(N__28932),
            .I(N__28923));
    Odrv4 I__6305 (
            .O(N__28929),
            .I(\b2v_inst.reg_ancho_3_i_1 ));
    LocalMux I__6304 (
            .O(N__28926),
            .I(\b2v_inst.reg_ancho_3_i_1 ));
    Odrv4 I__6303 (
            .O(N__28923),
            .I(\b2v_inst.reg_ancho_3_i_1 ));
    CascadeMux I__6302 (
            .O(N__28916),
            .I(N__28912));
    CascadeMux I__6301 (
            .O(N__28915),
            .I(N__28908));
    InMux I__6300 (
            .O(N__28912),
            .I(N__28905));
    CascadeMux I__6299 (
            .O(N__28911),
            .I(N__28902));
    InMux I__6298 (
            .O(N__28908),
            .I(N__28899));
    LocalMux I__6297 (
            .O(N__28905),
            .I(N__28896));
    InMux I__6296 (
            .O(N__28902),
            .I(N__28893));
    LocalMux I__6295 (
            .O(N__28899),
            .I(N__28890));
    Odrv4 I__6294 (
            .O(N__28896),
            .I(\b2v_inst.reg_ancho_3_i_2 ));
    LocalMux I__6293 (
            .O(N__28893),
            .I(\b2v_inst.reg_ancho_3_i_2 ));
    Odrv4 I__6292 (
            .O(N__28890),
            .I(\b2v_inst.reg_ancho_3_i_2 ));
    CascadeMux I__6291 (
            .O(N__28883),
            .I(N__28878));
    InMux I__6290 (
            .O(N__28882),
            .I(N__28875));
    CascadeMux I__6289 (
            .O(N__28881),
            .I(N__28872));
    InMux I__6288 (
            .O(N__28878),
            .I(N__28869));
    LocalMux I__6287 (
            .O(N__28875),
            .I(N__28866));
    InMux I__6286 (
            .O(N__28872),
            .I(N__28863));
    LocalMux I__6285 (
            .O(N__28869),
            .I(N__28860));
    Odrv4 I__6284 (
            .O(N__28866),
            .I(\b2v_inst.reg_ancho_3_i_3 ));
    LocalMux I__6283 (
            .O(N__28863),
            .I(\b2v_inst.reg_ancho_3_i_3 ));
    Odrv4 I__6282 (
            .O(N__28860),
            .I(\b2v_inst.reg_ancho_3_i_3 ));
    InMux I__6281 (
            .O(N__28853),
            .I(N__28849));
    InMux I__6280 (
            .O(N__28852),
            .I(N__28846));
    LocalMux I__6279 (
            .O(N__28849),
            .I(SYNTHESIZED_WIRE_5_7));
    LocalMux I__6278 (
            .O(N__28846),
            .I(SYNTHESIZED_WIRE_5_7));
    InMux I__6277 (
            .O(N__28841),
            .I(N__28836));
    InMux I__6276 (
            .O(N__28840),
            .I(N__28833));
    InMux I__6275 (
            .O(N__28839),
            .I(N__28830));
    LocalMux I__6274 (
            .O(N__28836),
            .I(SYNTHESIZED_WIRE_5_6));
    LocalMux I__6273 (
            .O(N__28833),
            .I(SYNTHESIZED_WIRE_5_6));
    LocalMux I__6272 (
            .O(N__28830),
            .I(SYNTHESIZED_WIRE_5_6));
    InMux I__6271 (
            .O(N__28823),
            .I(N__28820));
    LocalMux I__6270 (
            .O(N__28820),
            .I(\b2v_inst.un12_pix_count_intlto7_N_3LZ0Z3 ));
    InMux I__6269 (
            .O(N__28817),
            .I(N__28814));
    LocalMux I__6268 (
            .O(N__28814),
            .I(N__28810));
    InMux I__6267 (
            .O(N__28813),
            .I(N__28807));
    Odrv12 I__6266 (
            .O(N__28810),
            .I(SYNTHESIZED_WIRE_10_5));
    LocalMux I__6265 (
            .O(N__28807),
            .I(SYNTHESIZED_WIRE_10_5));
    InMux I__6264 (
            .O(N__28802),
            .I(N__28799));
    LocalMux I__6263 (
            .O(N__28799),
            .I(N__28796));
    Span4Mux_h I__6262 (
            .O(N__28796),
            .I(N__28792));
    InMux I__6261 (
            .O(N__28795),
            .I(N__28789));
    Odrv4 I__6260 (
            .O(N__28792),
            .I(SYNTHESIZED_WIRE_5_5));
    LocalMux I__6259 (
            .O(N__28789),
            .I(SYNTHESIZED_WIRE_5_5));
    CEMux I__6258 (
            .O(N__28784),
            .I(N__28780));
    CEMux I__6257 (
            .O(N__28783),
            .I(N__28776));
    LocalMux I__6256 (
            .O(N__28780),
            .I(N__28773));
    CEMux I__6255 (
            .O(N__28779),
            .I(N__28770));
    LocalMux I__6254 (
            .O(N__28776),
            .I(N__28767));
    Span4Mux_v I__6253 (
            .O(N__28773),
            .I(N__28764));
    LocalMux I__6252 (
            .O(N__28770),
            .I(N__28761));
    Sp12to4 I__6251 (
            .O(N__28767),
            .I(N__28757));
    Span4Mux_h I__6250 (
            .O(N__28764),
            .I(N__28752));
    Span4Mux_h I__6249 (
            .O(N__28761),
            .I(N__28752));
    CascadeMux I__6248 (
            .O(N__28760),
            .I(N__28748));
    Span12Mux_h I__6247 (
            .O(N__28757),
            .I(N__28745));
    Span4Mux_h I__6246 (
            .O(N__28752),
            .I(N__28742));
    InMux I__6245 (
            .O(N__28751),
            .I(N__28739));
    InMux I__6244 (
            .O(N__28748),
            .I(N__28736));
    Odrv12 I__6243 (
            .O(N__28745),
            .I(\b2v_inst4.pix_count_int_0_sqmuxa ));
    Odrv4 I__6242 (
            .O(N__28742),
            .I(\b2v_inst4.pix_count_int_0_sqmuxa ));
    LocalMux I__6241 (
            .O(N__28739),
            .I(\b2v_inst4.pix_count_int_0_sqmuxa ));
    LocalMux I__6240 (
            .O(N__28736),
            .I(\b2v_inst4.pix_count_int_0_sqmuxa ));
    CascadeMux I__6239 (
            .O(N__28727),
            .I(N__28723));
    InMux I__6238 (
            .O(N__28726),
            .I(N__28720));
    InMux I__6237 (
            .O(N__28723),
            .I(N__28717));
    LocalMux I__6236 (
            .O(N__28720),
            .I(N__28712));
    LocalMux I__6235 (
            .O(N__28717),
            .I(N__28712));
    Odrv4 I__6234 (
            .O(N__28712),
            .I(\b2v_inst9.N_175_i ));
    InMux I__6233 (
            .O(N__28709),
            .I(N__28704));
    InMux I__6232 (
            .O(N__28708),
            .I(N__28699));
    InMux I__6231 (
            .O(N__28707),
            .I(N__28699));
    LocalMux I__6230 (
            .O(N__28704),
            .I(\b2v_inst9.bit_counterZ0Z_0 ));
    LocalMux I__6229 (
            .O(N__28699),
            .I(\b2v_inst9.bit_counterZ0Z_0 ));
    InMux I__6228 (
            .O(N__28694),
            .I(N__28689));
    InMux I__6227 (
            .O(N__28693),
            .I(N__28684));
    InMux I__6226 (
            .O(N__28692),
            .I(N__28684));
    LocalMux I__6225 (
            .O(N__28689),
            .I(\b2v_inst9.bit_counterZ1Z_1 ));
    LocalMux I__6224 (
            .O(N__28684),
            .I(\b2v_inst9.bit_counterZ1Z_1 ));
    InMux I__6223 (
            .O(N__28679),
            .I(\b2v_inst9.un1_bit_counter_3_cry_0 ));
    CascadeMux I__6222 (
            .O(N__28676),
            .I(N__28672));
    InMux I__6221 (
            .O(N__28675),
            .I(N__28668));
    InMux I__6220 (
            .O(N__28672),
            .I(N__28663));
    InMux I__6219 (
            .O(N__28671),
            .I(N__28663));
    LocalMux I__6218 (
            .O(N__28668),
            .I(\b2v_inst9.bit_counterZ0Z_2 ));
    LocalMux I__6217 (
            .O(N__28663),
            .I(\b2v_inst9.bit_counterZ0Z_2 ));
    InMux I__6216 (
            .O(N__28658),
            .I(\b2v_inst9.un1_bit_counter_3_cry_1 ));
    InMux I__6215 (
            .O(N__28655),
            .I(N__28647));
    InMux I__6214 (
            .O(N__28654),
            .I(N__28647));
    InMux I__6213 (
            .O(N__28653),
            .I(N__28642));
    InMux I__6212 (
            .O(N__28652),
            .I(N__28642));
    LocalMux I__6211 (
            .O(N__28647),
            .I(\b2v_inst9.fsm_state_RNIND1P1Z0Z_0 ));
    LocalMux I__6210 (
            .O(N__28642),
            .I(\b2v_inst9.fsm_state_RNIND1P1Z0Z_0 ));
    InMux I__6209 (
            .O(N__28637),
            .I(\b2v_inst9.un1_bit_counter_3_cry_2 ));
    InMux I__6208 (
            .O(N__28634),
            .I(N__28629));
    InMux I__6207 (
            .O(N__28633),
            .I(N__28624));
    InMux I__6206 (
            .O(N__28632),
            .I(N__28624));
    LocalMux I__6205 (
            .O(N__28629),
            .I(\b2v_inst9.bit_counterZ0Z_3 ));
    LocalMux I__6204 (
            .O(N__28624),
            .I(\b2v_inst9.bit_counterZ0Z_3 ));
    InMux I__6203 (
            .O(N__28619),
            .I(N__28616));
    LocalMux I__6202 (
            .O(N__28616),
            .I(N__28611));
    InMux I__6201 (
            .O(N__28615),
            .I(N__28607));
    InMux I__6200 (
            .O(N__28614),
            .I(N__28604));
    Span4Mux_h I__6199 (
            .O(N__28611),
            .I(N__28601));
    InMux I__6198 (
            .O(N__28610),
            .I(N__28598));
    LocalMux I__6197 (
            .O(N__28607),
            .I(\b2v_inst.reg_anteriorZ0Z_0 ));
    LocalMux I__6196 (
            .O(N__28604),
            .I(\b2v_inst.reg_anteriorZ0Z_0 ));
    Odrv4 I__6195 (
            .O(N__28601),
            .I(\b2v_inst.reg_anteriorZ0Z_0 ));
    LocalMux I__6194 (
            .O(N__28598),
            .I(\b2v_inst.reg_anteriorZ0Z_0 ));
    InMux I__6193 (
            .O(N__28589),
            .I(N__28585));
    InMux I__6192 (
            .O(N__28588),
            .I(N__28581));
    LocalMux I__6191 (
            .O(N__28585),
            .I(N__28578));
    InMux I__6190 (
            .O(N__28584),
            .I(N__28575));
    LocalMux I__6189 (
            .O(N__28581),
            .I(N__28571));
    Span4Mux_h I__6188 (
            .O(N__28578),
            .I(N__28566));
    LocalMux I__6187 (
            .O(N__28575),
            .I(N__28566));
    InMux I__6186 (
            .O(N__28574),
            .I(N__28563));
    Span4Mux_h I__6185 (
            .O(N__28571),
            .I(N__28558));
    Span4Mux_v I__6184 (
            .O(N__28566),
            .I(N__28558));
    LocalMux I__6183 (
            .O(N__28563),
            .I(\b2v_inst.reg_anteriorZ0Z_1 ));
    Odrv4 I__6182 (
            .O(N__28558),
            .I(\b2v_inst.reg_anteriorZ0Z_1 ));
    InMux I__6181 (
            .O(N__28553),
            .I(N__28550));
    LocalMux I__6180 (
            .O(N__28550),
            .I(N__28547));
    Span4Mux_v I__6179 (
            .O(N__28547),
            .I(N__28543));
    InMux I__6178 (
            .O(N__28546),
            .I(N__28540));
    Span4Mux_h I__6177 (
            .O(N__28543),
            .I(N__28537));
    LocalMux I__6176 (
            .O(N__28540),
            .I(N__28534));
    Odrv4 I__6175 (
            .O(N__28537),
            .I(\b2v_inst.N_654_2 ));
    Odrv4 I__6174 (
            .O(N__28534),
            .I(\b2v_inst.N_654_2 ));
    CascadeMux I__6173 (
            .O(N__28529),
            .I(\b2v_inst.un1_reset_inv_0_0_tz_cascade_ ));
    InMux I__6172 (
            .O(N__28526),
            .I(N__28522));
    InMux I__6171 (
            .O(N__28525),
            .I(N__28518));
    LocalMux I__6170 (
            .O(N__28522),
            .I(N__28515));
    InMux I__6169 (
            .O(N__28521),
            .I(N__28511));
    LocalMux I__6168 (
            .O(N__28518),
            .I(N__28508));
    Span4Mux_h I__6167 (
            .O(N__28515),
            .I(N__28505));
    InMux I__6166 (
            .O(N__28514),
            .I(N__28502));
    LocalMux I__6165 (
            .O(N__28511),
            .I(N__28497));
    Span12Mux_h I__6164 (
            .O(N__28508),
            .I(N__28497));
    Odrv4 I__6163 (
            .O(N__28505),
            .I(\b2v_inst.N_482 ));
    LocalMux I__6162 (
            .O(N__28502),
            .I(\b2v_inst.N_482 ));
    Odrv12 I__6161 (
            .O(N__28497),
            .I(\b2v_inst.N_482 ));
    CascadeMux I__6160 (
            .O(N__28490),
            .I(N__28487));
    InMux I__6159 (
            .O(N__28487),
            .I(N__28484));
    LocalMux I__6158 (
            .O(N__28484),
            .I(N__28481));
    Span4Mux_h I__6157 (
            .O(N__28481),
            .I(N__28477));
    InMux I__6156 (
            .O(N__28480),
            .I(N__28474));
    Odrv4 I__6155 (
            .O(N__28477),
            .I(\b2v_inst.eventosZ0Z_7 ));
    LocalMux I__6154 (
            .O(N__28474),
            .I(\b2v_inst.eventosZ0Z_7 ));
    InMux I__6153 (
            .O(N__28469),
            .I(N__28466));
    LocalMux I__6152 (
            .O(N__28466),
            .I(\b2v_inst.data_a_escribir_RNO_2Z0Z_7 ));
    InMux I__6151 (
            .O(N__28463),
            .I(\b2v_inst9.un1_cycle_counter_2_cry_0 ));
    InMux I__6150 (
            .O(N__28460),
            .I(\b2v_inst9.un1_cycle_counter_2_cry_1 ));
    InMux I__6149 (
            .O(N__28457),
            .I(\b2v_inst9.un1_cycle_counter_2_cry_2 ));
    CascadeMux I__6148 (
            .O(N__28454),
            .I(N__28449));
    InMux I__6147 (
            .O(N__28453),
            .I(N__28446));
    InMux I__6146 (
            .O(N__28452),
            .I(N__28441));
    InMux I__6145 (
            .O(N__28449),
            .I(N__28441));
    LocalMux I__6144 (
            .O(N__28446),
            .I(\b2v_inst9.cycle_counterZ0Z_3 ));
    LocalMux I__6143 (
            .O(N__28441),
            .I(\b2v_inst9.cycle_counterZ0Z_3 ));
    CascadeMux I__6142 (
            .O(N__28436),
            .I(\b2v_inst9.cycle_counter_RNIQAGDZ0Z_3_cascade_ ));
    InMux I__6141 (
            .O(N__28433),
            .I(N__28430));
    LocalMux I__6140 (
            .O(N__28430),
            .I(\b2v_inst9.un1_cycle_counter_2_cry_0_THRU_CO ));
    CascadeMux I__6139 (
            .O(N__28427),
            .I(N__28422));
    CascadeMux I__6138 (
            .O(N__28426),
            .I(N__28419));
    InMux I__6137 (
            .O(N__28425),
            .I(N__28409));
    InMux I__6136 (
            .O(N__28422),
            .I(N__28409));
    InMux I__6135 (
            .O(N__28419),
            .I(N__28409));
    InMux I__6134 (
            .O(N__28418),
            .I(N__28409));
    LocalMux I__6133 (
            .O(N__28409),
            .I(\b2v_inst9.cycle_counterZ0Z_1 ));
    CascadeMux I__6132 (
            .O(N__28406),
            .I(N__28402));
    CascadeMux I__6131 (
            .O(N__28405),
            .I(N__28399));
    InMux I__6130 (
            .O(N__28402),
            .I(N__28396));
    InMux I__6129 (
            .O(N__28399),
            .I(N__28393));
    LocalMux I__6128 (
            .O(N__28396),
            .I(N__28390));
    LocalMux I__6127 (
            .O(N__28393),
            .I(\b2v_inst.reg_anterior_i_9 ));
    Odrv4 I__6126 (
            .O(N__28390),
            .I(\b2v_inst.reg_anterior_i_9 ));
    CascadeMux I__6125 (
            .O(N__28385),
            .I(N__28381));
    CascadeMux I__6124 (
            .O(N__28384),
            .I(N__28378));
    InMux I__6123 (
            .O(N__28381),
            .I(N__28375));
    InMux I__6122 (
            .O(N__28378),
            .I(N__28372));
    LocalMux I__6121 (
            .O(N__28375),
            .I(N__28369));
    LocalMux I__6120 (
            .O(N__28372),
            .I(\b2v_inst.reg_anterior_i_10 ));
    Odrv4 I__6119 (
            .O(N__28369),
            .I(\b2v_inst.reg_anterior_i_10 ));
    InMux I__6118 (
            .O(N__28364),
            .I(N__28361));
    LocalMux I__6117 (
            .O(N__28361),
            .I(N__28358));
    Odrv4 I__6116 (
            .O(N__28358),
            .I(\b2v_inst.valor_max_final43_THRU_CO ));
    CascadeMux I__6115 (
            .O(N__28355),
            .I(N__28352));
    InMux I__6114 (
            .O(N__28352),
            .I(N__28349));
    LocalMux I__6113 (
            .O(N__28349),
            .I(N__28346));
    Odrv12 I__6112 (
            .O(N__28346),
            .I(\b2v_inst.m54_ns_1 ));
    InMux I__6111 (
            .O(N__28343),
            .I(\b2v_inst.valor_max_final41 ));
    InMux I__6110 (
            .O(N__28340),
            .I(N__28334));
    InMux I__6109 (
            .O(N__28339),
            .I(N__28328));
    InMux I__6108 (
            .O(N__28338),
            .I(N__28325));
    InMux I__6107 (
            .O(N__28337),
            .I(N__28322));
    LocalMux I__6106 (
            .O(N__28334),
            .I(N__28319));
    InMux I__6105 (
            .O(N__28333),
            .I(N__28314));
    InMux I__6104 (
            .O(N__28332),
            .I(N__28314));
    InMux I__6103 (
            .O(N__28331),
            .I(N__28310));
    LocalMux I__6102 (
            .O(N__28328),
            .I(N__28307));
    LocalMux I__6101 (
            .O(N__28325),
            .I(N__28304));
    LocalMux I__6100 (
            .O(N__28322),
            .I(N__28301));
    Span4Mux_h I__6099 (
            .O(N__28319),
            .I(N__28298));
    LocalMux I__6098 (
            .O(N__28314),
            .I(N__28294));
    InMux I__6097 (
            .O(N__28313),
            .I(N__28290));
    LocalMux I__6096 (
            .O(N__28310),
            .I(N__28287));
    Span4Mux_h I__6095 (
            .O(N__28307),
            .I(N__28282));
    Span4Mux_h I__6094 (
            .O(N__28304),
            .I(N__28282));
    Span4Mux_h I__6093 (
            .O(N__28301),
            .I(N__28277));
    Span4Mux_h I__6092 (
            .O(N__28298),
            .I(N__28277));
    InMux I__6091 (
            .O(N__28297),
            .I(N__28274));
    Span4Mux_h I__6090 (
            .O(N__28294),
            .I(N__28271));
    InMux I__6089 (
            .O(N__28293),
            .I(N__28268));
    LocalMux I__6088 (
            .O(N__28290),
            .I(\b2v_inst.stateZ0Z_6 ));
    Odrv12 I__6087 (
            .O(N__28287),
            .I(\b2v_inst.stateZ0Z_6 ));
    Odrv4 I__6086 (
            .O(N__28282),
            .I(\b2v_inst.stateZ0Z_6 ));
    Odrv4 I__6085 (
            .O(N__28277),
            .I(\b2v_inst.stateZ0Z_6 ));
    LocalMux I__6084 (
            .O(N__28274),
            .I(\b2v_inst.stateZ0Z_6 ));
    Odrv4 I__6083 (
            .O(N__28271),
            .I(\b2v_inst.stateZ0Z_6 ));
    LocalMux I__6082 (
            .O(N__28268),
            .I(\b2v_inst.stateZ0Z_6 ));
    InMux I__6081 (
            .O(N__28253),
            .I(N__28249));
    CascadeMux I__6080 (
            .O(N__28252),
            .I(N__28246));
    LocalMux I__6079 (
            .O(N__28249),
            .I(N__28243));
    InMux I__6078 (
            .O(N__28246),
            .I(N__28240));
    Span4Mux_h I__6077 (
            .O(N__28243),
            .I(N__28235));
    LocalMux I__6076 (
            .O(N__28240),
            .I(N__28230));
    InMux I__6075 (
            .O(N__28239),
            .I(N__28225));
    InMux I__6074 (
            .O(N__28238),
            .I(N__28225));
    Span4Mux_h I__6073 (
            .O(N__28235),
            .I(N__28222));
    InMux I__6072 (
            .O(N__28234),
            .I(N__28217));
    InMux I__6071 (
            .O(N__28233),
            .I(N__28217));
    Odrv4 I__6070 (
            .O(N__28230),
            .I(\b2v_inst.stateZ0Z_10 ));
    LocalMux I__6069 (
            .O(N__28225),
            .I(\b2v_inst.stateZ0Z_10 ));
    Odrv4 I__6068 (
            .O(N__28222),
            .I(\b2v_inst.stateZ0Z_10 ));
    LocalMux I__6067 (
            .O(N__28217),
            .I(\b2v_inst.stateZ0Z_10 ));
    InMux I__6066 (
            .O(N__28208),
            .I(N__28198));
    InMux I__6065 (
            .O(N__28207),
            .I(N__28192));
    InMux I__6064 (
            .O(N__28206),
            .I(N__28192));
    InMux I__6063 (
            .O(N__28205),
            .I(N__28189));
    InMux I__6062 (
            .O(N__28204),
            .I(N__28186));
    InMux I__6061 (
            .O(N__28203),
            .I(N__28178));
    InMux I__6060 (
            .O(N__28202),
            .I(N__28178));
    CascadeMux I__6059 (
            .O(N__28201),
            .I(N__28175));
    LocalMux I__6058 (
            .O(N__28198),
            .I(N__28170));
    InMux I__6057 (
            .O(N__28197),
            .I(N__28167));
    LocalMux I__6056 (
            .O(N__28192),
            .I(N__28164));
    LocalMux I__6055 (
            .O(N__28189),
            .I(N__28161));
    LocalMux I__6054 (
            .O(N__28186),
            .I(N__28158));
    InMux I__6053 (
            .O(N__28185),
            .I(N__28151));
    InMux I__6052 (
            .O(N__28184),
            .I(N__28151));
    InMux I__6051 (
            .O(N__28183),
            .I(N__28151));
    LocalMux I__6050 (
            .O(N__28178),
            .I(N__28148));
    InMux I__6049 (
            .O(N__28175),
            .I(N__28145));
    InMux I__6048 (
            .O(N__28174),
            .I(N__28142));
    InMux I__6047 (
            .O(N__28173),
            .I(N__28139));
    Span4Mux_v I__6046 (
            .O(N__28170),
            .I(N__28133));
    LocalMux I__6045 (
            .O(N__28167),
            .I(N__28130));
    Span4Mux_h I__6044 (
            .O(N__28164),
            .I(N__28127));
    Span4Mux_v I__6043 (
            .O(N__28161),
            .I(N__28116));
    Span4Mux_v I__6042 (
            .O(N__28158),
            .I(N__28116));
    LocalMux I__6041 (
            .O(N__28151),
            .I(N__28116));
    Span4Mux_h I__6040 (
            .O(N__28148),
            .I(N__28116));
    LocalMux I__6039 (
            .O(N__28145),
            .I(N__28116));
    LocalMux I__6038 (
            .O(N__28142),
            .I(N__28113));
    LocalMux I__6037 (
            .O(N__28139),
            .I(N__28110));
    InMux I__6036 (
            .O(N__28138),
            .I(N__28107));
    InMux I__6035 (
            .O(N__28137),
            .I(N__28102));
    InMux I__6034 (
            .O(N__28136),
            .I(N__28102));
    Span4Mux_h I__6033 (
            .O(N__28133),
            .I(N__28099));
    Span4Mux_h I__6032 (
            .O(N__28130),
            .I(N__28096));
    Span4Mux_h I__6031 (
            .O(N__28127),
            .I(N__28091));
    Span4Mux_h I__6030 (
            .O(N__28116),
            .I(N__28091));
    Odrv12 I__6029 (
            .O(N__28113),
            .I(\b2v_inst.stateZ0Z_29 ));
    Odrv4 I__6028 (
            .O(N__28110),
            .I(\b2v_inst.stateZ0Z_29 ));
    LocalMux I__6027 (
            .O(N__28107),
            .I(\b2v_inst.stateZ0Z_29 ));
    LocalMux I__6026 (
            .O(N__28102),
            .I(\b2v_inst.stateZ0Z_29 ));
    Odrv4 I__6025 (
            .O(N__28099),
            .I(\b2v_inst.stateZ0Z_29 ));
    Odrv4 I__6024 (
            .O(N__28096),
            .I(\b2v_inst.stateZ0Z_29 ));
    Odrv4 I__6023 (
            .O(N__28091),
            .I(\b2v_inst.stateZ0Z_29 ));
    InMux I__6022 (
            .O(N__28076),
            .I(N__28073));
    LocalMux I__6021 (
            .O(N__28073),
            .I(N__28070));
    Odrv4 I__6020 (
            .O(N__28070),
            .I(\b2v_inst.state_ns_a3_i_0_a2_1_4_1 ));
    CascadeMux I__6019 (
            .O(N__28067),
            .I(N__28061));
    InMux I__6018 (
            .O(N__28066),
            .I(N__28058));
    InMux I__6017 (
            .O(N__28065),
            .I(N__28053));
    InMux I__6016 (
            .O(N__28064),
            .I(N__28053));
    InMux I__6015 (
            .O(N__28061),
            .I(N__28050));
    LocalMux I__6014 (
            .O(N__28058),
            .I(N__28047));
    LocalMux I__6013 (
            .O(N__28053),
            .I(N__28040));
    LocalMux I__6012 (
            .O(N__28050),
            .I(N__28040));
    Span4Mux_h I__6011 (
            .O(N__28047),
            .I(N__28037));
    InMux I__6010 (
            .O(N__28046),
            .I(N__28032));
    InMux I__6009 (
            .O(N__28045),
            .I(N__28032));
    Odrv12 I__6008 (
            .O(N__28040),
            .I(b2v_inst_state_3));
    Odrv4 I__6007 (
            .O(N__28037),
            .I(b2v_inst_state_3));
    LocalMux I__6006 (
            .O(N__28032),
            .I(b2v_inst_state_3));
    InMux I__6005 (
            .O(N__28025),
            .I(N__28022));
    LocalMux I__6004 (
            .O(N__28022),
            .I(\b2v_inst.N_694 ));
    CascadeMux I__6003 (
            .O(N__28019),
            .I(\b2v_inst.N_695_cascade_ ));
    InMux I__6002 (
            .O(N__28016),
            .I(N__28013));
    LocalMux I__6001 (
            .O(N__28013),
            .I(N__28010));
    Span4Mux_h I__6000 (
            .O(N__28010),
            .I(N__28007));
    Odrv4 I__5999 (
            .O(N__28007),
            .I(\b2v_inst.state_ns_a3_i_0_1_1 ));
    InMux I__5998 (
            .O(N__28004),
            .I(N__27998));
    InMux I__5997 (
            .O(N__28003),
            .I(N__27998));
    LocalMux I__5996 (
            .O(N__27998),
            .I(N__27994));
    InMux I__5995 (
            .O(N__27997),
            .I(N__27990));
    Span4Mux_h I__5994 (
            .O(N__27994),
            .I(N__27987));
    InMux I__5993 (
            .O(N__27993),
            .I(N__27984));
    LocalMux I__5992 (
            .O(N__27990),
            .I(N__27980));
    Span4Mux_h I__5991 (
            .O(N__27987),
            .I(N__27975));
    LocalMux I__5990 (
            .O(N__27984),
            .I(N__27975));
    InMux I__5989 (
            .O(N__27983),
            .I(N__27972));
    Span4Mux_v I__5988 (
            .O(N__27980),
            .I(N__27967));
    Span4Mux_h I__5987 (
            .O(N__27975),
            .I(N__27967));
    LocalMux I__5986 (
            .O(N__27972),
            .I(\b2v_inst.un2_cuentalto10_i_a2_8 ));
    Odrv4 I__5985 (
            .O(N__27967),
            .I(\b2v_inst.un2_cuentalto10_i_a2_8 ));
    InMux I__5984 (
            .O(N__27962),
            .I(N__27954));
    InMux I__5983 (
            .O(N__27961),
            .I(N__27954));
    InMux I__5982 (
            .O(N__27960),
            .I(N__27951));
    InMux I__5981 (
            .O(N__27959),
            .I(N__27947));
    LocalMux I__5980 (
            .O(N__27954),
            .I(N__27944));
    LocalMux I__5979 (
            .O(N__27951),
            .I(N__27941));
    InMux I__5978 (
            .O(N__27950),
            .I(N__27938));
    LocalMux I__5977 (
            .O(N__27947),
            .I(N__27935));
    Span4Mux_h I__5976 (
            .O(N__27944),
            .I(N__27932));
    Span4Mux_v I__5975 (
            .O(N__27941),
            .I(N__27925));
    LocalMux I__5974 (
            .O(N__27938),
            .I(N__27925));
    Span4Mux_h I__5973 (
            .O(N__27935),
            .I(N__27925));
    Odrv4 I__5972 (
            .O(N__27932),
            .I(\b2v_inst.un2_cuentalto10_i_a2_7 ));
    Odrv4 I__5971 (
            .O(N__27925),
            .I(\b2v_inst.un2_cuentalto10_i_a2_7 ));
    CascadeMux I__5970 (
            .O(N__27920),
            .I(N__27914));
    InMux I__5969 (
            .O(N__27919),
            .I(N__27911));
    InMux I__5968 (
            .O(N__27918),
            .I(N__27902));
    InMux I__5967 (
            .O(N__27917),
            .I(N__27902));
    InMux I__5966 (
            .O(N__27914),
            .I(N__27902));
    LocalMux I__5965 (
            .O(N__27911),
            .I(N__27899));
    InMux I__5964 (
            .O(N__27910),
            .I(N__27896));
    CascadeMux I__5963 (
            .O(N__27909),
            .I(N__27893));
    LocalMux I__5962 (
            .O(N__27902),
            .I(N__27890));
    Span4Mux_h I__5961 (
            .O(N__27899),
            .I(N__27887));
    LocalMux I__5960 (
            .O(N__27896),
            .I(N__27883));
    InMux I__5959 (
            .O(N__27893),
            .I(N__27880));
    Span4Mux_v I__5958 (
            .O(N__27890),
            .I(N__27877));
    Span4Mux_v I__5957 (
            .O(N__27887),
            .I(N__27874));
    InMux I__5956 (
            .O(N__27886),
            .I(N__27871));
    Span4Mux_v I__5955 (
            .O(N__27883),
            .I(N__27866));
    LocalMux I__5954 (
            .O(N__27880),
            .I(N__27866));
    Sp12to4 I__5953 (
            .O(N__27877),
            .I(N__27859));
    Sp12to4 I__5952 (
            .O(N__27874),
            .I(N__27859));
    LocalMux I__5951 (
            .O(N__27871),
            .I(N__27859));
    Span4Mux_h I__5950 (
            .O(N__27866),
            .I(N__27856));
    Span12Mux_h I__5949 (
            .O(N__27859),
            .I(N__27853));
    Span4Mux_h I__5948 (
            .O(N__27856),
            .I(N__27850));
    Odrv12 I__5947 (
            .O(N__27853),
            .I(\b2v_inst.state_32_repZ0Z1 ));
    Odrv4 I__5946 (
            .O(N__27850),
            .I(\b2v_inst.state_32_repZ0Z1 ));
    CascadeMux I__5945 (
            .O(N__27845),
            .I(N__27841));
    InMux I__5944 (
            .O(N__27844),
            .I(N__27834));
    InMux I__5943 (
            .O(N__27841),
            .I(N__27830));
    InMux I__5942 (
            .O(N__27840),
            .I(N__27827));
    InMux I__5941 (
            .O(N__27839),
            .I(N__27822));
    InMux I__5940 (
            .O(N__27838),
            .I(N__27822));
    InMux I__5939 (
            .O(N__27837),
            .I(N__27819));
    LocalMux I__5938 (
            .O(N__27834),
            .I(N__27816));
    InMux I__5937 (
            .O(N__27833),
            .I(N__27813));
    LocalMux I__5936 (
            .O(N__27830),
            .I(N__27808));
    LocalMux I__5935 (
            .O(N__27827),
            .I(N__27808));
    LocalMux I__5934 (
            .O(N__27822),
            .I(N__27805));
    LocalMux I__5933 (
            .O(N__27819),
            .I(N__27802));
    Span4Mux_v I__5932 (
            .O(N__27816),
            .I(N__27799));
    LocalMux I__5931 (
            .O(N__27813),
            .I(N__27796));
    Span4Mux_v I__5930 (
            .O(N__27808),
            .I(N__27793));
    Span4Mux_h I__5929 (
            .O(N__27805),
            .I(N__27788));
    Span4Mux_v I__5928 (
            .O(N__27802),
            .I(N__27788));
    Span4Mux_v I__5927 (
            .O(N__27799),
            .I(N__27782));
    Span4Mux_v I__5926 (
            .O(N__27796),
            .I(N__27782));
    Span4Mux_v I__5925 (
            .O(N__27793),
            .I(N__27779));
    Span4Mux_h I__5924 (
            .O(N__27788),
            .I(N__27776));
    InMux I__5923 (
            .O(N__27787),
            .I(N__27773));
    Sp12to4 I__5922 (
            .O(N__27782),
            .I(N__27768));
    Sp12to4 I__5921 (
            .O(N__27779),
            .I(N__27768));
    Span4Mux_h I__5920 (
            .O(N__27776),
            .I(N__27763));
    LocalMux I__5919 (
            .O(N__27773),
            .I(N__27763));
    Span12Mux_h I__5918 (
            .O(N__27768),
            .I(N__27760));
    Sp12to4 I__5917 (
            .O(N__27763),
            .I(N__27757));
    Span12Mux_v I__5916 (
            .O(N__27760),
            .I(N__27754));
    Span12Mux_v I__5915 (
            .O(N__27757),
            .I(N__27751));
    Odrv12 I__5914 (
            .O(N__27754),
            .I(reset_c));
    Odrv12 I__5913 (
            .O(N__27751),
            .I(reset_c));
    CascadeMux I__5912 (
            .O(N__27746),
            .I(N__27742));
    InMux I__5911 (
            .O(N__27745),
            .I(N__27739));
    InMux I__5910 (
            .O(N__27742),
            .I(N__27736));
    LocalMux I__5909 (
            .O(N__27739),
            .I(N__27733));
    LocalMux I__5908 (
            .O(N__27736),
            .I(\b2v_inst.reg_anterior_i_1 ));
    Odrv4 I__5907 (
            .O(N__27733),
            .I(\b2v_inst.reg_anterior_i_1 ));
    CascadeMux I__5906 (
            .O(N__27728),
            .I(N__27724));
    InMux I__5905 (
            .O(N__27727),
            .I(N__27721));
    InMux I__5904 (
            .O(N__27724),
            .I(N__27718));
    LocalMux I__5903 (
            .O(N__27721),
            .I(N__27715));
    LocalMux I__5902 (
            .O(N__27718),
            .I(\b2v_inst.reg_anterior_i_2 ));
    Odrv4 I__5901 (
            .O(N__27715),
            .I(\b2v_inst.reg_anterior_i_2 ));
    CascadeMux I__5900 (
            .O(N__27710),
            .I(N__27706));
    InMux I__5899 (
            .O(N__27709),
            .I(N__27703));
    InMux I__5898 (
            .O(N__27706),
            .I(N__27700));
    LocalMux I__5897 (
            .O(N__27703),
            .I(N__27697));
    LocalMux I__5896 (
            .O(N__27700),
            .I(\b2v_inst.reg_anterior_i_3 ));
    Odrv4 I__5895 (
            .O(N__27697),
            .I(\b2v_inst.reg_anterior_i_3 ));
    CascadeMux I__5894 (
            .O(N__27692),
            .I(N__27688));
    CascadeMux I__5893 (
            .O(N__27691),
            .I(N__27685));
    InMux I__5892 (
            .O(N__27688),
            .I(N__27682));
    InMux I__5891 (
            .O(N__27685),
            .I(N__27679));
    LocalMux I__5890 (
            .O(N__27682),
            .I(N__27676));
    LocalMux I__5889 (
            .O(N__27679),
            .I(\b2v_inst.reg_anterior_i_4 ));
    Odrv4 I__5888 (
            .O(N__27676),
            .I(\b2v_inst.reg_anterior_i_4 ));
    CascadeMux I__5887 (
            .O(N__27671),
            .I(N__27667));
    CascadeMux I__5886 (
            .O(N__27670),
            .I(N__27664));
    InMux I__5885 (
            .O(N__27667),
            .I(N__27661));
    InMux I__5884 (
            .O(N__27664),
            .I(N__27658));
    LocalMux I__5883 (
            .O(N__27661),
            .I(N__27655));
    LocalMux I__5882 (
            .O(N__27658),
            .I(\b2v_inst.reg_anterior_i_5 ));
    Odrv4 I__5881 (
            .O(N__27655),
            .I(\b2v_inst.reg_anterior_i_5 ));
    CascadeMux I__5880 (
            .O(N__27650),
            .I(N__27646));
    InMux I__5879 (
            .O(N__27649),
            .I(N__27643));
    InMux I__5878 (
            .O(N__27646),
            .I(N__27640));
    LocalMux I__5877 (
            .O(N__27643),
            .I(N__27637));
    LocalMux I__5876 (
            .O(N__27640),
            .I(\b2v_inst.reg_anterior_i_6 ));
    Odrv4 I__5875 (
            .O(N__27637),
            .I(\b2v_inst.reg_anterior_i_6 ));
    CascadeMux I__5874 (
            .O(N__27632),
            .I(N__27628));
    CascadeMux I__5873 (
            .O(N__27631),
            .I(N__27625));
    InMux I__5872 (
            .O(N__27628),
            .I(N__27622));
    InMux I__5871 (
            .O(N__27625),
            .I(N__27619));
    LocalMux I__5870 (
            .O(N__27622),
            .I(N__27616));
    LocalMux I__5869 (
            .O(N__27619),
            .I(\b2v_inst.reg_anterior_i_7 ));
    Odrv4 I__5868 (
            .O(N__27616),
            .I(\b2v_inst.reg_anterior_i_7 ));
    CascadeMux I__5867 (
            .O(N__27611),
            .I(N__27607));
    CascadeMux I__5866 (
            .O(N__27610),
            .I(N__27604));
    InMux I__5865 (
            .O(N__27607),
            .I(N__27601));
    InMux I__5864 (
            .O(N__27604),
            .I(N__27598));
    LocalMux I__5863 (
            .O(N__27601),
            .I(N__27595));
    LocalMux I__5862 (
            .O(N__27598),
            .I(\b2v_inst.reg_anterior_i_8 ));
    Odrv4 I__5861 (
            .O(N__27595),
            .I(\b2v_inst.reg_anterior_i_8 ));
    CascadeMux I__5860 (
            .O(N__27590),
            .I(N__27587));
    InMux I__5859 (
            .O(N__27587),
            .I(N__27582));
    InMux I__5858 (
            .O(N__27586),
            .I(N__27579));
    InMux I__5857 (
            .O(N__27585),
            .I(N__27576));
    LocalMux I__5856 (
            .O(N__27582),
            .I(N__27572));
    LocalMux I__5855 (
            .O(N__27579),
            .I(N__27569));
    LocalMux I__5854 (
            .O(N__27576),
            .I(N__27566));
    InMux I__5853 (
            .O(N__27575),
            .I(N__27563));
    Span4Mux_h I__5852 (
            .O(N__27572),
            .I(N__27559));
    Span4Mux_v I__5851 (
            .O(N__27569),
            .I(N__27552));
    Span4Mux_h I__5850 (
            .O(N__27566),
            .I(N__27552));
    LocalMux I__5849 (
            .O(N__27563),
            .I(N__27552));
    InMux I__5848 (
            .O(N__27562),
            .I(N__27549));
    Odrv4 I__5847 (
            .O(N__27559),
            .I(\b2v_inst.reg_ancho_2Z0Z_7 ));
    Odrv4 I__5846 (
            .O(N__27552),
            .I(\b2v_inst.reg_ancho_2Z0Z_7 ));
    LocalMux I__5845 (
            .O(N__27549),
            .I(\b2v_inst.reg_ancho_2Z0Z_7 ));
    InMux I__5844 (
            .O(N__27542),
            .I(\b2v_inst.valor_max_final43 ));
    InMux I__5843 (
            .O(N__27539),
            .I(N__27536));
    LocalMux I__5842 (
            .O(N__27536),
            .I(\b2v_inst.data_a_escribir_RNO_0Z0Z_0 ));
    InMux I__5841 (
            .O(N__27533),
            .I(N__27530));
    LocalMux I__5840 (
            .O(N__27530),
            .I(\b2v_inst.data_a_escribir_RNO_0Z0Z_1 ));
    InMux I__5839 (
            .O(N__27527),
            .I(N__27524));
    LocalMux I__5838 (
            .O(N__27524),
            .I(N__27521));
    Span4Mux_v I__5837 (
            .O(N__27521),
            .I(N__27517));
    InMux I__5836 (
            .O(N__27520),
            .I(N__27514));
    Sp12to4 I__5835 (
            .O(N__27517),
            .I(N__27511));
    LocalMux I__5834 (
            .O(N__27514),
            .I(\b2v_inst.eventosZ0Z_5 ));
    Odrv12 I__5833 (
            .O(N__27511),
            .I(\b2v_inst.eventosZ0Z_5 ));
    CascadeMux I__5832 (
            .O(N__27506),
            .I(N__27502));
    InMux I__5831 (
            .O(N__27505),
            .I(N__27499));
    InMux I__5830 (
            .O(N__27502),
            .I(N__27496));
    LocalMux I__5829 (
            .O(N__27499),
            .I(N__27493));
    LocalMux I__5828 (
            .O(N__27496),
            .I(\b2v_inst.reg_anterior_i_0 ));
    Odrv4 I__5827 (
            .O(N__27493),
            .I(\b2v_inst.reg_anterior_i_0 ));
    InMux I__5826 (
            .O(N__27488),
            .I(N__27483));
    InMux I__5825 (
            .O(N__27487),
            .I(N__27480));
    InMux I__5824 (
            .O(N__27486),
            .I(N__27476));
    LocalMux I__5823 (
            .O(N__27483),
            .I(N__27471));
    LocalMux I__5822 (
            .O(N__27480),
            .I(N__27471));
    InMux I__5821 (
            .O(N__27479),
            .I(N__27468));
    LocalMux I__5820 (
            .O(N__27476),
            .I(N__27465));
    Span4Mux_v I__5819 (
            .O(N__27471),
            .I(N__27460));
    LocalMux I__5818 (
            .O(N__27468),
            .I(N__27460));
    Span4Mux_v I__5817 (
            .O(N__27465),
            .I(N__27455));
    Span4Mux_h I__5816 (
            .O(N__27460),
            .I(N__27455));
    Span4Mux_h I__5815 (
            .O(N__27455),
            .I(N__27452));
    Odrv4 I__5814 (
            .O(N__27452),
            .I(SYNTHESIZED_WIRE_3_0));
    InMux I__5813 (
            .O(N__27449),
            .I(N__27445));
    CascadeMux I__5812 (
            .O(N__27448),
            .I(N__27442));
    LocalMux I__5811 (
            .O(N__27445),
            .I(N__27438));
    InMux I__5810 (
            .O(N__27442),
            .I(N__27435));
    CascadeMux I__5809 (
            .O(N__27441),
            .I(N__27431));
    Span4Mux_v I__5808 (
            .O(N__27438),
            .I(N__27425));
    LocalMux I__5807 (
            .O(N__27435),
            .I(N__27425));
    CascadeMux I__5806 (
            .O(N__27434),
            .I(N__27422));
    InMux I__5805 (
            .O(N__27431),
            .I(N__27419));
    InMux I__5804 (
            .O(N__27430),
            .I(N__27416));
    Span4Mux_v I__5803 (
            .O(N__27425),
            .I(N__27413));
    InMux I__5802 (
            .O(N__27422),
            .I(N__27410));
    LocalMux I__5801 (
            .O(N__27419),
            .I(N__27405));
    LocalMux I__5800 (
            .O(N__27416),
            .I(N__27405));
    Odrv4 I__5799 (
            .O(N__27413),
            .I(\b2v_inst.reg_ancho_2Z0Z_0 ));
    LocalMux I__5798 (
            .O(N__27410),
            .I(\b2v_inst.reg_ancho_2Z0Z_0 ));
    Odrv4 I__5797 (
            .O(N__27405),
            .I(\b2v_inst.reg_ancho_2Z0Z_0 ));
    InMux I__5796 (
            .O(N__27398),
            .I(N__27395));
    LocalMux I__5795 (
            .O(N__27395),
            .I(N__27390));
    CascadeMux I__5794 (
            .O(N__27394),
            .I(N__27387));
    InMux I__5793 (
            .O(N__27393),
            .I(N__27384));
    Span4Mux_v I__5792 (
            .O(N__27390),
            .I(N__27380));
    InMux I__5791 (
            .O(N__27387),
            .I(N__27377));
    LocalMux I__5790 (
            .O(N__27384),
            .I(N__27374));
    InMux I__5789 (
            .O(N__27383),
            .I(N__27371));
    Span4Mux_h I__5788 (
            .O(N__27380),
            .I(N__27365));
    LocalMux I__5787 (
            .O(N__27377),
            .I(N__27365));
    Span4Mux_h I__5786 (
            .O(N__27374),
            .I(N__27360));
    LocalMux I__5785 (
            .O(N__27371),
            .I(N__27360));
    InMux I__5784 (
            .O(N__27370),
            .I(N__27357));
    Odrv4 I__5783 (
            .O(N__27365),
            .I(\b2v_inst.reg_ancho_2Z0Z_5 ));
    Odrv4 I__5782 (
            .O(N__27360),
            .I(\b2v_inst.reg_ancho_2Z0Z_5 ));
    LocalMux I__5781 (
            .O(N__27357),
            .I(\b2v_inst.reg_ancho_2Z0Z_5 ));
    InMux I__5780 (
            .O(N__27350),
            .I(N__27345));
    CascadeMux I__5779 (
            .O(N__27349),
            .I(N__27342));
    CascadeMux I__5778 (
            .O(N__27348),
            .I(N__27339));
    LocalMux I__5777 (
            .O(N__27345),
            .I(N__27336));
    InMux I__5776 (
            .O(N__27342),
            .I(N__27333));
    InMux I__5775 (
            .O(N__27339),
            .I(N__27330));
    Span4Mux_h I__5774 (
            .O(N__27336),
            .I(N__27327));
    LocalMux I__5773 (
            .O(N__27333),
            .I(N__27324));
    LocalMux I__5772 (
            .O(N__27330),
            .I(N__27321));
    Span4Mux_v I__5771 (
            .O(N__27327),
            .I(N__27312));
    Span4Mux_v I__5770 (
            .O(N__27324),
            .I(N__27312));
    Span4Mux_v I__5769 (
            .O(N__27321),
            .I(N__27312));
    InMux I__5768 (
            .O(N__27320),
            .I(N__27309));
    InMux I__5767 (
            .O(N__27319),
            .I(N__27306));
    Odrv4 I__5766 (
            .O(N__27312),
            .I(\b2v_inst.reg_ancho_2Z0Z_6 ));
    LocalMux I__5765 (
            .O(N__27309),
            .I(\b2v_inst.reg_ancho_2Z0Z_6 ));
    LocalMux I__5764 (
            .O(N__27306),
            .I(\b2v_inst.reg_ancho_2Z0Z_6 ));
    InMux I__5763 (
            .O(N__27299),
            .I(\b2v_inst.valor_max_final42 ));
    InMux I__5762 (
            .O(N__27296),
            .I(N__27293));
    LocalMux I__5761 (
            .O(N__27293),
            .I(N__27290));
    Span4Mux_h I__5760 (
            .O(N__27290),
            .I(N__27287));
    Odrv4 I__5759 (
            .O(N__27287),
            .I(\b2v_inst.data_a_escribir11_7_and ));
    InMux I__5758 (
            .O(N__27284),
            .I(N__27280));
    InMux I__5757 (
            .O(N__27283),
            .I(N__27277));
    LocalMux I__5756 (
            .O(N__27280),
            .I(N__27271));
    LocalMux I__5755 (
            .O(N__27277),
            .I(N__27271));
    InMux I__5754 (
            .O(N__27276),
            .I(N__27267));
    Span4Mux_v I__5753 (
            .O(N__27271),
            .I(N__27264));
    InMux I__5752 (
            .O(N__27270),
            .I(N__27261));
    LocalMux I__5751 (
            .O(N__27267),
            .I(N__27254));
    Sp12to4 I__5750 (
            .O(N__27264),
            .I(N__27254));
    LocalMux I__5749 (
            .O(N__27261),
            .I(N__27254));
    Odrv12 I__5748 (
            .O(N__27254),
            .I(SYNTHESIZED_WIRE_3_7));
    InMux I__5747 (
            .O(N__27251),
            .I(N__27245));
    InMux I__5746 (
            .O(N__27250),
            .I(N__27242));
    InMux I__5745 (
            .O(N__27249),
            .I(N__27239));
    InMux I__5744 (
            .O(N__27248),
            .I(N__27236));
    LocalMux I__5743 (
            .O(N__27245),
            .I(N__27233));
    LocalMux I__5742 (
            .O(N__27242),
            .I(N__27228));
    LocalMux I__5741 (
            .O(N__27239),
            .I(N__27228));
    LocalMux I__5740 (
            .O(N__27236),
            .I(N__27225));
    Span4Mux_v I__5739 (
            .O(N__27233),
            .I(N__27222));
    Span4Mux_v I__5738 (
            .O(N__27228),
            .I(N__27217));
    Span4Mux_h I__5737 (
            .O(N__27225),
            .I(N__27217));
    Span4Mux_h I__5736 (
            .O(N__27222),
            .I(N__27214));
    Span4Mux_h I__5735 (
            .O(N__27217),
            .I(N__27211));
    Odrv4 I__5734 (
            .O(N__27214),
            .I(SYNTHESIZED_WIRE_3_8));
    Odrv4 I__5733 (
            .O(N__27211),
            .I(SYNTHESIZED_WIRE_3_8));
    CascadeMux I__5732 (
            .O(N__27206),
            .I(N__27200));
    CascadeMux I__5731 (
            .O(N__27205),
            .I(N__27197));
    CascadeMux I__5730 (
            .O(N__27204),
            .I(N__27193));
    InMux I__5729 (
            .O(N__27203),
            .I(N__27183));
    InMux I__5728 (
            .O(N__27200),
            .I(N__27183));
    InMux I__5727 (
            .O(N__27197),
            .I(N__27179));
    InMux I__5726 (
            .O(N__27196),
            .I(N__27174));
    InMux I__5725 (
            .O(N__27193),
            .I(N__27174));
    InMux I__5724 (
            .O(N__27192),
            .I(N__27171));
    InMux I__5723 (
            .O(N__27191),
            .I(N__27168));
    InMux I__5722 (
            .O(N__27190),
            .I(N__27163));
    InMux I__5721 (
            .O(N__27189),
            .I(N__27163));
    CascadeMux I__5720 (
            .O(N__27188),
            .I(N__27159));
    LocalMux I__5719 (
            .O(N__27183),
            .I(N__27156));
    CascadeMux I__5718 (
            .O(N__27182),
            .I(N__27153));
    LocalMux I__5717 (
            .O(N__27179),
            .I(N__27150));
    LocalMux I__5716 (
            .O(N__27174),
            .I(N__27147));
    LocalMux I__5715 (
            .O(N__27171),
            .I(N__27143));
    LocalMux I__5714 (
            .O(N__27168),
            .I(N__27138));
    LocalMux I__5713 (
            .O(N__27163),
            .I(N__27138));
    InMux I__5712 (
            .O(N__27162),
            .I(N__27133));
    InMux I__5711 (
            .O(N__27159),
            .I(N__27133));
    Span4Mux_h I__5710 (
            .O(N__27156),
            .I(N__27130));
    InMux I__5709 (
            .O(N__27153),
            .I(N__27127));
    Span4Mux_v I__5708 (
            .O(N__27150),
            .I(N__27122));
    Span4Mux_v I__5707 (
            .O(N__27147),
            .I(N__27122));
    InMux I__5706 (
            .O(N__27146),
            .I(N__27119));
    Odrv12 I__5705 (
            .O(N__27143),
            .I(\b2v_inst9.fsm_stateZ0Z_1 ));
    Odrv4 I__5704 (
            .O(N__27138),
            .I(\b2v_inst9.fsm_stateZ0Z_1 ));
    LocalMux I__5703 (
            .O(N__27133),
            .I(\b2v_inst9.fsm_stateZ0Z_1 ));
    Odrv4 I__5702 (
            .O(N__27130),
            .I(\b2v_inst9.fsm_stateZ0Z_1 ));
    LocalMux I__5701 (
            .O(N__27127),
            .I(\b2v_inst9.fsm_stateZ0Z_1 ));
    Odrv4 I__5700 (
            .O(N__27122),
            .I(\b2v_inst9.fsm_stateZ0Z_1 ));
    LocalMux I__5699 (
            .O(N__27119),
            .I(\b2v_inst9.fsm_stateZ0Z_1 ));
    CascadeMux I__5698 (
            .O(N__27104),
            .I(\b2v_inst9.N_84_2_cascade_ ));
    InMux I__5697 (
            .O(N__27101),
            .I(N__27098));
    LocalMux I__5696 (
            .O(N__27098),
            .I(N__27094));
    InMux I__5695 (
            .O(N__27097),
            .I(N__27091));
    Odrv4 I__5694 (
            .O(N__27094),
            .I(\b2v_inst9.N_582 ));
    LocalMux I__5693 (
            .O(N__27091),
            .I(\b2v_inst9.N_582 ));
    InMux I__5692 (
            .O(N__27086),
            .I(N__27083));
    LocalMux I__5691 (
            .O(N__27083),
            .I(N__27080));
    Span4Mux_v I__5690 (
            .O(N__27080),
            .I(N__27077));
    Sp12to4 I__5689 (
            .O(N__27077),
            .I(N__27074));
    Span12Mux_h I__5688 (
            .O(N__27074),
            .I(N__27070));
    InMux I__5687 (
            .O(N__27073),
            .I(N__27067));
    Odrv12 I__5686 (
            .O(N__27070),
            .I(SYNTHESIZED_WIRE_5_4));
    LocalMux I__5685 (
            .O(N__27067),
            .I(SYNTHESIZED_WIRE_5_4));
    CascadeMux I__5684 (
            .O(N__27062),
            .I(\b2v_inst.un12_pix_count_intlto7_N_2LZ0Z1_cascade_ ));
    InMux I__5683 (
            .O(N__27059),
            .I(N__27055));
    InMux I__5682 (
            .O(N__27058),
            .I(N__27052));
    LocalMux I__5681 (
            .O(N__27055),
            .I(N__27049));
    LocalMux I__5680 (
            .O(N__27052),
            .I(N__27046));
    Span4Mux_h I__5679 (
            .O(N__27049),
            .I(N__27043));
    Span4Mux_v I__5678 (
            .O(N__27046),
            .I(N__27040));
    Span4Mux_v I__5677 (
            .O(N__27043),
            .I(N__27035));
    Span4Mux_h I__5676 (
            .O(N__27040),
            .I(N__27035));
    Odrv4 I__5675 (
            .O(N__27035),
            .I(\b2v_inst.un13_pix_count_int_li_0 ));
    CascadeMux I__5674 (
            .O(N__27032),
            .I(\b2v_inst.un13_pix_count_int_li_0_cascade_ ));
    InMux I__5673 (
            .O(N__27029),
            .I(N__27026));
    LocalMux I__5672 (
            .O(N__27026),
            .I(N__27023));
    Span4Mux_v I__5671 (
            .O(N__27023),
            .I(N__27019));
    CascadeMux I__5670 (
            .O(N__27022),
            .I(N__27015));
    Sp12to4 I__5669 (
            .O(N__27019),
            .I(N__27012));
    InMux I__5668 (
            .O(N__27018),
            .I(N__27009));
    InMux I__5667 (
            .O(N__27015),
            .I(N__27006));
    Odrv12 I__5666 (
            .O(N__27012),
            .I(SYNTHESIZED_WIRE_10_1));
    LocalMux I__5665 (
            .O(N__27009),
            .I(SYNTHESIZED_WIRE_10_1));
    LocalMux I__5664 (
            .O(N__27006),
            .I(SYNTHESIZED_WIRE_10_1));
    InMux I__5663 (
            .O(N__26999),
            .I(N__26995));
    InMux I__5662 (
            .O(N__26998),
            .I(N__26992));
    LocalMux I__5661 (
            .O(N__26995),
            .I(SYNTHESIZED_WIRE_5_1));
    LocalMux I__5660 (
            .O(N__26992),
            .I(SYNTHESIZED_WIRE_5_1));
    InMux I__5659 (
            .O(N__26987),
            .I(N__26983));
    CascadeMux I__5658 (
            .O(N__26986),
            .I(N__26979));
    LocalMux I__5657 (
            .O(N__26983),
            .I(N__26976));
    InMux I__5656 (
            .O(N__26982),
            .I(N__26971));
    InMux I__5655 (
            .O(N__26979),
            .I(N__26971));
    Odrv12 I__5654 (
            .O(N__26976),
            .I(SYNTHESIZED_WIRE_10_2));
    LocalMux I__5653 (
            .O(N__26971),
            .I(SYNTHESIZED_WIRE_10_2));
    InMux I__5652 (
            .O(N__26966),
            .I(N__26962));
    InMux I__5651 (
            .O(N__26965),
            .I(N__26959));
    LocalMux I__5650 (
            .O(N__26962),
            .I(SYNTHESIZED_WIRE_5_2));
    LocalMux I__5649 (
            .O(N__26959),
            .I(SYNTHESIZED_WIRE_5_2));
    CascadeMux I__5648 (
            .O(N__26954),
            .I(N__26951));
    InMux I__5647 (
            .O(N__26951),
            .I(N__26947));
    InMux I__5646 (
            .O(N__26950),
            .I(N__26944));
    LocalMux I__5645 (
            .O(N__26947),
            .I(N__26941));
    LocalMux I__5644 (
            .O(N__26944),
            .I(N__26938));
    Span4Mux_h I__5643 (
            .O(N__26941),
            .I(N__26935));
    Span4Mux_h I__5642 (
            .O(N__26938),
            .I(N__26929));
    Span4Mux_h I__5641 (
            .O(N__26935),
            .I(N__26929));
    InMux I__5640 (
            .O(N__26934),
            .I(N__26926));
    Odrv4 I__5639 (
            .O(N__26929),
            .I(\b2v_inst.state_fastZ0Z_19 ));
    LocalMux I__5638 (
            .O(N__26926),
            .I(\b2v_inst.state_fastZ0Z_19 ));
    InMux I__5637 (
            .O(N__26921),
            .I(N__26918));
    LocalMux I__5636 (
            .O(N__26918),
            .I(\b2v_inst9.fsm_state_srsts_1_0 ));
    CascadeMux I__5635 (
            .O(N__26915),
            .I(N__26912));
    InMux I__5634 (
            .O(N__26912),
            .I(N__26909));
    LocalMux I__5633 (
            .O(N__26909),
            .I(\b2v_inst9.N_522 ));
    CascadeMux I__5632 (
            .O(N__26906),
            .I(\b2v_inst9.N_522_cascade_ ));
    InMux I__5631 (
            .O(N__26903),
            .I(N__26894));
    InMux I__5630 (
            .O(N__26902),
            .I(N__26891));
    InMux I__5629 (
            .O(N__26901),
            .I(N__26886));
    InMux I__5628 (
            .O(N__26900),
            .I(N__26886));
    InMux I__5627 (
            .O(N__26899),
            .I(N__26878));
    InMux I__5626 (
            .O(N__26898),
            .I(N__26875));
    InMux I__5625 (
            .O(N__26897),
            .I(N__26871));
    LocalMux I__5624 (
            .O(N__26894),
            .I(N__26866));
    LocalMux I__5623 (
            .O(N__26891),
            .I(N__26866));
    LocalMux I__5622 (
            .O(N__26886),
            .I(N__26863));
    InMux I__5621 (
            .O(N__26885),
            .I(N__26856));
    InMux I__5620 (
            .O(N__26884),
            .I(N__26856));
    InMux I__5619 (
            .O(N__26883),
            .I(N__26856));
    InMux I__5618 (
            .O(N__26882),
            .I(N__26851));
    InMux I__5617 (
            .O(N__26881),
            .I(N__26851));
    LocalMux I__5616 (
            .O(N__26878),
            .I(N__26848));
    LocalMux I__5615 (
            .O(N__26875),
            .I(N__26845));
    InMux I__5614 (
            .O(N__26874),
            .I(N__26842));
    LocalMux I__5613 (
            .O(N__26871),
            .I(N__26837));
    Span4Mux_v I__5612 (
            .O(N__26866),
            .I(N__26837));
    Span4Mux_v I__5611 (
            .O(N__26863),
            .I(N__26828));
    LocalMux I__5610 (
            .O(N__26856),
            .I(N__26828));
    LocalMux I__5609 (
            .O(N__26851),
            .I(N__26828));
    Span4Mux_h I__5608 (
            .O(N__26848),
            .I(N__26828));
    Odrv4 I__5607 (
            .O(N__26845),
            .I(\b2v_inst9.fsm_stateZ0Z_0 ));
    LocalMux I__5606 (
            .O(N__26842),
            .I(\b2v_inst9.fsm_stateZ0Z_0 ));
    Odrv4 I__5605 (
            .O(N__26837),
            .I(\b2v_inst9.fsm_stateZ0Z_0 ));
    Odrv4 I__5604 (
            .O(N__26828),
            .I(\b2v_inst9.fsm_stateZ0Z_0 ));
    InMux I__5603 (
            .O(N__26819),
            .I(N__26816));
    LocalMux I__5602 (
            .O(N__26816),
            .I(\b2v_inst.N_268 ));
    InMux I__5601 (
            .O(N__26813),
            .I(N__26810));
    LocalMux I__5600 (
            .O(N__26810),
            .I(\b2v_inst.un1_reg_anterior_iv_0_1_10 ));
    InMux I__5599 (
            .O(N__26807),
            .I(N__26804));
    LocalMux I__5598 (
            .O(N__26804),
            .I(N__26801));
    Span4Mux_h I__5597 (
            .O(N__26801),
            .I(N__26797));
    CascadeMux I__5596 (
            .O(N__26800),
            .I(N__26793));
    Span4Mux_h I__5595 (
            .O(N__26797),
            .I(N__26790));
    InMux I__5594 (
            .O(N__26796),
            .I(N__26785));
    InMux I__5593 (
            .O(N__26793),
            .I(N__26785));
    Odrv4 I__5592 (
            .O(N__26790),
            .I(SYNTHESIZED_WIRE_10_3));
    LocalMux I__5591 (
            .O(N__26785),
            .I(SYNTHESIZED_WIRE_10_3));
    InMux I__5590 (
            .O(N__26780),
            .I(N__26777));
    LocalMux I__5589 (
            .O(N__26777),
            .I(N__26774));
    Span12Mux_h I__5588 (
            .O(N__26774),
            .I(N__26770));
    InMux I__5587 (
            .O(N__26773),
            .I(N__26767));
    Odrv12 I__5586 (
            .O(N__26770),
            .I(SYNTHESIZED_WIRE_10_4));
    LocalMux I__5585 (
            .O(N__26767),
            .I(SYNTHESIZED_WIRE_10_4));
    InMux I__5584 (
            .O(N__26762),
            .I(N__26758));
    CascadeMux I__5583 (
            .O(N__26761),
            .I(N__26755));
    LocalMux I__5582 (
            .O(N__26758),
            .I(N__26752));
    InMux I__5581 (
            .O(N__26755),
            .I(N__26749));
    Odrv12 I__5580 (
            .O(N__26752),
            .I(SYNTHESIZED_WIRE_10_6));
    LocalMux I__5579 (
            .O(N__26749),
            .I(SYNTHESIZED_WIRE_10_6));
    InMux I__5578 (
            .O(N__26744),
            .I(N__26741));
    LocalMux I__5577 (
            .O(N__26741),
            .I(N__26738));
    Span4Mux_h I__5576 (
            .O(N__26738),
            .I(N__26734));
    CascadeMux I__5575 (
            .O(N__26737),
            .I(N__26731));
    Span4Mux_h I__5574 (
            .O(N__26734),
            .I(N__26728));
    InMux I__5573 (
            .O(N__26731),
            .I(N__26725));
    Odrv4 I__5572 (
            .O(N__26728),
            .I(SYNTHESIZED_WIRE_10_7));
    LocalMux I__5571 (
            .O(N__26725),
            .I(SYNTHESIZED_WIRE_10_7));
    InMux I__5570 (
            .O(N__26720),
            .I(N__26717));
    LocalMux I__5569 (
            .O(N__26717),
            .I(N__26713));
    CascadeMux I__5568 (
            .O(N__26716),
            .I(N__26709));
    Sp12to4 I__5567 (
            .O(N__26713),
            .I(N__26706));
    InMux I__5566 (
            .O(N__26712),
            .I(N__26703));
    InMux I__5565 (
            .O(N__26709),
            .I(N__26700));
    Span12Mux_v I__5564 (
            .O(N__26706),
            .I(N__26697));
    LocalMux I__5563 (
            .O(N__26703),
            .I(SYNTHESIZED_WIRE_10_0));
    LocalMux I__5562 (
            .O(N__26700),
            .I(SYNTHESIZED_WIRE_10_0));
    Odrv12 I__5561 (
            .O(N__26697),
            .I(SYNTHESIZED_WIRE_10_0));
    InMux I__5560 (
            .O(N__26690),
            .I(N__26686));
    InMux I__5559 (
            .O(N__26689),
            .I(N__26683));
    LocalMux I__5558 (
            .O(N__26686),
            .I(SYNTHESIZED_WIRE_5_0));
    LocalMux I__5557 (
            .O(N__26683),
            .I(SYNTHESIZED_WIRE_5_0));
    InMux I__5556 (
            .O(N__26678),
            .I(N__26675));
    LocalMux I__5555 (
            .O(N__26675),
            .I(N__26671));
    InMux I__5554 (
            .O(N__26674),
            .I(N__26668));
    Span4Mux_h I__5553 (
            .O(N__26671),
            .I(N__26665));
    LocalMux I__5552 (
            .O(N__26668),
            .I(\b2v_inst.eventosZ0Z_6 ));
    Odrv4 I__5551 (
            .O(N__26665),
            .I(\b2v_inst.eventosZ0Z_6 ));
    CascadeMux I__5550 (
            .O(N__26660),
            .I(\b2v_inst.un1_reg_anterior_iv_0_0_6_cascade_ ));
    InMux I__5549 (
            .O(N__26657),
            .I(N__26654));
    LocalMux I__5548 (
            .O(N__26654),
            .I(\b2v_inst.N_272 ));
    CEMux I__5547 (
            .O(N__26651),
            .I(N__26648));
    LocalMux I__5546 (
            .O(N__26648),
            .I(N__26644));
    CEMux I__5545 (
            .O(N__26647),
            .I(N__26641));
    Span4Mux_h I__5544 (
            .O(N__26644),
            .I(N__26638));
    LocalMux I__5543 (
            .O(N__26641),
            .I(N__26635));
    Odrv4 I__5542 (
            .O(N__26638),
            .I(\b2v_inst.data_a_escribir_1_sqmuxa ));
    Odrv12 I__5541 (
            .O(N__26635),
            .I(\b2v_inst.data_a_escribir_1_sqmuxa ));
    InMux I__5540 (
            .O(N__26630),
            .I(N__26627));
    LocalMux I__5539 (
            .O(N__26627),
            .I(N__26624));
    Span4Mux_h I__5538 (
            .O(N__26624),
            .I(N__26621));
    Odrv4 I__5537 (
            .O(N__26621),
            .I(\b2v_inst.data_a_escribir11_1_and ));
    InMux I__5536 (
            .O(N__26618),
            .I(N__26614));
    InMux I__5535 (
            .O(N__26617),
            .I(N__26611));
    LocalMux I__5534 (
            .O(N__26614),
            .I(N__26608));
    LocalMux I__5533 (
            .O(N__26611),
            .I(\b2v_inst.eventosZ0Z_4 ));
    Odrv4 I__5532 (
            .O(N__26608),
            .I(\b2v_inst.eventosZ0Z_4 ));
    CascadeMux I__5531 (
            .O(N__26603),
            .I(\b2v_inst.un1_reg_anterior_iv_0_0_4_cascade_ ));
    CascadeMux I__5530 (
            .O(N__26600),
            .I(\b2v_inst.un1_reg_anterior_iv_0_1_4_cascade_ ));
    InMux I__5529 (
            .O(N__26597),
            .I(N__26594));
    LocalMux I__5528 (
            .O(N__26594),
            .I(\b2v_inst.N_274 ));
    InMux I__5527 (
            .O(N__26591),
            .I(N__26587));
    InMux I__5526 (
            .O(N__26590),
            .I(N__26584));
    LocalMux I__5525 (
            .O(N__26587),
            .I(\b2v_inst.eventosZ0Z_0 ));
    LocalMux I__5524 (
            .O(N__26584),
            .I(\b2v_inst.eventosZ0Z_0 ));
    CascadeMux I__5523 (
            .O(N__26579),
            .I(\b2v_inst.data_a_escribir_RNO_2Z0Z_0_cascade_ ));
    CascadeMux I__5522 (
            .O(N__26576),
            .I(\b2v_inst.un1_reg_anterior_0_i_1_0_cascade_ ));
    InMux I__5521 (
            .O(N__26573),
            .I(N__26570));
    LocalMux I__5520 (
            .O(N__26570),
            .I(N__26566));
    InMux I__5519 (
            .O(N__26569),
            .I(N__26563));
    Odrv4 I__5518 (
            .O(N__26566),
            .I(\b2v_inst.eventosZ0Z_1 ));
    LocalMux I__5517 (
            .O(N__26563),
            .I(\b2v_inst.eventosZ0Z_1 ));
    CascadeMux I__5516 (
            .O(N__26558),
            .I(\b2v_inst.data_a_escribir_RNO_2Z0Z_1_cascade_ ));
    CascadeMux I__5515 (
            .O(N__26555),
            .I(\b2v_inst.un1_reg_anterior_0_i_1_1_cascade_ ));
    InMux I__5514 (
            .O(N__26552),
            .I(N__26548));
    InMux I__5513 (
            .O(N__26551),
            .I(N__26545));
    LocalMux I__5512 (
            .O(N__26548),
            .I(\b2v_inst.eventosZ0Z_10 ));
    LocalMux I__5511 (
            .O(N__26545),
            .I(\b2v_inst.eventosZ0Z_10 ));
    InMux I__5510 (
            .O(N__26540),
            .I(N__26537));
    LocalMux I__5509 (
            .O(N__26537),
            .I(\b2v_inst.N_269 ));
    CascadeMux I__5508 (
            .O(N__26534),
            .I(\b2v_inst.un1_reg_anterior_iv_0_0_10_cascade_ ));
    InMux I__5507 (
            .O(N__26531),
            .I(\b2v_inst.un2_valor_max1 ));
    InMux I__5506 (
            .O(N__26528),
            .I(N__26503));
    InMux I__5505 (
            .O(N__26527),
            .I(N__26503));
    InMux I__5504 (
            .O(N__26526),
            .I(N__26503));
    InMux I__5503 (
            .O(N__26525),
            .I(N__26503));
    InMux I__5502 (
            .O(N__26524),
            .I(N__26503));
    InMux I__5501 (
            .O(N__26523),
            .I(N__26503));
    InMux I__5500 (
            .O(N__26522),
            .I(N__26503));
    InMux I__5499 (
            .O(N__26521),
            .I(N__26500));
    InMux I__5498 (
            .O(N__26520),
            .I(N__26493));
    InMux I__5497 (
            .O(N__26519),
            .I(N__26493));
    InMux I__5496 (
            .O(N__26518),
            .I(N__26493));
    LocalMux I__5495 (
            .O(N__26503),
            .I(N__26490));
    LocalMux I__5494 (
            .O(N__26500),
            .I(N__26485));
    LocalMux I__5493 (
            .O(N__26493),
            .I(N__26485));
    Span4Mux_v I__5492 (
            .O(N__26490),
            .I(N__26482));
    Span4Mux_h I__5491 (
            .O(N__26485),
            .I(N__26479));
    Sp12to4 I__5490 (
            .O(N__26482),
            .I(N__26476));
    Span4Mux_h I__5489 (
            .O(N__26479),
            .I(N__26473));
    Span12Mux_h I__5488 (
            .O(N__26476),
            .I(N__26470));
    Span4Mux_h I__5487 (
            .O(N__26473),
            .I(N__26467));
    Odrv12 I__5486 (
            .O(N__26470),
            .I(\b2v_inst.ignorar_anchoZ0Z_1 ));
    Odrv4 I__5485 (
            .O(N__26467),
            .I(\b2v_inst.ignorar_anchoZ0Z_1 ));
    CEMux I__5484 (
            .O(N__26462),
            .I(N__26459));
    LocalMux I__5483 (
            .O(N__26459),
            .I(N__26455));
    CEMux I__5482 (
            .O(N__26458),
            .I(N__26452));
    Span4Mux_h I__5481 (
            .O(N__26455),
            .I(N__26446));
    LocalMux I__5480 (
            .O(N__26452),
            .I(N__26443));
    InMux I__5479 (
            .O(N__26451),
            .I(N__26436));
    InMux I__5478 (
            .O(N__26450),
            .I(N__26436));
    InMux I__5477 (
            .O(N__26449),
            .I(N__26433));
    Span4Mux_v I__5476 (
            .O(N__26446),
            .I(N__26430));
    Span4Mux_h I__5475 (
            .O(N__26443),
            .I(N__26427));
    InMux I__5474 (
            .O(N__26442),
            .I(N__26422));
    InMux I__5473 (
            .O(N__26441),
            .I(N__26422));
    LocalMux I__5472 (
            .O(N__26436),
            .I(N__26417));
    LocalMux I__5471 (
            .O(N__26433),
            .I(N__26417));
    Odrv4 I__5470 (
            .O(N__26430),
            .I(\b2v_inst.stateZ0Z_25 ));
    Odrv4 I__5469 (
            .O(N__26427),
            .I(\b2v_inst.stateZ0Z_25 ));
    LocalMux I__5468 (
            .O(N__26422),
            .I(\b2v_inst.stateZ0Z_25 ));
    Odrv4 I__5467 (
            .O(N__26417),
            .I(\b2v_inst.stateZ0Z_25 ));
    InMux I__5466 (
            .O(N__26408),
            .I(N__26405));
    LocalMux I__5465 (
            .O(N__26405),
            .I(N__26402));
    Odrv4 I__5464 (
            .O(N__26402),
            .I(\b2v_inst.data_a_escribir11_0_and ));
    CascadeMux I__5463 (
            .O(N__26399),
            .I(N__26396));
    InMux I__5462 (
            .O(N__26396),
            .I(N__26393));
    LocalMux I__5461 (
            .O(N__26393),
            .I(\b2v_inst.reg_ancho_1_i_3 ));
    CascadeMux I__5460 (
            .O(N__26390),
            .I(N__26387));
    InMux I__5459 (
            .O(N__26387),
            .I(N__26384));
    LocalMux I__5458 (
            .O(N__26384),
            .I(\b2v_inst.reg_ancho_1_i_4 ));
    CascadeMux I__5457 (
            .O(N__26381),
            .I(N__26378));
    InMux I__5456 (
            .O(N__26378),
            .I(N__26375));
    LocalMux I__5455 (
            .O(N__26375),
            .I(\b2v_inst.reg_ancho_1_i_5 ));
    CascadeMux I__5454 (
            .O(N__26372),
            .I(N__26369));
    InMux I__5453 (
            .O(N__26369),
            .I(N__26366));
    LocalMux I__5452 (
            .O(N__26366),
            .I(\b2v_inst.reg_ancho_1_i_6 ));
    CascadeMux I__5451 (
            .O(N__26363),
            .I(N__26360));
    InMux I__5450 (
            .O(N__26360),
            .I(N__26357));
    LocalMux I__5449 (
            .O(N__26357),
            .I(\b2v_inst.reg_ancho_1_i_7 ));
    CascadeMux I__5448 (
            .O(N__26354),
            .I(N__26351));
    InMux I__5447 (
            .O(N__26351),
            .I(N__26348));
    LocalMux I__5446 (
            .O(N__26348),
            .I(\b2v_inst.reg_ancho_1_i_8 ));
    CascadeMux I__5445 (
            .O(N__26345),
            .I(N__26342));
    InMux I__5444 (
            .O(N__26342),
            .I(N__26339));
    LocalMux I__5443 (
            .O(N__26339),
            .I(\b2v_inst.reg_ancho_1_i_9 ));
    CascadeMux I__5442 (
            .O(N__26336),
            .I(N__26333));
    InMux I__5441 (
            .O(N__26333),
            .I(N__26330));
    LocalMux I__5440 (
            .O(N__26330),
            .I(\b2v_inst.reg_ancho_1_i_10 ));
    CascadeMux I__5439 (
            .O(N__26327),
            .I(N__26324));
    InMux I__5438 (
            .O(N__26324),
            .I(N__26321));
    LocalMux I__5437 (
            .O(N__26321),
            .I(\b2v_inst.reg_ancho_1_i_0 ));
    CascadeMux I__5436 (
            .O(N__26318),
            .I(N__26315));
    InMux I__5435 (
            .O(N__26315),
            .I(N__26312));
    LocalMux I__5434 (
            .O(N__26312),
            .I(\b2v_inst.reg_ancho_1_i_1 ));
    CascadeMux I__5433 (
            .O(N__26309),
            .I(N__26306));
    InMux I__5432 (
            .O(N__26306),
            .I(N__26303));
    LocalMux I__5431 (
            .O(N__26303),
            .I(\b2v_inst.reg_ancho_1_i_2 ));
    InMux I__5430 (
            .O(N__26300),
            .I(N__26297));
    LocalMux I__5429 (
            .O(N__26297),
            .I(\b2v_inst.pix_data_regZ0Z_2 ));
    CascadeMux I__5428 (
            .O(N__26294),
            .I(N__26291));
    InMux I__5427 (
            .O(N__26291),
            .I(N__26288));
    LocalMux I__5426 (
            .O(N__26288),
            .I(\b2v_inst.pix_data_regZ0Z_5 ));
    InMux I__5425 (
            .O(N__26285),
            .I(N__26282));
    LocalMux I__5424 (
            .O(N__26282),
            .I(\b2v_inst.pix_data_regZ0Z_6 ));
    InMux I__5423 (
            .O(N__26279),
            .I(N__26276));
    LocalMux I__5422 (
            .O(N__26276),
            .I(\b2v_inst.pix_data_regZ0Z_7 ));
    InMux I__5421 (
            .O(N__26273),
            .I(N__26270));
    LocalMux I__5420 (
            .O(N__26270),
            .I(N__26267));
    Span4Mux_v I__5419 (
            .O(N__26267),
            .I(N__26264));
    Odrv4 I__5418 (
            .O(N__26264),
            .I(\b2v_inst9.N_583 ));
    IoInMux I__5417 (
            .O(N__26261),
            .I(N__26257));
    InMux I__5416 (
            .O(N__26260),
            .I(N__26254));
    LocalMux I__5415 (
            .O(N__26257),
            .I(N__26251));
    LocalMux I__5414 (
            .O(N__26254),
            .I(N__26248));
    IoSpan4Mux I__5413 (
            .O(N__26251),
            .I(N__26245));
    Span4Mux_h I__5412 (
            .O(N__26248),
            .I(N__26242));
    Span4Mux_s3_h I__5411 (
            .O(N__26245),
            .I(N__26239));
    Span4Mux_h I__5410 (
            .O(N__26242),
            .I(N__26236));
    Span4Mux_h I__5409 (
            .O(N__26239),
            .I(N__26233));
    Span4Mux_h I__5408 (
            .O(N__26236),
            .I(N__26230));
    Odrv4 I__5407 (
            .O(N__26233),
            .I(leds_c_9));
    Odrv4 I__5406 (
            .O(N__26230),
            .I(leds_c_9));
    InMux I__5405 (
            .O(N__26225),
            .I(N__26222));
    LocalMux I__5404 (
            .O(N__26222),
            .I(N__26218));
    InMux I__5403 (
            .O(N__26221),
            .I(N__26215));
    Span4Mux_h I__5402 (
            .O(N__26218),
            .I(N__26210));
    LocalMux I__5401 (
            .O(N__26215),
            .I(N__26210));
    Odrv4 I__5400 (
            .O(N__26210),
            .I(b2v_inst_energia_temp_9));
    CEMux I__5399 (
            .O(N__26207),
            .I(N__26202));
    CEMux I__5398 (
            .O(N__26206),
            .I(N__26199));
    CEMux I__5397 (
            .O(N__26205),
            .I(N__26194));
    LocalMux I__5396 (
            .O(N__26202),
            .I(N__26191));
    LocalMux I__5395 (
            .O(N__26199),
            .I(N__26187));
    CEMux I__5394 (
            .O(N__26198),
            .I(N__26184));
    CEMux I__5393 (
            .O(N__26197),
            .I(N__26181));
    LocalMux I__5392 (
            .O(N__26194),
            .I(N__26177));
    Span4Mux_v I__5391 (
            .O(N__26191),
            .I(N__26174));
    CEMux I__5390 (
            .O(N__26190),
            .I(N__26171));
    Span4Mux_v I__5389 (
            .O(N__26187),
            .I(N__26168));
    LocalMux I__5388 (
            .O(N__26184),
            .I(N__26163));
    LocalMux I__5387 (
            .O(N__26181),
            .I(N__26163));
    CEMux I__5386 (
            .O(N__26180),
            .I(N__26160));
    Span4Mux_v I__5385 (
            .O(N__26177),
            .I(N__26153));
    Span4Mux_h I__5384 (
            .O(N__26174),
            .I(N__26153));
    LocalMux I__5383 (
            .O(N__26171),
            .I(N__26153));
    Span4Mux_h I__5382 (
            .O(N__26168),
            .I(N__26150));
    Span4Mux_h I__5381 (
            .O(N__26163),
            .I(N__26145));
    LocalMux I__5380 (
            .O(N__26160),
            .I(N__26145));
    Span4Mux_v I__5379 (
            .O(N__26153),
            .I(N__26141));
    Span4Mux_v I__5378 (
            .O(N__26150),
            .I(N__26136));
    Span4Mux_v I__5377 (
            .O(N__26145),
            .I(N__26136));
    CEMux I__5376 (
            .O(N__26144),
            .I(N__26133));
    Span4Mux_v I__5375 (
            .O(N__26141),
            .I(N__26130));
    Span4Mux_v I__5374 (
            .O(N__26136),
            .I(N__26127));
    LocalMux I__5373 (
            .O(N__26133),
            .I(N__26124));
    Span4Mux_h I__5372 (
            .O(N__26130),
            .I(N__26121));
    Span4Mux_h I__5371 (
            .O(N__26127),
            .I(N__26116));
    Span4Mux_v I__5370 (
            .O(N__26124),
            .I(N__26116));
    Odrv4 I__5369 (
            .O(N__26121),
            .I(\b2v_inst.N_577_i ));
    Odrv4 I__5368 (
            .O(N__26116),
            .I(\b2v_inst.N_577_i ));
    InMux I__5367 (
            .O(N__26111),
            .I(N__26108));
    LocalMux I__5366 (
            .O(N__26108),
            .I(N__26105));
    Span4Mux_v I__5365 (
            .O(N__26105),
            .I(N__26102));
    Odrv4 I__5364 (
            .O(N__26102),
            .I(\b2v_inst9.data_to_sendZ0Z_0 ));
    IoInMux I__5363 (
            .O(N__26099),
            .I(N__26096));
    LocalMux I__5362 (
            .O(N__26096),
            .I(N__26093));
    IoSpan4Mux I__5361 (
            .O(N__26093),
            .I(N__26090));
    Span4Mux_s2_v I__5360 (
            .O(N__26090),
            .I(N__26087));
    Sp12to4 I__5359 (
            .O(N__26087),
            .I(N__26084));
    Span12Mux_s10_v I__5358 (
            .O(N__26084),
            .I(N__26081));
    Span12Mux_h I__5357 (
            .O(N__26081),
            .I(N__26078));
    Odrv12 I__5356 (
            .O(N__26078),
            .I(uart_tx_o_c));
    InMux I__5355 (
            .O(N__26075),
            .I(N__26071));
    InMux I__5354 (
            .O(N__26074),
            .I(N__26068));
    LocalMux I__5353 (
            .O(N__26071),
            .I(N__26062));
    LocalMux I__5352 (
            .O(N__26068),
            .I(N__26062));
    InMux I__5351 (
            .O(N__26067),
            .I(N__26057));
    Span4Mux_h I__5350 (
            .O(N__26062),
            .I(N__26054));
    InMux I__5349 (
            .O(N__26061),
            .I(N__26051));
    InMux I__5348 (
            .O(N__26060),
            .I(N__26048));
    LocalMux I__5347 (
            .O(N__26057),
            .I(N__26045));
    Span4Mux_h I__5346 (
            .O(N__26054),
            .I(N__26042));
    LocalMux I__5345 (
            .O(N__26051),
            .I(b2v_inst_state_2));
    LocalMux I__5344 (
            .O(N__26048),
            .I(b2v_inst_state_2));
    Odrv4 I__5343 (
            .O(N__26045),
            .I(b2v_inst_state_2));
    Odrv4 I__5342 (
            .O(N__26042),
            .I(b2v_inst_state_2));
    CascadeMux I__5341 (
            .O(N__26033),
            .I(N__26028));
    InMux I__5340 (
            .O(N__26032),
            .I(N__26025));
    CascadeMux I__5339 (
            .O(N__26031),
            .I(N__26022));
    InMux I__5338 (
            .O(N__26028),
            .I(N__26018));
    LocalMux I__5337 (
            .O(N__26025),
            .I(N__26015));
    InMux I__5336 (
            .O(N__26022),
            .I(N__26011));
    CascadeMux I__5335 (
            .O(N__26021),
            .I(N__26008));
    LocalMux I__5334 (
            .O(N__26018),
            .I(N__26005));
    Span4Mux_v I__5333 (
            .O(N__26015),
            .I(N__26001));
    InMux I__5332 (
            .O(N__26014),
            .I(N__25998));
    LocalMux I__5331 (
            .O(N__26011),
            .I(N__25995));
    InMux I__5330 (
            .O(N__26008),
            .I(N__25992));
    Span4Mux_v I__5329 (
            .O(N__26005),
            .I(N__25989));
    InMux I__5328 (
            .O(N__26004),
            .I(N__25986));
    Span4Mux_v I__5327 (
            .O(N__26001),
            .I(N__25981));
    LocalMux I__5326 (
            .O(N__25998),
            .I(N__25981));
    Span4Mux_v I__5325 (
            .O(N__25995),
            .I(N__25978));
    LocalMux I__5324 (
            .O(N__25992),
            .I(N__25975));
    Sp12to4 I__5323 (
            .O(N__25989),
            .I(N__25970));
    LocalMux I__5322 (
            .O(N__25986),
            .I(N__25970));
    Span4Mux_h I__5321 (
            .O(N__25981),
            .I(N__25963));
    Span4Mux_v I__5320 (
            .O(N__25978),
            .I(N__25963));
    Span4Mux_h I__5319 (
            .O(N__25975),
            .I(N__25963));
    Odrv12 I__5318 (
            .O(N__25970),
            .I(\b2v_inst.stateZ0Z_11 ));
    Odrv4 I__5317 (
            .O(N__25963),
            .I(\b2v_inst.stateZ0Z_11 ));
    InMux I__5316 (
            .O(N__25958),
            .I(N__25942));
    InMux I__5315 (
            .O(N__25957),
            .I(N__25942));
    InMux I__5314 (
            .O(N__25956),
            .I(N__25942));
    InMux I__5313 (
            .O(N__25955),
            .I(N__25942));
    InMux I__5312 (
            .O(N__25954),
            .I(N__25939));
    InMux I__5311 (
            .O(N__25953),
            .I(N__25936));
    InMux I__5310 (
            .O(N__25952),
            .I(N__25930));
    CascadeMux I__5309 (
            .O(N__25951),
            .I(N__25927));
    LocalMux I__5308 (
            .O(N__25942),
            .I(N__25922));
    LocalMux I__5307 (
            .O(N__25939),
            .I(N__25922));
    LocalMux I__5306 (
            .O(N__25936),
            .I(N__25919));
    CascadeMux I__5305 (
            .O(N__25935),
            .I(N__25916));
    CascadeMux I__5304 (
            .O(N__25934),
            .I(N__25913));
    CascadeMux I__5303 (
            .O(N__25933),
            .I(N__25906));
    LocalMux I__5302 (
            .O(N__25930),
            .I(N__25903));
    InMux I__5301 (
            .O(N__25927),
            .I(N__25900));
    Span4Mux_h I__5300 (
            .O(N__25922),
            .I(N__25896));
    Span4Mux_v I__5299 (
            .O(N__25919),
            .I(N__25893));
    InMux I__5298 (
            .O(N__25916),
            .I(N__25890));
    InMux I__5297 (
            .O(N__25913),
            .I(N__25887));
    InMux I__5296 (
            .O(N__25912),
            .I(N__25876));
    InMux I__5295 (
            .O(N__25911),
            .I(N__25876));
    InMux I__5294 (
            .O(N__25910),
            .I(N__25876));
    InMux I__5293 (
            .O(N__25909),
            .I(N__25876));
    InMux I__5292 (
            .O(N__25906),
            .I(N__25876));
    Span4Mux_h I__5291 (
            .O(N__25903),
            .I(N__25873));
    LocalMux I__5290 (
            .O(N__25900),
            .I(N__25870));
    CascadeMux I__5289 (
            .O(N__25899),
            .I(N__25867));
    Span4Mux_v I__5288 (
            .O(N__25896),
            .I(N__25864));
    Span4Mux_v I__5287 (
            .O(N__25893),
            .I(N__25861));
    LocalMux I__5286 (
            .O(N__25890),
            .I(N__25858));
    LocalMux I__5285 (
            .O(N__25887),
            .I(N__25853));
    LocalMux I__5284 (
            .O(N__25876),
            .I(N__25853));
    Span4Mux_v I__5283 (
            .O(N__25873),
            .I(N__25850));
    Span12Mux_v I__5282 (
            .O(N__25870),
            .I(N__25847));
    InMux I__5281 (
            .O(N__25867),
            .I(N__25844));
    Odrv4 I__5280 (
            .O(N__25864),
            .I(\b2v_inst.stateZ0Z_32 ));
    Odrv4 I__5279 (
            .O(N__25861),
            .I(\b2v_inst.stateZ0Z_32 ));
    Odrv4 I__5278 (
            .O(N__25858),
            .I(\b2v_inst.stateZ0Z_32 ));
    Odrv4 I__5277 (
            .O(N__25853),
            .I(\b2v_inst.stateZ0Z_32 ));
    Odrv4 I__5276 (
            .O(N__25850),
            .I(\b2v_inst.stateZ0Z_32 ));
    Odrv12 I__5275 (
            .O(N__25847),
            .I(\b2v_inst.stateZ0Z_32 ));
    LocalMux I__5274 (
            .O(N__25844),
            .I(\b2v_inst.stateZ0Z_32 ));
    InMux I__5273 (
            .O(N__25829),
            .I(N__25824));
    InMux I__5272 (
            .O(N__25828),
            .I(N__25821));
    InMux I__5271 (
            .O(N__25827),
            .I(N__25818));
    LocalMux I__5270 (
            .O(N__25824),
            .I(N__25807));
    LocalMux I__5269 (
            .O(N__25821),
            .I(N__25807));
    LocalMux I__5268 (
            .O(N__25818),
            .I(N__25807));
    InMux I__5267 (
            .O(N__25817),
            .I(N__25804));
    InMux I__5266 (
            .O(N__25816),
            .I(N__25799));
    InMux I__5265 (
            .O(N__25815),
            .I(N__25799));
    InMux I__5264 (
            .O(N__25814),
            .I(N__25796));
    Span4Mux_h I__5263 (
            .O(N__25807),
            .I(N__25793));
    LocalMux I__5262 (
            .O(N__25804),
            .I(b2v_inst_state_14));
    LocalMux I__5261 (
            .O(N__25799),
            .I(b2v_inst_state_14));
    LocalMux I__5260 (
            .O(N__25796),
            .I(b2v_inst_state_14));
    Odrv4 I__5259 (
            .O(N__25793),
            .I(b2v_inst_state_14));
    InMux I__5258 (
            .O(N__25784),
            .I(N__25781));
    LocalMux I__5257 (
            .O(N__25781),
            .I(\b2v_inst.state_ns_a3_i_0_a2_6_1 ));
    CascadeMux I__5256 (
            .O(N__25778),
            .I(\b2v_inst9.fsm_state_ns_i_0_i_0_1_cascade_ ));
    InMux I__5255 (
            .O(N__25775),
            .I(N__25771));
    InMux I__5254 (
            .O(N__25774),
            .I(N__25768));
    LocalMux I__5253 (
            .O(N__25771),
            .I(\b2v_inst9.N_832 ));
    LocalMux I__5252 (
            .O(N__25768),
            .I(\b2v_inst9.N_832 ));
    CascadeMux I__5251 (
            .O(N__25763),
            .I(N__25760));
    InMux I__5250 (
            .O(N__25760),
            .I(N__25757));
    LocalMux I__5249 (
            .O(N__25757),
            .I(N__25754));
    Span4Mux_h I__5248 (
            .O(N__25754),
            .I(N__25751));
    Odrv4 I__5247 (
            .O(N__25751),
            .I(\b2v_inst9.data_to_sendZ0Z_3 ));
    InMux I__5246 (
            .O(N__25748),
            .I(N__25745));
    LocalMux I__5245 (
            .O(N__25745),
            .I(\b2v_inst9.data_to_send_10_0_0_0_2 ));
    CascadeMux I__5244 (
            .O(N__25742),
            .I(N__25739));
    InMux I__5243 (
            .O(N__25739),
            .I(N__25735));
    InMux I__5242 (
            .O(N__25738),
            .I(N__25732));
    LocalMux I__5241 (
            .O(N__25735),
            .I(N__25728));
    LocalMux I__5240 (
            .O(N__25732),
            .I(N__25725));
    CascadeMux I__5239 (
            .O(N__25731),
            .I(N__25718));
    Span4Mux_h I__5238 (
            .O(N__25728),
            .I(N__25713));
    Span4Mux_h I__5237 (
            .O(N__25725),
            .I(N__25713));
    InMux I__5236 (
            .O(N__25724),
            .I(N__25708));
    InMux I__5235 (
            .O(N__25723),
            .I(N__25708));
    InMux I__5234 (
            .O(N__25722),
            .I(N__25701));
    InMux I__5233 (
            .O(N__25721),
            .I(N__25701));
    InMux I__5232 (
            .O(N__25718),
            .I(N__25701));
    Span4Mux_h I__5231 (
            .O(N__25713),
            .I(N__25698));
    LocalMux I__5230 (
            .O(N__25708),
            .I(b2v_inst_state_12));
    LocalMux I__5229 (
            .O(N__25701),
            .I(b2v_inst_state_12));
    Odrv4 I__5228 (
            .O(N__25698),
            .I(b2v_inst_state_12));
    InMux I__5227 (
            .O(N__25691),
            .I(N__25688));
    LocalMux I__5226 (
            .O(N__25688),
            .I(N__25682));
    InMux I__5225 (
            .O(N__25687),
            .I(N__25679));
    InMux I__5224 (
            .O(N__25686),
            .I(N__25676));
    InMux I__5223 (
            .O(N__25685),
            .I(N__25673));
    Span4Mux_v I__5222 (
            .O(N__25682),
            .I(N__25667));
    LocalMux I__5221 (
            .O(N__25679),
            .I(N__25667));
    LocalMux I__5220 (
            .O(N__25676),
            .I(N__25664));
    LocalMux I__5219 (
            .O(N__25673),
            .I(N__25661));
    CascadeMux I__5218 (
            .O(N__25672),
            .I(N__25658));
    Span4Mux_h I__5217 (
            .O(N__25667),
            .I(N__25655));
    Span4Mux_h I__5216 (
            .O(N__25664),
            .I(N__25650));
    Span4Mux_h I__5215 (
            .O(N__25661),
            .I(N__25650));
    InMux I__5214 (
            .O(N__25658),
            .I(N__25647));
    Odrv4 I__5213 (
            .O(N__25655),
            .I(b2v_inst_state_13));
    Odrv4 I__5212 (
            .O(N__25650),
            .I(b2v_inst_state_13));
    LocalMux I__5211 (
            .O(N__25647),
            .I(b2v_inst_state_13));
    InMux I__5210 (
            .O(N__25640),
            .I(N__25636));
    CascadeMux I__5209 (
            .O(N__25639),
            .I(N__25629));
    LocalMux I__5208 (
            .O(N__25636),
            .I(N__25625));
    InMux I__5207 (
            .O(N__25635),
            .I(N__25617));
    InMux I__5206 (
            .O(N__25634),
            .I(N__25617));
    InMux I__5205 (
            .O(N__25633),
            .I(N__25617));
    InMux I__5204 (
            .O(N__25632),
            .I(N__25614));
    InMux I__5203 (
            .O(N__25629),
            .I(N__25609));
    InMux I__5202 (
            .O(N__25628),
            .I(N__25609));
    Span4Mux_h I__5201 (
            .O(N__25625),
            .I(N__25606));
    InMux I__5200 (
            .O(N__25624),
            .I(N__25603));
    LocalMux I__5199 (
            .O(N__25617),
            .I(N__25598));
    LocalMux I__5198 (
            .O(N__25614),
            .I(N__25598));
    LocalMux I__5197 (
            .O(N__25609),
            .I(N__25595));
    Span4Mux_v I__5196 (
            .O(N__25606),
            .I(N__25590));
    LocalMux I__5195 (
            .O(N__25603),
            .I(N__25590));
    Span4Mux_h I__5194 (
            .O(N__25598),
            .I(N__25587));
    Span4Mux_h I__5193 (
            .O(N__25595),
            .I(N__25584));
    Odrv4 I__5192 (
            .O(N__25590),
            .I(\b2v_inst9.N_739 ));
    Odrv4 I__5191 (
            .O(N__25587),
            .I(\b2v_inst9.N_739 ));
    Odrv4 I__5190 (
            .O(N__25584),
            .I(\b2v_inst9.N_739 ));
    InMux I__5189 (
            .O(N__25577),
            .I(N__25574));
    LocalMux I__5188 (
            .O(N__25574),
            .I(\b2v_inst.pix_data_regZ0Z_0 ));
    InMux I__5187 (
            .O(N__25571),
            .I(N__25568));
    LocalMux I__5186 (
            .O(N__25568),
            .I(\b2v_inst.pix_data_regZ0Z_1 ));
    InMux I__5185 (
            .O(N__25565),
            .I(\b2v_inst.eventos_cry_6 ));
    InMux I__5184 (
            .O(N__25562),
            .I(bfn_15_11_0_));
    InMux I__5183 (
            .O(N__25559),
            .I(\b2v_inst.eventos_cry_8 ));
    InMux I__5182 (
            .O(N__25556),
            .I(\b2v_inst.eventos_cry_9 ));
    InMux I__5181 (
            .O(N__25553),
            .I(N__25550));
    LocalMux I__5180 (
            .O(N__25550),
            .I(N__25547));
    Span4Mux_h I__5179 (
            .O(N__25547),
            .I(N__25544));
    Odrv4 I__5178 (
            .O(N__25544),
            .I(\b2v_inst.state_ns_a3_i_0_a2_5_1 ));
    CascadeMux I__5177 (
            .O(N__25541),
            .I(\b2v_inst.state_ns_a3_i_0_a2_4_1_cascade_ ));
    InMux I__5176 (
            .O(N__25538),
            .I(N__25532));
    InMux I__5175 (
            .O(N__25537),
            .I(N__25532));
    LocalMux I__5174 (
            .O(N__25532),
            .I(N__25525));
    CascadeMux I__5173 (
            .O(N__25531),
            .I(N__25521));
    InMux I__5172 (
            .O(N__25530),
            .I(N__25516));
    InMux I__5171 (
            .O(N__25529),
            .I(N__25516));
    InMux I__5170 (
            .O(N__25528),
            .I(N__25513));
    Span4Mux_v I__5169 (
            .O(N__25525),
            .I(N__25510));
    InMux I__5168 (
            .O(N__25524),
            .I(N__25505));
    InMux I__5167 (
            .O(N__25521),
            .I(N__25505));
    LocalMux I__5166 (
            .O(N__25516),
            .I(N__25502));
    LocalMux I__5165 (
            .O(N__25513),
            .I(N__25495));
    Span4Mux_h I__5164 (
            .O(N__25510),
            .I(N__25495));
    LocalMux I__5163 (
            .O(N__25505),
            .I(N__25495));
    Span4Mux_h I__5162 (
            .O(N__25502),
            .I(N__25492));
    Span4Mux_h I__5161 (
            .O(N__25495),
            .I(N__25489));
    Odrv4 I__5160 (
            .O(N__25492),
            .I(\b2v_inst.stateZ0Z_31 ));
    Odrv4 I__5159 (
            .O(N__25489),
            .I(\b2v_inst.stateZ0Z_31 ));
    InMux I__5158 (
            .O(N__25484),
            .I(N__25480));
    CascadeMux I__5157 (
            .O(N__25483),
            .I(N__25477));
    LocalMux I__5156 (
            .O(N__25480),
            .I(N__25474));
    InMux I__5155 (
            .O(N__25477),
            .I(N__25471));
    Span4Mux_h I__5154 (
            .O(N__25474),
            .I(N__25464));
    LocalMux I__5153 (
            .O(N__25471),
            .I(N__25464));
    InMux I__5152 (
            .O(N__25470),
            .I(N__25459));
    InMux I__5151 (
            .O(N__25469),
            .I(N__25459));
    Span4Mux_h I__5150 (
            .O(N__25464),
            .I(N__25454));
    LocalMux I__5149 (
            .O(N__25459),
            .I(N__25451));
    InMux I__5148 (
            .O(N__25458),
            .I(N__25446));
    InMux I__5147 (
            .O(N__25457),
            .I(N__25446));
    Odrv4 I__5146 (
            .O(N__25454),
            .I(b2v_inst_state_7));
    Odrv12 I__5145 (
            .O(N__25451),
            .I(b2v_inst_state_7));
    LocalMux I__5144 (
            .O(N__25446),
            .I(b2v_inst_state_7));
    InMux I__5143 (
            .O(N__25439),
            .I(N__25434));
    InMux I__5142 (
            .O(N__25438),
            .I(N__25431));
    InMux I__5141 (
            .O(N__25437),
            .I(N__25428));
    LocalMux I__5140 (
            .O(N__25434),
            .I(N__25423));
    LocalMux I__5139 (
            .O(N__25431),
            .I(N__25423));
    LocalMux I__5138 (
            .O(N__25428),
            .I(N__25420));
    Span4Mux_h I__5137 (
            .O(N__25423),
            .I(N__25413));
    Span4Mux_v I__5136 (
            .O(N__25420),
            .I(N__25410));
    InMux I__5135 (
            .O(N__25419),
            .I(N__25407));
    InMux I__5134 (
            .O(N__25418),
            .I(N__25400));
    InMux I__5133 (
            .O(N__25417),
            .I(N__25400));
    InMux I__5132 (
            .O(N__25416),
            .I(N__25400));
    Span4Mux_h I__5131 (
            .O(N__25413),
            .I(N__25397));
    Odrv4 I__5130 (
            .O(N__25410),
            .I(b2v_inst_state_1));
    LocalMux I__5129 (
            .O(N__25407),
            .I(b2v_inst_state_1));
    LocalMux I__5128 (
            .O(N__25400),
            .I(b2v_inst_state_1));
    Odrv4 I__5127 (
            .O(N__25397),
            .I(b2v_inst_state_1));
    InMux I__5126 (
            .O(N__25388),
            .I(N__25385));
    LocalMux I__5125 (
            .O(N__25385),
            .I(\b2v_inst.data_a_escribir11_8_and ));
    InMux I__5124 (
            .O(N__25382),
            .I(N__25379));
    LocalMux I__5123 (
            .O(N__25379),
            .I(N__25376));
    Span4Mux_h I__5122 (
            .O(N__25376),
            .I(N__25373));
    Span4Mux_h I__5121 (
            .O(N__25373),
            .I(N__25370));
    Odrv4 I__5120 (
            .O(N__25370),
            .I(\b2v_inst.dir_mem_1Z0Z_10 ));
    InMux I__5119 (
            .O(N__25367),
            .I(N__25360));
    CascadeMux I__5118 (
            .O(N__25366),
            .I(N__25355));
    InMux I__5117 (
            .O(N__25365),
            .I(N__25350));
    InMux I__5116 (
            .O(N__25364),
            .I(N__25350));
    CascadeMux I__5115 (
            .O(N__25363),
            .I(N__25344));
    LocalMux I__5114 (
            .O(N__25360),
            .I(N__25341));
    InMux I__5113 (
            .O(N__25359),
            .I(N__25336));
    InMux I__5112 (
            .O(N__25358),
            .I(N__25333));
    InMux I__5111 (
            .O(N__25355),
            .I(N__25330));
    LocalMux I__5110 (
            .O(N__25350),
            .I(N__25327));
    InMux I__5109 (
            .O(N__25349),
            .I(N__25324));
    InMux I__5108 (
            .O(N__25348),
            .I(N__25321));
    InMux I__5107 (
            .O(N__25347),
            .I(N__25316));
    InMux I__5106 (
            .O(N__25344),
            .I(N__25316));
    Span4Mux_h I__5105 (
            .O(N__25341),
            .I(N__25313));
    InMux I__5104 (
            .O(N__25340),
            .I(N__25308));
    InMux I__5103 (
            .O(N__25339),
            .I(N__25308));
    LocalMux I__5102 (
            .O(N__25336),
            .I(N__25301));
    LocalMux I__5101 (
            .O(N__25333),
            .I(N__25301));
    LocalMux I__5100 (
            .O(N__25330),
            .I(N__25301));
    Odrv4 I__5099 (
            .O(N__25327),
            .I(\b2v_inst.N_490 ));
    LocalMux I__5098 (
            .O(N__25324),
            .I(\b2v_inst.N_490 ));
    LocalMux I__5097 (
            .O(N__25321),
            .I(\b2v_inst.N_490 ));
    LocalMux I__5096 (
            .O(N__25316),
            .I(\b2v_inst.N_490 ));
    Odrv4 I__5095 (
            .O(N__25313),
            .I(\b2v_inst.N_490 ));
    LocalMux I__5094 (
            .O(N__25308),
            .I(\b2v_inst.N_490 ));
    Odrv4 I__5093 (
            .O(N__25301),
            .I(\b2v_inst.N_490 ));
    CascadeMux I__5092 (
            .O(N__25286),
            .I(N__25283));
    InMux I__5091 (
            .O(N__25283),
            .I(N__25280));
    LocalMux I__5090 (
            .O(N__25280),
            .I(N__25277));
    Span4Mux_v I__5089 (
            .O(N__25277),
            .I(N__25274));
    Span4Mux_h I__5088 (
            .O(N__25274),
            .I(N__25271));
    Odrv4 I__5087 (
            .O(N__25271),
            .I(\b2v_inst.dir_mem_3Z0Z_10 ));
    InMux I__5086 (
            .O(N__25268),
            .I(N__25264));
    InMux I__5085 (
            .O(N__25267),
            .I(N__25261));
    LocalMux I__5084 (
            .O(N__25264),
            .I(N__25250));
    LocalMux I__5083 (
            .O(N__25261),
            .I(N__25245));
    InMux I__5082 (
            .O(N__25260),
            .I(N__25242));
    InMux I__5081 (
            .O(N__25259),
            .I(N__25237));
    InMux I__5080 (
            .O(N__25258),
            .I(N__25237));
    InMux I__5079 (
            .O(N__25257),
            .I(N__25234));
    InMux I__5078 (
            .O(N__25256),
            .I(N__25231));
    InMux I__5077 (
            .O(N__25255),
            .I(N__25228));
    InMux I__5076 (
            .O(N__25254),
            .I(N__25225));
    InMux I__5075 (
            .O(N__25253),
            .I(N__25222));
    Span4Mux_h I__5074 (
            .O(N__25250),
            .I(N__25219));
    InMux I__5073 (
            .O(N__25249),
            .I(N__25214));
    InMux I__5072 (
            .O(N__25248),
            .I(N__25214));
    Span4Mux_h I__5071 (
            .O(N__25245),
            .I(N__25207));
    LocalMux I__5070 (
            .O(N__25242),
            .I(N__25207));
    LocalMux I__5069 (
            .O(N__25237),
            .I(N__25207));
    LocalMux I__5068 (
            .O(N__25234),
            .I(N__25202));
    LocalMux I__5067 (
            .O(N__25231),
            .I(N__25202));
    LocalMux I__5066 (
            .O(N__25228),
            .I(\b2v_inst.N_488 ));
    LocalMux I__5065 (
            .O(N__25225),
            .I(\b2v_inst.N_488 ));
    LocalMux I__5064 (
            .O(N__25222),
            .I(\b2v_inst.N_488 ));
    Odrv4 I__5063 (
            .O(N__25219),
            .I(\b2v_inst.N_488 ));
    LocalMux I__5062 (
            .O(N__25214),
            .I(\b2v_inst.N_488 ));
    Odrv4 I__5061 (
            .O(N__25207),
            .I(\b2v_inst.N_488 ));
    Odrv4 I__5060 (
            .O(N__25202),
            .I(\b2v_inst.N_488 ));
    InMux I__5059 (
            .O(N__25187),
            .I(bfn_15_10_0_));
    InMux I__5058 (
            .O(N__25184),
            .I(\b2v_inst.eventos_cry_0 ));
    InMux I__5057 (
            .O(N__25181),
            .I(\b2v_inst.eventos_cry_1 ));
    InMux I__5056 (
            .O(N__25178),
            .I(\b2v_inst.eventos_cry_2 ));
    InMux I__5055 (
            .O(N__25175),
            .I(\b2v_inst.eventos_cry_3 ));
    InMux I__5054 (
            .O(N__25172),
            .I(\b2v_inst.eventos_cry_4 ));
    InMux I__5053 (
            .O(N__25169),
            .I(\b2v_inst.eventos_cry_5 ));
    InMux I__5052 (
            .O(N__25166),
            .I(N__25163));
    LocalMux I__5051 (
            .O(N__25163),
            .I(\b2v_inst.data_a_escribir11_4_and ));
    InMux I__5050 (
            .O(N__25160),
            .I(\b2v_inst.data_a_escribir12 ));
    InMux I__5049 (
            .O(N__25157),
            .I(N__25154));
    LocalMux I__5048 (
            .O(N__25154),
            .I(\b2v_inst.data_a_escribir11_9_and ));
    InMux I__5047 (
            .O(N__25151),
            .I(N__25148));
    LocalMux I__5046 (
            .O(N__25148),
            .I(\b2v_inst.data_a_escribir11_2_and ));
    CascadeMux I__5045 (
            .O(N__25145),
            .I(N__25142));
    InMux I__5044 (
            .O(N__25142),
            .I(N__25138));
    InMux I__5043 (
            .O(N__25141),
            .I(N__25135));
    LocalMux I__5042 (
            .O(N__25138),
            .I(N__25132));
    LocalMux I__5041 (
            .O(N__25135),
            .I(N__25129));
    Span4Mux_v I__5040 (
            .O(N__25132),
            .I(N__25126));
    Span4Mux_h I__5039 (
            .O(N__25129),
            .I(N__25123));
    Span4Mux_h I__5038 (
            .O(N__25126),
            .I(N__25120));
    Span4Mux_h I__5037 (
            .O(N__25123),
            .I(N__25117));
    Odrv4 I__5036 (
            .O(N__25120),
            .I(b2v_inst_energia_temp_10));
    Odrv4 I__5035 (
            .O(N__25117),
            .I(b2v_inst_energia_temp_10));
    InMux I__5034 (
            .O(N__25112),
            .I(\b2v_inst.un14_data_ram_energia_o_cry_9 ));
    InMux I__5033 (
            .O(N__25109),
            .I(N__25106));
    LocalMux I__5032 (
            .O(N__25106),
            .I(N__25102));
    InMux I__5031 (
            .O(N__25105),
            .I(N__25099));
    Span4Mux_v I__5030 (
            .O(N__25102),
            .I(N__25096));
    LocalMux I__5029 (
            .O(N__25099),
            .I(N__25093));
    Span4Mux_v I__5028 (
            .O(N__25096),
            .I(N__25088));
    Span4Mux_h I__5027 (
            .O(N__25093),
            .I(N__25088));
    Span4Mux_h I__5026 (
            .O(N__25088),
            .I(N__25085));
    Odrv4 I__5025 (
            .O(N__25085),
            .I(b2v_inst_energia_temp_11));
    InMux I__5024 (
            .O(N__25082),
            .I(N__25079));
    LocalMux I__5023 (
            .O(N__25079),
            .I(N__25076));
    Span4Mux_v I__5022 (
            .O(N__25076),
            .I(N__25073));
    Span4Mux_h I__5021 (
            .O(N__25073),
            .I(N__25070));
    Span4Mux_h I__5020 (
            .O(N__25070),
            .I(N__25067));
    Odrv4 I__5019 (
            .O(N__25067),
            .I(SYNTHESIZED_WIRE_13_11));
    InMux I__5018 (
            .O(N__25064),
            .I(\b2v_inst.un14_data_ram_energia_o_cry_10 ));
    InMux I__5017 (
            .O(N__25061),
            .I(N__25058));
    LocalMux I__5016 (
            .O(N__25058),
            .I(N__25054));
    InMux I__5015 (
            .O(N__25057),
            .I(N__25051));
    Span4Mux_h I__5014 (
            .O(N__25054),
            .I(N__25048));
    LocalMux I__5013 (
            .O(N__25051),
            .I(N__25045));
    Span4Mux_v I__5012 (
            .O(N__25048),
            .I(N__25042));
    Span4Mux_h I__5011 (
            .O(N__25045),
            .I(N__25039));
    Odrv4 I__5010 (
            .O(N__25042),
            .I(b2v_inst_energia_temp_12));
    Odrv4 I__5009 (
            .O(N__25039),
            .I(b2v_inst_energia_temp_12));
    InMux I__5008 (
            .O(N__25034),
            .I(N__25031));
    LocalMux I__5007 (
            .O(N__25031),
            .I(N__25028));
    Span4Mux_v I__5006 (
            .O(N__25028),
            .I(N__25025));
    Span4Mux_v I__5005 (
            .O(N__25025),
            .I(N__25022));
    Sp12to4 I__5004 (
            .O(N__25022),
            .I(N__25019));
    Odrv12 I__5003 (
            .O(N__25019),
            .I(SYNTHESIZED_WIRE_13_12));
    InMux I__5002 (
            .O(N__25016),
            .I(\b2v_inst.un14_data_ram_energia_o_cry_11 ));
    InMux I__5001 (
            .O(N__25013),
            .I(N__25010));
    LocalMux I__5000 (
            .O(N__25010),
            .I(N__25006));
    InMux I__4999 (
            .O(N__25009),
            .I(N__25003));
    Span4Mux_h I__4998 (
            .O(N__25006),
            .I(N__25000));
    LocalMux I__4997 (
            .O(N__25003),
            .I(b2v_inst_energia_temp_13));
    Odrv4 I__4996 (
            .O(N__25000),
            .I(b2v_inst_energia_temp_13));
    InMux I__4995 (
            .O(N__24995),
            .I(\b2v_inst.un14_data_ram_energia_o_cry_12 ));
    InMux I__4994 (
            .O(N__24992),
            .I(N__24989));
    LocalMux I__4993 (
            .O(N__24989),
            .I(N__24986));
    Span4Mux_v I__4992 (
            .O(N__24986),
            .I(N__24983));
    Sp12to4 I__4991 (
            .O(N__24983),
            .I(N__24980));
    Odrv12 I__4990 (
            .O(N__24980),
            .I(SYNTHESIZED_WIRE_13_13));
    IoInMux I__4989 (
            .O(N__24977),
            .I(N__24973));
    InMux I__4988 (
            .O(N__24976),
            .I(N__24970));
    LocalMux I__4987 (
            .O(N__24973),
            .I(N__24967));
    LocalMux I__4986 (
            .O(N__24970),
            .I(N__24964));
    Span4Mux_s3_h I__4985 (
            .O(N__24967),
            .I(N__24961));
    Span4Mux_v I__4984 (
            .O(N__24964),
            .I(N__24958));
    Span4Mux_h I__4983 (
            .O(N__24961),
            .I(N__24955));
    Sp12to4 I__4982 (
            .O(N__24958),
            .I(N__24952));
    Odrv4 I__4981 (
            .O(N__24955),
            .I(leds_c_8));
    Odrv12 I__4980 (
            .O(N__24952),
            .I(leds_c_8));
    InMux I__4979 (
            .O(N__24947),
            .I(N__24944));
    LocalMux I__4978 (
            .O(N__24944),
            .I(N__24940));
    InMux I__4977 (
            .O(N__24943),
            .I(N__24937));
    Odrv4 I__4976 (
            .O(N__24940),
            .I(b2v_inst_energia_temp_8));
    LocalMux I__4975 (
            .O(N__24937),
            .I(b2v_inst_energia_temp_8));
    InMux I__4974 (
            .O(N__24932),
            .I(N__24929));
    LocalMux I__4973 (
            .O(N__24929),
            .I(\b2v_inst.un14_data_ram_energia_o_cry_9_c_RNI28GBZ0 ));
    InMux I__4972 (
            .O(N__24926),
            .I(N__24923));
    LocalMux I__4971 (
            .O(N__24923),
            .I(N__24920));
    Span4Mux_h I__4970 (
            .O(N__24920),
            .I(N__24917));
    Span4Mux_h I__4969 (
            .O(N__24917),
            .I(N__24914));
    Span4Mux_h I__4968 (
            .O(N__24914),
            .I(N__24911));
    Odrv4 I__4967 (
            .O(N__24911),
            .I(N_461_i));
    CascadeMux I__4966 (
            .O(N__24908),
            .I(N__24904));
    InMux I__4965 (
            .O(N__24907),
            .I(N__24901));
    InMux I__4964 (
            .O(N__24904),
            .I(N__24898));
    LocalMux I__4963 (
            .O(N__24901),
            .I(b2v_inst_energia_temp_2));
    LocalMux I__4962 (
            .O(N__24898),
            .I(b2v_inst_energia_temp_2));
    InMux I__4961 (
            .O(N__24893),
            .I(N__24890));
    LocalMux I__4960 (
            .O(N__24890),
            .I(N__24887));
    Odrv4 I__4959 (
            .O(N__24887),
            .I(\b2v_inst.un14_data_ram_energia_o_cry_1_c_RNIHM5MZ0 ));
    InMux I__4958 (
            .O(N__24884),
            .I(\b2v_inst.un14_data_ram_energia_o_cry_1 ));
    CascadeMux I__4957 (
            .O(N__24881),
            .I(N__24877));
    InMux I__4956 (
            .O(N__24880),
            .I(N__24874));
    InMux I__4955 (
            .O(N__24877),
            .I(N__24871));
    LocalMux I__4954 (
            .O(N__24874),
            .I(b2v_inst_energia_temp_3));
    LocalMux I__4953 (
            .O(N__24871),
            .I(b2v_inst_energia_temp_3));
    InMux I__4952 (
            .O(N__24866),
            .I(N__24863));
    LocalMux I__4951 (
            .O(N__24863),
            .I(N__24860));
    Odrv4 I__4950 (
            .O(N__24860),
            .I(\b2v_inst.un14_data_ram_energia_o_cry_2_c_RNIKQ6MZ0 ));
    InMux I__4949 (
            .O(N__24857),
            .I(\b2v_inst.un14_data_ram_energia_o_cry_2 ));
    InMux I__4948 (
            .O(N__24854),
            .I(N__24851));
    LocalMux I__4947 (
            .O(N__24851),
            .I(N__24848));
    Span4Mux_v I__4946 (
            .O(N__24848),
            .I(N__24845));
    Span4Mux_h I__4945 (
            .O(N__24845),
            .I(N__24842));
    Span4Mux_h I__4944 (
            .O(N__24842),
            .I(N__24839));
    Odrv4 I__4943 (
            .O(N__24839),
            .I(\b2v_inst.pix_data_regZ0Z_4 ));
    CascadeMux I__4942 (
            .O(N__24836),
            .I(N__24832));
    InMux I__4941 (
            .O(N__24835),
            .I(N__24829));
    InMux I__4940 (
            .O(N__24832),
            .I(N__24826));
    LocalMux I__4939 (
            .O(N__24829),
            .I(N__24823));
    LocalMux I__4938 (
            .O(N__24826),
            .I(N__24820));
    Span4Mux_v I__4937 (
            .O(N__24823),
            .I(N__24815));
    Span4Mux_v I__4936 (
            .O(N__24820),
            .I(N__24815));
    Span4Mux_h I__4935 (
            .O(N__24815),
            .I(N__24812));
    Span4Mux_v I__4934 (
            .O(N__24812),
            .I(N__24809));
    Odrv4 I__4933 (
            .O(N__24809),
            .I(b2v_inst_energia_temp_4));
    InMux I__4932 (
            .O(N__24806),
            .I(N__24803));
    LocalMux I__4931 (
            .O(N__24803),
            .I(N__24800));
    Span4Mux_h I__4930 (
            .O(N__24800),
            .I(N__24797));
    Odrv4 I__4929 (
            .O(N__24797),
            .I(\b2v_inst.un14_data_ram_energia_o_cry_3_c_RNINU7MZ0 ));
    InMux I__4928 (
            .O(N__24794),
            .I(\b2v_inst.un14_data_ram_energia_o_cry_3 ));
    InMux I__4927 (
            .O(N__24791),
            .I(N__24787));
    InMux I__4926 (
            .O(N__24790),
            .I(N__24784));
    LocalMux I__4925 (
            .O(N__24787),
            .I(N__24779));
    LocalMux I__4924 (
            .O(N__24784),
            .I(N__24779));
    Span12Mux_v I__4923 (
            .O(N__24779),
            .I(N__24776));
    Odrv12 I__4922 (
            .O(N__24776),
            .I(b2v_inst_energia_temp_5));
    InMux I__4921 (
            .O(N__24773),
            .I(N__24770));
    LocalMux I__4920 (
            .O(N__24770),
            .I(\b2v_inst.un14_data_ram_energia_o_cry_4_c_RNIQ29MZ0 ));
    InMux I__4919 (
            .O(N__24767),
            .I(\b2v_inst.un14_data_ram_energia_o_cry_4 ));
    InMux I__4918 (
            .O(N__24764),
            .I(N__24760));
    CascadeMux I__4917 (
            .O(N__24763),
            .I(N__24757));
    LocalMux I__4916 (
            .O(N__24760),
            .I(N__24754));
    InMux I__4915 (
            .O(N__24757),
            .I(N__24751));
    Span4Mux_v I__4914 (
            .O(N__24754),
            .I(N__24746));
    LocalMux I__4913 (
            .O(N__24751),
            .I(N__24746));
    Span4Mux_h I__4912 (
            .O(N__24746),
            .I(N__24743));
    Odrv4 I__4911 (
            .O(N__24743),
            .I(b2v_inst_energia_temp_6));
    InMux I__4910 (
            .O(N__24740),
            .I(N__24737));
    LocalMux I__4909 (
            .O(N__24737),
            .I(N__24734));
    Odrv12 I__4908 (
            .O(N__24734),
            .I(\b2v_inst.un14_data_ram_energia_o_cry_5_c_RNIT6AMZ0 ));
    InMux I__4907 (
            .O(N__24731),
            .I(\b2v_inst.un14_data_ram_energia_o_cry_5 ));
    InMux I__4906 (
            .O(N__24728),
            .I(N__24724));
    CascadeMux I__4905 (
            .O(N__24727),
            .I(N__24721));
    LocalMux I__4904 (
            .O(N__24724),
            .I(N__24718));
    InMux I__4903 (
            .O(N__24721),
            .I(N__24715));
    Span4Mux_v I__4902 (
            .O(N__24718),
            .I(N__24710));
    LocalMux I__4901 (
            .O(N__24715),
            .I(N__24710));
    Span4Mux_v I__4900 (
            .O(N__24710),
            .I(N__24707));
    Span4Mux_h I__4899 (
            .O(N__24707),
            .I(N__24704));
    Odrv4 I__4898 (
            .O(N__24704),
            .I(b2v_inst_energia_temp_7));
    InMux I__4897 (
            .O(N__24701),
            .I(N__24698));
    LocalMux I__4896 (
            .O(N__24698),
            .I(\b2v_inst.un14_data_ram_energia_o_cry_6_c_RNI0BBMZ0 ));
    InMux I__4895 (
            .O(N__24695),
            .I(\b2v_inst.un14_data_ram_energia_o_cry_6 ));
    InMux I__4894 (
            .O(N__24692),
            .I(N__24689));
    LocalMux I__4893 (
            .O(N__24689),
            .I(N__24686));
    Span4Mux_h I__4892 (
            .O(N__24686),
            .I(N__24683));
    Odrv4 I__4891 (
            .O(N__24683),
            .I(\b2v_inst.un14_data_ram_energia_o_cry_7_c_RNIN84CZ0 ));
    InMux I__4890 (
            .O(N__24680),
            .I(bfn_14_15_0_));
    InMux I__4889 (
            .O(N__24677),
            .I(N__24674));
    LocalMux I__4888 (
            .O(N__24674),
            .I(N__24671));
    Span4Mux_h I__4887 (
            .O(N__24671),
            .I(N__24668));
    Odrv4 I__4886 (
            .O(N__24668),
            .I(\b2v_inst.un14_data_ram_energia_o_cry_8_c_RNIPB5CZ0 ));
    InMux I__4885 (
            .O(N__24665),
            .I(\b2v_inst.un14_data_ram_energia_o_cry_8 ));
    InMux I__4884 (
            .O(N__24662),
            .I(N__24653));
    InMux I__4883 (
            .O(N__24661),
            .I(N__24653));
    InMux I__4882 (
            .O(N__24660),
            .I(N__24650));
    InMux I__4881 (
            .O(N__24659),
            .I(N__24647));
    InMux I__4880 (
            .O(N__24658),
            .I(N__24644));
    LocalMux I__4879 (
            .O(N__24653),
            .I(N__24639));
    LocalMux I__4878 (
            .O(N__24650),
            .I(N__24639));
    LocalMux I__4877 (
            .O(N__24647),
            .I(N__24634));
    LocalMux I__4876 (
            .O(N__24644),
            .I(N__24634));
    Span4Mux_h I__4875 (
            .O(N__24639),
            .I(N__24629));
    Span4Mux_h I__4874 (
            .O(N__24634),
            .I(N__24629));
    Odrv4 I__4873 (
            .O(N__24629),
            .I(b2v_inst_state_15));
    CascadeMux I__4872 (
            .O(N__24626),
            .I(\b2v_inst9.N_832_cascade_ ));
    InMux I__4871 (
            .O(N__24623),
            .I(N__24620));
    LocalMux I__4870 (
            .O(N__24620),
            .I(N__24617));
    Odrv12 I__4869 (
            .O(N__24617),
            .I(\b2v_inst9.data_to_send_10_0_0_0_1 ));
    InMux I__4868 (
            .O(N__24614),
            .I(N__24611));
    LocalMux I__4867 (
            .O(N__24611),
            .I(N__24608));
    Odrv12 I__4866 (
            .O(N__24608),
            .I(\b2v_inst9.data_to_send_10_0_0_1_1 ));
    CascadeMux I__4865 (
            .O(N__24605),
            .I(\b2v_inst9.data_to_send_10_0_0_2_2_cascade_ ));
    InMux I__4864 (
            .O(N__24602),
            .I(N__24599));
    LocalMux I__4863 (
            .O(N__24599),
            .I(N__24596));
    Odrv4 I__4862 (
            .O(N__24596),
            .I(\b2v_inst9.data_to_sendZ0Z_2 ));
    CEMux I__4861 (
            .O(N__24593),
            .I(N__24587));
    CEMux I__4860 (
            .O(N__24592),
            .I(N__24584));
    CEMux I__4859 (
            .O(N__24591),
            .I(N__24581));
    CEMux I__4858 (
            .O(N__24590),
            .I(N__24578));
    LocalMux I__4857 (
            .O(N__24587),
            .I(N__24575));
    LocalMux I__4856 (
            .O(N__24584),
            .I(N__24570));
    LocalMux I__4855 (
            .O(N__24581),
            .I(N__24570));
    LocalMux I__4854 (
            .O(N__24578),
            .I(N__24567));
    Odrv4 I__4853 (
            .O(N__24575),
            .I(\b2v_inst9.un2_n_fsm_state_0_sqmuxa_2_0_i_0 ));
    Odrv4 I__4852 (
            .O(N__24570),
            .I(\b2v_inst9.un2_n_fsm_state_0_sqmuxa_2_0_i_0 ));
    Odrv4 I__4851 (
            .O(N__24567),
            .I(\b2v_inst9.un2_n_fsm_state_0_sqmuxa_2_0_i_0 ));
    InMux I__4850 (
            .O(N__24560),
            .I(N__24551));
    InMux I__4849 (
            .O(N__24559),
            .I(N__24551));
    InMux I__4848 (
            .O(N__24558),
            .I(N__24551));
    LocalMux I__4847 (
            .O(N__24551),
            .I(N__24545));
    InMux I__4846 (
            .O(N__24550),
            .I(N__24540));
    InMux I__4845 (
            .O(N__24549),
            .I(N__24540));
    InMux I__4844 (
            .O(N__24548),
            .I(N__24537));
    Odrv12 I__4843 (
            .O(N__24545),
            .I(\b2v_inst9.N_740 ));
    LocalMux I__4842 (
            .O(N__24540),
            .I(\b2v_inst9.N_740 ));
    LocalMux I__4841 (
            .O(N__24537),
            .I(\b2v_inst9.N_740 ));
    InMux I__4840 (
            .O(N__24530),
            .I(N__24527));
    LocalMux I__4839 (
            .O(N__24527),
            .I(\b2v_inst9.data_to_send_10_0_0_1_2 ));
    InMux I__4838 (
            .O(N__24524),
            .I(N__24516));
    InMux I__4837 (
            .O(N__24523),
            .I(N__24516));
    InMux I__4836 (
            .O(N__24522),
            .I(N__24508));
    InMux I__4835 (
            .O(N__24521),
            .I(N__24508));
    LocalMux I__4834 (
            .O(N__24516),
            .I(N__24505));
    InMux I__4833 (
            .O(N__24515),
            .I(N__24500));
    InMux I__4832 (
            .O(N__24514),
            .I(N__24500));
    InMux I__4831 (
            .O(N__24513),
            .I(N__24497));
    LocalMux I__4830 (
            .O(N__24508),
            .I(\b2v_inst9.N_738 ));
    Odrv4 I__4829 (
            .O(N__24505),
            .I(\b2v_inst9.N_738 ));
    LocalMux I__4828 (
            .O(N__24500),
            .I(\b2v_inst9.N_738 ));
    LocalMux I__4827 (
            .O(N__24497),
            .I(\b2v_inst9.N_738 ));
    CascadeMux I__4826 (
            .O(N__24488),
            .I(N__24484));
    InMux I__4825 (
            .O(N__24487),
            .I(N__24481));
    InMux I__4824 (
            .O(N__24484),
            .I(N__24478));
    LocalMux I__4823 (
            .O(N__24481),
            .I(N__24470));
    LocalMux I__4822 (
            .O(N__24478),
            .I(N__24470));
    CascadeMux I__4821 (
            .O(N__24477),
            .I(N__24467));
    CascadeMux I__4820 (
            .O(N__24476),
            .I(N__24463));
    CascadeMux I__4819 (
            .O(N__24475),
            .I(N__24460));
    Span4Mux_h I__4818 (
            .O(N__24470),
            .I(N__24457));
    InMux I__4817 (
            .O(N__24467),
            .I(N__24452));
    InMux I__4816 (
            .O(N__24466),
            .I(N__24452));
    InMux I__4815 (
            .O(N__24463),
            .I(N__24449));
    InMux I__4814 (
            .O(N__24460),
            .I(N__24446));
    Odrv4 I__4813 (
            .O(N__24457),
            .I(\b2v_inst9.N_741 ));
    LocalMux I__4812 (
            .O(N__24452),
            .I(\b2v_inst9.N_741 ));
    LocalMux I__4811 (
            .O(N__24449),
            .I(\b2v_inst9.N_741 ));
    LocalMux I__4810 (
            .O(N__24446),
            .I(\b2v_inst9.N_741 ));
    InMux I__4809 (
            .O(N__24437),
            .I(N__24434));
    LocalMux I__4808 (
            .O(N__24434),
            .I(N__24431));
    Span4Mux_h I__4807 (
            .O(N__24431),
            .I(N__24428));
    Odrv4 I__4806 (
            .O(N__24428),
            .I(\b2v_inst9.data_to_send_10_0_0_1_3 ));
    InMux I__4805 (
            .O(N__24425),
            .I(N__24422));
    LocalMux I__4804 (
            .O(N__24422),
            .I(N__24418));
    CascadeMux I__4803 (
            .O(N__24421),
            .I(N__24415));
    Span4Mux_h I__4802 (
            .O(N__24418),
            .I(N__24412));
    InMux I__4801 (
            .O(N__24415),
            .I(N__24409));
    Odrv4 I__4800 (
            .O(N__24412),
            .I(b2v_inst_energia_temp_0));
    LocalMux I__4799 (
            .O(N__24409),
            .I(b2v_inst_energia_temp_0));
    InMux I__4798 (
            .O(N__24404),
            .I(N__24401));
    LocalMux I__4797 (
            .O(N__24401),
            .I(N__24398));
    Span4Mux_h I__4796 (
            .O(N__24398),
            .I(N__24395));
    Span4Mux_v I__4795 (
            .O(N__24395),
            .I(N__24392));
    Odrv4 I__4794 (
            .O(N__24392),
            .I(\b2v_inst.un14_data_ram_energia_o_axb_0 ));
    InMux I__4793 (
            .O(N__24389),
            .I(N__24385));
    CascadeMux I__4792 (
            .O(N__24388),
            .I(N__24382));
    LocalMux I__4791 (
            .O(N__24385),
            .I(N__24379));
    InMux I__4790 (
            .O(N__24382),
            .I(N__24376));
    Odrv4 I__4789 (
            .O(N__24379),
            .I(b2v_inst_energia_temp_1));
    LocalMux I__4788 (
            .O(N__24376),
            .I(b2v_inst_energia_temp_1));
    InMux I__4787 (
            .O(N__24371),
            .I(N__24368));
    LocalMux I__4786 (
            .O(N__24368),
            .I(N__24365));
    Span4Mux_v I__4785 (
            .O(N__24365),
            .I(N__24362));
    Span4Mux_v I__4784 (
            .O(N__24362),
            .I(N__24359));
    Odrv4 I__4783 (
            .O(N__24359),
            .I(\b2v_inst.un14_data_ram_energia_o_cry_0_c_RNIEI4MZ0 ));
    InMux I__4782 (
            .O(N__24356),
            .I(\b2v_inst.un14_data_ram_energia_o_cry_0 ));
    InMux I__4781 (
            .O(N__24353),
            .I(N__24350));
    LocalMux I__4780 (
            .O(N__24350),
            .I(\b2v_inst9.data_to_send_10_0_0_0_6 ));
    CascadeMux I__4779 (
            .O(N__24347),
            .I(\b2v_inst9.data_to_send_10_0_0_0_7_cascade_ ));
    CascadeMux I__4778 (
            .O(N__24344),
            .I(N__24340));
    InMux I__4777 (
            .O(N__24343),
            .I(N__24335));
    InMux I__4776 (
            .O(N__24340),
            .I(N__24335));
    LocalMux I__4775 (
            .O(N__24335),
            .I(\b2v_inst9.data_to_sendZ0Z_7 ));
    InMux I__4774 (
            .O(N__24332),
            .I(N__24329));
    LocalMux I__4773 (
            .O(N__24329),
            .I(\b2v_inst9.data_to_send_10_0_0_2_0 ));
    InMux I__4772 (
            .O(N__24326),
            .I(N__24323));
    LocalMux I__4771 (
            .O(N__24323),
            .I(N__24320));
    Span4Mux_v I__4770 (
            .O(N__24320),
            .I(N__24317));
    Odrv4 I__4769 (
            .O(N__24317),
            .I(\b2v_inst9.data_to_send_10_0_0_1_0 ));
    CascadeMux I__4768 (
            .O(N__24314),
            .I(\b2v_inst9.N_738_cascade_ ));
    InMux I__4767 (
            .O(N__24311),
            .I(N__24308));
    LocalMux I__4766 (
            .O(N__24308),
            .I(N__24305));
    Odrv4 I__4765 (
            .O(N__24305),
            .I(\b2v_inst9.data_to_send_10_0_0_2_1 ));
    InMux I__4764 (
            .O(N__24302),
            .I(N__24299));
    LocalMux I__4763 (
            .O(N__24299),
            .I(N__24296));
    Span4Mux_v I__4762 (
            .O(N__24296),
            .I(N__24293));
    Odrv4 I__4761 (
            .O(N__24293),
            .I(\b2v_inst9.data_to_sendZ0Z_1 ));
    CascadeMux I__4760 (
            .O(N__24290),
            .I(N_478_cascade_));
    InMux I__4759 (
            .O(N__24287),
            .I(N__24284));
    LocalMux I__4758 (
            .O(N__24284),
            .I(\b2v_inst9.data_to_send_10_0_0_0_0 ));
    InMux I__4757 (
            .O(N__24281),
            .I(N__24277));
    InMux I__4756 (
            .O(N__24280),
            .I(N__24270));
    LocalMux I__4755 (
            .O(N__24277),
            .I(N__24267));
    InMux I__4754 (
            .O(N__24276),
            .I(N__24258));
    InMux I__4753 (
            .O(N__24275),
            .I(N__24258));
    InMux I__4752 (
            .O(N__24274),
            .I(N__24258));
    InMux I__4751 (
            .O(N__24273),
            .I(N__24258));
    LocalMux I__4750 (
            .O(N__24270),
            .I(N__24251));
    Span4Mux_h I__4749 (
            .O(N__24267),
            .I(N__24246));
    LocalMux I__4748 (
            .O(N__24258),
            .I(N__24246));
    InMux I__4747 (
            .O(N__24257),
            .I(N__24237));
    InMux I__4746 (
            .O(N__24256),
            .I(N__24237));
    InMux I__4745 (
            .O(N__24255),
            .I(N__24237));
    InMux I__4744 (
            .O(N__24254),
            .I(N__24237));
    Odrv4 I__4743 (
            .O(N__24251),
            .I(\b2v_inst.N_655 ));
    Odrv4 I__4742 (
            .O(N__24246),
            .I(\b2v_inst.N_655 ));
    LocalMux I__4741 (
            .O(N__24237),
            .I(\b2v_inst.N_655 ));
    InMux I__4740 (
            .O(N__24230),
            .I(N__24227));
    LocalMux I__4739 (
            .O(N__24227),
            .I(N__24223));
    CascadeMux I__4738 (
            .O(N__24226),
            .I(N__24220));
    Span4Mux_h I__4737 (
            .O(N__24223),
            .I(N__24217));
    InMux I__4736 (
            .O(N__24220),
            .I(N__24214));
    Odrv4 I__4735 (
            .O(N__24217),
            .I(\b2v_inst.un4_cuenta_cry_4_c_RNIFZ0Z888 ));
    LocalMux I__4734 (
            .O(N__24214),
            .I(\b2v_inst.un4_cuenta_cry_4_c_RNIFZ0Z888 ));
    CascadeMux I__4733 (
            .O(N__24209),
            .I(N__24206));
    InMux I__4732 (
            .O(N__24206),
            .I(N__24202));
    InMux I__4731 (
            .O(N__24205),
            .I(N__24199));
    LocalMux I__4730 (
            .O(N__24202),
            .I(N__24196));
    LocalMux I__4729 (
            .O(N__24199),
            .I(N__24193));
    Span4Mux_h I__4728 (
            .O(N__24196),
            .I(N__24188));
    Span4Mux_v I__4727 (
            .O(N__24193),
            .I(N__24188));
    Odrv4 I__4726 (
            .O(N__24188),
            .I(\b2v_inst.cuentaZ0Z_5 ));
    CEMux I__4725 (
            .O(N__24185),
            .I(N__24182));
    LocalMux I__4724 (
            .O(N__24182),
            .I(N__24176));
    CEMux I__4723 (
            .O(N__24181),
            .I(N__24173));
    CEMux I__4722 (
            .O(N__24180),
            .I(N__24170));
    CEMux I__4721 (
            .O(N__24179),
            .I(N__24167));
    Span4Mux_v I__4720 (
            .O(N__24176),
            .I(N__24162));
    LocalMux I__4719 (
            .O(N__24173),
            .I(N__24162));
    LocalMux I__4718 (
            .O(N__24170),
            .I(N__24159));
    LocalMux I__4717 (
            .O(N__24167),
            .I(N__24156));
    Span4Mux_v I__4716 (
            .O(N__24162),
            .I(N__24153));
    Span4Mux_v I__4715 (
            .O(N__24159),
            .I(N__24150));
    Span4Mux_h I__4714 (
            .O(N__24156),
            .I(N__24147));
    Span4Mux_h I__4713 (
            .O(N__24153),
            .I(N__24144));
    Odrv4 I__4712 (
            .O(N__24150),
            .I(\b2v_inst.N_547_i_0 ));
    Odrv4 I__4711 (
            .O(N__24147),
            .I(\b2v_inst.N_547_i_0 ));
    Odrv4 I__4710 (
            .O(N__24144),
            .I(\b2v_inst.N_547_i_0 ));
    InMux I__4709 (
            .O(N__24137),
            .I(N__24134));
    LocalMux I__4708 (
            .O(N__24134),
            .I(N__24131));
    Odrv4 I__4707 (
            .O(N__24131),
            .I(\b2v_inst9.data_to_send_10_0_0_0_4 ));
    CascadeMux I__4706 (
            .O(N__24128),
            .I(N__24125));
    InMux I__4705 (
            .O(N__24125),
            .I(N__24122));
    LocalMux I__4704 (
            .O(N__24122),
            .I(\b2v_inst9.data_to_sendZ0Z_4 ));
    InMux I__4703 (
            .O(N__24119),
            .I(N__24116));
    LocalMux I__4702 (
            .O(N__24116),
            .I(\b2v_inst9.data_to_send_10_0_0_1_4 ));
    InMux I__4701 (
            .O(N__24113),
            .I(N__24110));
    LocalMux I__4700 (
            .O(N__24110),
            .I(N__24107));
    Odrv4 I__4699 (
            .O(N__24107),
            .I(\b2v_inst9.data_to_send_10_0_0_1_5 ));
    InMux I__4698 (
            .O(N__24104),
            .I(N__24101));
    LocalMux I__4697 (
            .O(N__24101),
            .I(N__24098));
    Span4Mux_h I__4696 (
            .O(N__24098),
            .I(N__24095));
    Odrv4 I__4695 (
            .O(N__24095),
            .I(\b2v_inst9.fsm_state_ns_i_i_0_a2_2_2Z0Z_0 ));
    CascadeMux I__4694 (
            .O(N__24092),
            .I(\b2v_inst9.N_583_cascade_ ));
    InMux I__4693 (
            .O(N__24089),
            .I(N__24085));
    IoInMux I__4692 (
            .O(N__24088),
            .I(N__24082));
    LocalMux I__4691 (
            .O(N__24085),
            .I(N__24079));
    LocalMux I__4690 (
            .O(N__24082),
            .I(N__24076));
    Span12Mux_v I__4689 (
            .O(N__24079),
            .I(N__24073));
    Span4Mux_s3_h I__4688 (
            .O(N__24076),
            .I(N__24070));
    Span12Mux_h I__4687 (
            .O(N__24073),
            .I(N__24067));
    Span4Mux_v I__4686 (
            .O(N__24070),
            .I(N__24064));
    Odrv12 I__4685 (
            .O(N__24067),
            .I(reset_c_i));
    Odrv4 I__4684 (
            .O(N__24064),
            .I(reset_c_i));
    CascadeMux I__4683 (
            .O(N__24059),
            .I(\b2v_inst9.un2_n_fsm_state_0_sqmuxa_2_0_i_cascade_ ));
    InMux I__4682 (
            .O(N__24056),
            .I(N__24053));
    LocalMux I__4681 (
            .O(N__24053),
            .I(N__24050));
    Span4Mux_h I__4680 (
            .O(N__24050),
            .I(N__24047));
    Odrv4 I__4679 (
            .O(N__24047),
            .I(\b2v_inst.dir_energia_s_6 ));
    InMux I__4678 (
            .O(N__24044),
            .I(\b2v_inst.dir_energia_cry_5 ));
    InMux I__4677 (
            .O(N__24041),
            .I(N__24038));
    LocalMux I__4676 (
            .O(N__24038),
            .I(N__24035));
    Span4Mux_h I__4675 (
            .O(N__24035),
            .I(N__24032));
    Odrv4 I__4674 (
            .O(N__24032),
            .I(\b2v_inst.dir_energia_s_7 ));
    InMux I__4673 (
            .O(N__24029),
            .I(\b2v_inst.dir_energia_cry_6 ));
    InMux I__4672 (
            .O(N__24026),
            .I(N__24023));
    LocalMux I__4671 (
            .O(N__24023),
            .I(N__24020));
    Span4Mux_h I__4670 (
            .O(N__24020),
            .I(N__24017));
    Odrv4 I__4669 (
            .O(N__24017),
            .I(\b2v_inst.dir_energia_s_8 ));
    InMux I__4668 (
            .O(N__24014),
            .I(bfn_13_17_0_));
    InMux I__4667 (
            .O(N__24011),
            .I(N__24008));
    LocalMux I__4666 (
            .O(N__24008),
            .I(N__24005));
    Span4Mux_h I__4665 (
            .O(N__24005),
            .I(N__24002));
    Odrv4 I__4664 (
            .O(N__24002),
            .I(\b2v_inst.dir_energia_s_9 ));
    InMux I__4663 (
            .O(N__23999),
            .I(\b2v_inst.dir_energia_cry_8 ));
    InMux I__4662 (
            .O(N__23996),
            .I(N__23993));
    LocalMux I__4661 (
            .O(N__23993),
            .I(N__23990));
    Span4Mux_v I__4660 (
            .O(N__23990),
            .I(N__23987));
    Span4Mux_h I__4659 (
            .O(N__23987),
            .I(N__23984));
    Odrv4 I__4658 (
            .O(N__23984),
            .I(\b2v_inst.dir_energia_s_10 ));
    InMux I__4657 (
            .O(N__23981),
            .I(\b2v_inst.dir_energia_cry_9 ));
    InMux I__4656 (
            .O(N__23978),
            .I(N__23973));
    CascadeMux I__4655 (
            .O(N__23977),
            .I(N__23970));
    CascadeMux I__4654 (
            .O(N__23976),
            .I(N__23963));
    LocalMux I__4653 (
            .O(N__23973),
            .I(N__23960));
    InMux I__4652 (
            .O(N__23970),
            .I(N__23951));
    InMux I__4651 (
            .O(N__23969),
            .I(N__23951));
    InMux I__4650 (
            .O(N__23968),
            .I(N__23951));
    InMux I__4649 (
            .O(N__23967),
            .I(N__23951));
    InMux I__4648 (
            .O(N__23966),
            .I(N__23945));
    InMux I__4647 (
            .O(N__23963),
            .I(N__23942));
    Span4Mux_v I__4646 (
            .O(N__23960),
            .I(N__23939));
    LocalMux I__4645 (
            .O(N__23951),
            .I(N__23936));
    InMux I__4644 (
            .O(N__23950),
            .I(N__23929));
    InMux I__4643 (
            .O(N__23949),
            .I(N__23929));
    InMux I__4642 (
            .O(N__23948),
            .I(N__23929));
    LocalMux I__4641 (
            .O(N__23945),
            .I(N__23926));
    LocalMux I__4640 (
            .O(N__23942),
            .I(N__23921));
    Span4Mux_h I__4639 (
            .O(N__23939),
            .I(N__23921));
    Span4Mux_v I__4638 (
            .O(N__23936),
            .I(N__23916));
    LocalMux I__4637 (
            .O(N__23929),
            .I(N__23916));
    Span4Mux_v I__4636 (
            .O(N__23926),
            .I(N__23909));
    Span4Mux_v I__4635 (
            .O(N__23921),
            .I(N__23904));
    Span4Mux_v I__4634 (
            .O(N__23916),
            .I(N__23904));
    InMux I__4633 (
            .O(N__23915),
            .I(N__23899));
    InMux I__4632 (
            .O(N__23914),
            .I(N__23899));
    InMux I__4631 (
            .O(N__23913),
            .I(N__23894));
    InMux I__4630 (
            .O(N__23912),
            .I(N__23894));
    Sp12to4 I__4629 (
            .O(N__23909),
            .I(N__23885));
    Sp12to4 I__4628 (
            .O(N__23904),
            .I(N__23885));
    LocalMux I__4627 (
            .O(N__23899),
            .I(N__23885));
    LocalMux I__4626 (
            .O(N__23894),
            .I(N__23885));
    Odrv12 I__4625 (
            .O(N__23885),
            .I(\b2v_inst.stateZ0Z_19 ));
    CascadeMux I__4624 (
            .O(N__23882),
            .I(N__23879));
    InMux I__4623 (
            .O(N__23879),
            .I(N__23876));
    LocalMux I__4622 (
            .O(N__23876),
            .I(N__23862));
    InMux I__4621 (
            .O(N__23875),
            .I(N__23847));
    InMux I__4620 (
            .O(N__23874),
            .I(N__23847));
    InMux I__4619 (
            .O(N__23873),
            .I(N__23847));
    InMux I__4618 (
            .O(N__23872),
            .I(N__23847));
    InMux I__4617 (
            .O(N__23871),
            .I(N__23847));
    InMux I__4616 (
            .O(N__23870),
            .I(N__23847));
    InMux I__4615 (
            .O(N__23869),
            .I(N__23847));
    InMux I__4614 (
            .O(N__23868),
            .I(N__23838));
    InMux I__4613 (
            .O(N__23867),
            .I(N__23838));
    InMux I__4612 (
            .O(N__23866),
            .I(N__23838));
    InMux I__4611 (
            .O(N__23865),
            .I(N__23838));
    Span4Mux_v I__4610 (
            .O(N__23862),
            .I(N__23835));
    LocalMux I__4609 (
            .O(N__23847),
            .I(\b2v_inst.N_352_0 ));
    LocalMux I__4608 (
            .O(N__23838),
            .I(\b2v_inst.N_352_0 ));
    Odrv4 I__4607 (
            .O(N__23835),
            .I(\b2v_inst.N_352_0 ));
    InMux I__4606 (
            .O(N__23828),
            .I(\b2v_inst.dir_energia_cry_10 ));
    CascadeMux I__4605 (
            .O(N__23825),
            .I(N__23822));
    InMux I__4604 (
            .O(N__23822),
            .I(N__23819));
    LocalMux I__4603 (
            .O(N__23819),
            .I(N__23815));
    InMux I__4602 (
            .O(N__23818),
            .I(N__23812));
    Span4Mux_h I__4601 (
            .O(N__23815),
            .I(N__23809));
    LocalMux I__4600 (
            .O(N__23812),
            .I(\b2v_inst.dir_energiaZ0Z_11 ));
    Odrv4 I__4599 (
            .O(N__23809),
            .I(\b2v_inst.dir_energiaZ0Z_11 ));
    CEMux I__4598 (
            .O(N__23804),
            .I(N__23801));
    LocalMux I__4597 (
            .O(N__23801),
            .I(N__23796));
    CEMux I__4596 (
            .O(N__23800),
            .I(N__23793));
    CEMux I__4595 (
            .O(N__23799),
            .I(N__23790));
    Span4Mux_v I__4594 (
            .O(N__23796),
            .I(N__23785));
    LocalMux I__4593 (
            .O(N__23793),
            .I(N__23785));
    LocalMux I__4592 (
            .O(N__23790),
            .I(N__23782));
    Span4Mux_h I__4591 (
            .O(N__23785),
            .I(N__23779));
    Odrv4 I__4590 (
            .O(N__23782),
            .I(\b2v_inst.N_430_i ));
    Odrv4 I__4589 (
            .O(N__23779),
            .I(\b2v_inst.N_430_i ));
    InMux I__4588 (
            .O(N__23774),
            .I(N__23771));
    LocalMux I__4587 (
            .O(N__23771),
            .I(N__23768));
    Odrv4 I__4586 (
            .O(N__23768),
            .I(\b2v_inst.N_648_5 ));
    InMux I__4585 (
            .O(N__23765),
            .I(N__23756));
    InMux I__4584 (
            .O(N__23764),
            .I(N__23756));
    InMux I__4583 (
            .O(N__23763),
            .I(N__23756));
    LocalMux I__4582 (
            .O(N__23756),
            .I(N__23753));
    Span4Mux_h I__4581 (
            .O(N__23753),
            .I(N__23750));
    Span4Mux_v I__4580 (
            .O(N__23750),
            .I(N__23745));
    InMux I__4579 (
            .O(N__23749),
            .I(N__23742));
    InMux I__4578 (
            .O(N__23748),
            .I(N__23739));
    Span4Mux_v I__4577 (
            .O(N__23745),
            .I(N__23736));
    LocalMux I__4576 (
            .O(N__23742),
            .I(N__23733));
    LocalMux I__4575 (
            .O(N__23739),
            .I(\b2v_inst.un9_indice_0_a2_5_1 ));
    Odrv4 I__4574 (
            .O(N__23736),
            .I(\b2v_inst.un9_indice_0_a2_5_1 ));
    Odrv4 I__4573 (
            .O(N__23733),
            .I(\b2v_inst.un9_indice_0_a2_5_1 ));
    InMux I__4572 (
            .O(N__23726),
            .I(N__23723));
    LocalMux I__4571 (
            .O(N__23723),
            .I(N__23720));
    Span4Mux_v I__4570 (
            .O(N__23720),
            .I(N__23715));
    InMux I__4569 (
            .O(N__23719),
            .I(N__23710));
    InMux I__4568 (
            .O(N__23718),
            .I(N__23710));
    Odrv4 I__4567 (
            .O(N__23715),
            .I(\b2v_inst.un4_cuenta_cry_9_c_RNI01TZ0Z9 ));
    LocalMux I__4566 (
            .O(N__23710),
            .I(\b2v_inst.un4_cuenta_cry_9_c_RNI01TZ0Z9 ));
    InMux I__4565 (
            .O(N__23705),
            .I(N__23701));
    CascadeMux I__4564 (
            .O(N__23704),
            .I(N__23698));
    LocalMux I__4563 (
            .O(N__23701),
            .I(N__23695));
    InMux I__4562 (
            .O(N__23698),
            .I(N__23692));
    Span4Mux_v I__4561 (
            .O(N__23695),
            .I(N__23687));
    LocalMux I__4560 (
            .O(N__23692),
            .I(N__23687));
    Span4Mux_v I__4559 (
            .O(N__23687),
            .I(N__23684));
    Odrv4 I__4558 (
            .O(N__23684),
            .I(\b2v_inst.cuentaZ0Z_10 ));
    InMux I__4557 (
            .O(N__23681),
            .I(N__23678));
    LocalMux I__4556 (
            .O(N__23678),
            .I(N__23675));
    Span4Mux_h I__4555 (
            .O(N__23675),
            .I(N__23671));
    IoInMux I__4554 (
            .O(N__23674),
            .I(N__23668));
    Span4Mux_v I__4553 (
            .O(N__23671),
            .I(N__23665));
    LocalMux I__4552 (
            .O(N__23668),
            .I(N__23662));
    Span4Mux_h I__4551 (
            .O(N__23665),
            .I(N__23659));
    Odrv12 I__4550 (
            .O(N__23662),
            .I(leds_c_2));
    Odrv4 I__4549 (
            .O(N__23659),
            .I(leds_c_2));
    InMux I__4548 (
            .O(N__23654),
            .I(N__23650));
    IoInMux I__4547 (
            .O(N__23653),
            .I(N__23647));
    LocalMux I__4546 (
            .O(N__23650),
            .I(N__23644));
    LocalMux I__4545 (
            .O(N__23647),
            .I(N__23641));
    Span4Mux_v I__4544 (
            .O(N__23644),
            .I(N__23638));
    Span4Mux_s3_h I__4543 (
            .O(N__23641),
            .I(N__23635));
    Span4Mux_h I__4542 (
            .O(N__23638),
            .I(N__23632));
    Span4Mux_h I__4541 (
            .O(N__23635),
            .I(N__23629));
    Span4Mux_h I__4540 (
            .O(N__23632),
            .I(N__23626));
    Odrv4 I__4539 (
            .O(N__23629),
            .I(leds_c_3));
    Odrv4 I__4538 (
            .O(N__23626),
            .I(leds_c_3));
    InMux I__4537 (
            .O(N__23621),
            .I(N__23618));
    LocalMux I__4536 (
            .O(N__23618),
            .I(N__23615));
    Span4Mux_h I__4535 (
            .O(N__23615),
            .I(N__23612));
    Span4Mux_h I__4534 (
            .O(N__23612),
            .I(N__23609));
    Span4Mux_h I__4533 (
            .O(N__23609),
            .I(N__23606));
    Odrv4 I__4532 (
            .O(N__23606),
            .I(N_546_i));
    InMux I__4531 (
            .O(N__23603),
            .I(N__23600));
    LocalMux I__4530 (
            .O(N__23600),
            .I(N__23597));
    Span4Mux_h I__4529 (
            .O(N__23597),
            .I(N__23594));
    Odrv4 I__4528 (
            .O(N__23594),
            .I(\b2v_inst.dir_energia_s_1 ));
    InMux I__4527 (
            .O(N__23591),
            .I(\b2v_inst.dir_energia_cry_0 ));
    CascadeMux I__4526 (
            .O(N__23588),
            .I(N__23585));
    InMux I__4525 (
            .O(N__23585),
            .I(N__23582));
    LocalMux I__4524 (
            .O(N__23582),
            .I(N__23579));
    Span4Mux_v I__4523 (
            .O(N__23579),
            .I(N__23576));
    Odrv4 I__4522 (
            .O(N__23576),
            .I(\b2v_inst.dir_energia_s_2 ));
    InMux I__4521 (
            .O(N__23573),
            .I(\b2v_inst.dir_energia_cry_1 ));
    InMux I__4520 (
            .O(N__23570),
            .I(N__23567));
    LocalMux I__4519 (
            .O(N__23567),
            .I(N__23564));
    Span4Mux_v I__4518 (
            .O(N__23564),
            .I(N__23561));
    Odrv4 I__4517 (
            .O(N__23561),
            .I(\b2v_inst.dir_energia_s_3 ));
    InMux I__4516 (
            .O(N__23558),
            .I(\b2v_inst.dir_energia_cry_2 ));
    CascadeMux I__4515 (
            .O(N__23555),
            .I(N__23552));
    InMux I__4514 (
            .O(N__23552),
            .I(N__23549));
    LocalMux I__4513 (
            .O(N__23549),
            .I(N__23546));
    Span4Mux_v I__4512 (
            .O(N__23546),
            .I(N__23543));
    Span4Mux_h I__4511 (
            .O(N__23543),
            .I(N__23540));
    Odrv4 I__4510 (
            .O(N__23540),
            .I(\b2v_inst.dir_energia_s_4 ));
    InMux I__4509 (
            .O(N__23537),
            .I(\b2v_inst.dir_energia_cry_3 ));
    InMux I__4508 (
            .O(N__23534),
            .I(N__23531));
    LocalMux I__4507 (
            .O(N__23531),
            .I(N__23528));
    Span4Mux_h I__4506 (
            .O(N__23528),
            .I(N__23525));
    Odrv4 I__4505 (
            .O(N__23525),
            .I(\b2v_inst.dir_energia_s_5 ));
    InMux I__4504 (
            .O(N__23522),
            .I(\b2v_inst.dir_energia_cry_4 ));
    InMux I__4503 (
            .O(N__23519),
            .I(N__23516));
    LocalMux I__4502 (
            .O(N__23516),
            .I(N__23513));
    Span4Mux_v I__4501 (
            .O(N__23513),
            .I(N__23509));
    InMux I__4500 (
            .O(N__23512),
            .I(N__23506));
    Odrv4 I__4499 (
            .O(N__23509),
            .I(\b2v_inst.cuentaZ0Z_9 ));
    LocalMux I__4498 (
            .O(N__23506),
            .I(\b2v_inst.cuentaZ0Z_9 ));
    InMux I__4497 (
            .O(N__23501),
            .I(N__23498));
    LocalMux I__4496 (
            .O(N__23498),
            .I(N__23493));
    InMux I__4495 (
            .O(N__23497),
            .I(N__23488));
    InMux I__4494 (
            .O(N__23496),
            .I(N__23488));
    Odrv12 I__4493 (
            .O(N__23493),
            .I(\b2v_inst.un4_cuenta_cry_8_c_RNINKCZ0Z8 ));
    LocalMux I__4492 (
            .O(N__23488),
            .I(\b2v_inst.un4_cuenta_cry_8_c_RNINKCZ0Z8 ));
    InMux I__4491 (
            .O(N__23483),
            .I(bfn_13_13_0_));
    InMux I__4490 (
            .O(N__23480),
            .I(\b2v_inst.un4_cuenta_cry_9 ));
    InMux I__4489 (
            .O(N__23477),
            .I(N__23474));
    LocalMux I__4488 (
            .O(N__23474),
            .I(N__23471));
    Span4Mux_h I__4487 (
            .O(N__23471),
            .I(N__23468));
    Span4Mux_h I__4486 (
            .O(N__23468),
            .I(N__23465));
    Odrv4 I__4485 (
            .O(N__23465),
            .I(N_458_i));
    InMux I__4484 (
            .O(N__23462),
            .I(N__23459));
    LocalMux I__4483 (
            .O(N__23459),
            .I(N__23455));
    CascadeMux I__4482 (
            .O(N__23458),
            .I(N__23452));
    Span4Mux_h I__4481 (
            .O(N__23455),
            .I(N__23447));
    InMux I__4480 (
            .O(N__23452),
            .I(N__23440));
    InMux I__4479 (
            .O(N__23451),
            .I(N__23440));
    InMux I__4478 (
            .O(N__23450),
            .I(N__23440));
    Odrv4 I__4477 (
            .O(N__23447),
            .I(b2v_inst_state_4));
    LocalMux I__4476 (
            .O(N__23440),
            .I(b2v_inst_state_4));
    InMux I__4475 (
            .O(N__23435),
            .I(N__23432));
    LocalMux I__4474 (
            .O(N__23432),
            .I(N__23427));
    CascadeMux I__4473 (
            .O(N__23431),
            .I(N__23424));
    CascadeMux I__4472 (
            .O(N__23430),
            .I(N__23420));
    Span4Mux_v I__4471 (
            .O(N__23427),
            .I(N__23417));
    InMux I__4470 (
            .O(N__23424),
            .I(N__23410));
    InMux I__4469 (
            .O(N__23423),
            .I(N__23410));
    InMux I__4468 (
            .O(N__23420),
            .I(N__23410));
    Odrv4 I__4467 (
            .O(N__23417),
            .I(b2v_inst_state_8));
    LocalMux I__4466 (
            .O(N__23410),
            .I(b2v_inst_state_8));
    InMux I__4465 (
            .O(N__23405),
            .I(N__23401));
    IoInMux I__4464 (
            .O(N__23404),
            .I(N__23398));
    LocalMux I__4463 (
            .O(N__23401),
            .I(N__23395));
    LocalMux I__4462 (
            .O(N__23398),
            .I(N__23392));
    Span4Mux_v I__4461 (
            .O(N__23395),
            .I(N__23389));
    Span12Mux_s6_v I__4460 (
            .O(N__23392),
            .I(N__23386));
    Span4Mux_h I__4459 (
            .O(N__23389),
            .I(N__23383));
    Span12Mux_v I__4458 (
            .O(N__23386),
            .I(N__23380));
    Span4Mux_h I__4457 (
            .O(N__23383),
            .I(N__23377));
    Odrv12 I__4456 (
            .O(N__23380),
            .I(leds_c_0));
    Odrv4 I__4455 (
            .O(N__23377),
            .I(leds_c_0));
    IoInMux I__4454 (
            .O(N__23372),
            .I(N__23368));
    InMux I__4453 (
            .O(N__23371),
            .I(N__23365));
    LocalMux I__4452 (
            .O(N__23368),
            .I(N__23362));
    LocalMux I__4451 (
            .O(N__23365),
            .I(N__23359));
    Span4Mux_s3_h I__4450 (
            .O(N__23362),
            .I(N__23356));
    Span4Mux_h I__4449 (
            .O(N__23359),
            .I(N__23353));
    Span4Mux_v I__4448 (
            .O(N__23356),
            .I(N__23350));
    Span4Mux_h I__4447 (
            .O(N__23353),
            .I(N__23347));
    Span4Mux_v I__4446 (
            .O(N__23350),
            .I(N__23344));
    Span4Mux_h I__4445 (
            .O(N__23347),
            .I(N__23341));
    Span4Mux_h I__4444 (
            .O(N__23344),
            .I(N__23336));
    Span4Mux_v I__4443 (
            .O(N__23341),
            .I(N__23336));
    Odrv4 I__4442 (
            .O(N__23336),
            .I(leds_c_1));
    InMux I__4441 (
            .O(N__23333),
            .I(N__23329));
    IoInMux I__4440 (
            .O(N__23332),
            .I(N__23326));
    LocalMux I__4439 (
            .O(N__23329),
            .I(N__23323));
    LocalMux I__4438 (
            .O(N__23326),
            .I(N__23320));
    Span4Mux_v I__4437 (
            .O(N__23323),
            .I(N__23317));
    Span4Mux_s3_h I__4436 (
            .O(N__23320),
            .I(N__23314));
    Span4Mux_h I__4435 (
            .O(N__23317),
            .I(N__23311));
    Span4Mux_h I__4434 (
            .O(N__23314),
            .I(N__23308));
    Span4Mux_h I__4433 (
            .O(N__23311),
            .I(N__23305));
    Odrv4 I__4432 (
            .O(N__23308),
            .I(leds_c_13));
    Odrv4 I__4431 (
            .O(N__23305),
            .I(leds_c_13));
    InMux I__4430 (
            .O(N__23300),
            .I(N__23293));
    InMux I__4429 (
            .O(N__23299),
            .I(N__23288));
    InMux I__4428 (
            .O(N__23298),
            .I(N__23288));
    InMux I__4427 (
            .O(N__23297),
            .I(N__23285));
    InMux I__4426 (
            .O(N__23296),
            .I(N__23282));
    LocalMux I__4425 (
            .O(N__23293),
            .I(\b2v_inst.cuentaZ0Z_0 ));
    LocalMux I__4424 (
            .O(N__23288),
            .I(\b2v_inst.cuentaZ0Z_0 ));
    LocalMux I__4423 (
            .O(N__23285),
            .I(\b2v_inst.cuentaZ0Z_0 ));
    LocalMux I__4422 (
            .O(N__23282),
            .I(\b2v_inst.cuentaZ0Z_0 ));
    InMux I__4421 (
            .O(N__23273),
            .I(N__23269));
    CascadeMux I__4420 (
            .O(N__23272),
            .I(N__23265));
    LocalMux I__4419 (
            .O(N__23269),
            .I(N__23262));
    InMux I__4418 (
            .O(N__23268),
            .I(N__23259));
    InMux I__4417 (
            .O(N__23265),
            .I(N__23256));
    Odrv4 I__4416 (
            .O(N__23262),
            .I(\b2v_inst.cuentaZ0Z_1 ));
    LocalMux I__4415 (
            .O(N__23259),
            .I(\b2v_inst.cuentaZ0Z_1 ));
    LocalMux I__4414 (
            .O(N__23256),
            .I(\b2v_inst.cuentaZ0Z_1 ));
    CascadeMux I__4413 (
            .O(N__23249),
            .I(N__23245));
    InMux I__4412 (
            .O(N__23248),
            .I(N__23242));
    InMux I__4411 (
            .O(N__23245),
            .I(N__23239));
    LocalMux I__4410 (
            .O(N__23242),
            .I(\b2v_inst.cuentaZ0Z_2 ));
    LocalMux I__4409 (
            .O(N__23239),
            .I(\b2v_inst.cuentaZ0Z_2 ));
    InMux I__4408 (
            .O(N__23234),
            .I(N__23230));
    InMux I__4407 (
            .O(N__23233),
            .I(N__23227));
    LocalMux I__4406 (
            .O(N__23230),
            .I(N__23224));
    LocalMux I__4405 (
            .O(N__23227),
            .I(\b2v_inst.un4_cuenta_cry_1_c_RNI9VZ0Z48 ));
    Odrv4 I__4404 (
            .O(N__23224),
            .I(\b2v_inst.un4_cuenta_cry_1_c_RNI9VZ0Z48 ));
    InMux I__4403 (
            .O(N__23219),
            .I(\b2v_inst.un4_cuenta_cry_1 ));
    CascadeMux I__4402 (
            .O(N__23216),
            .I(N__23212));
    InMux I__4401 (
            .O(N__23215),
            .I(N__23209));
    InMux I__4400 (
            .O(N__23212),
            .I(N__23206));
    LocalMux I__4399 (
            .O(N__23209),
            .I(\b2v_inst.cuentaZ0Z_3 ));
    LocalMux I__4398 (
            .O(N__23206),
            .I(\b2v_inst.cuentaZ0Z_3 ));
    InMux I__4397 (
            .O(N__23201),
            .I(N__23197));
    InMux I__4396 (
            .O(N__23200),
            .I(N__23194));
    LocalMux I__4395 (
            .O(N__23197),
            .I(\b2v_inst.un4_cuenta_cry_2_c_RNIBZ0Z268 ));
    LocalMux I__4394 (
            .O(N__23194),
            .I(\b2v_inst.un4_cuenta_cry_2_c_RNIBZ0Z268 ));
    InMux I__4393 (
            .O(N__23189),
            .I(\b2v_inst.un4_cuenta_cry_2 ));
    CascadeMux I__4392 (
            .O(N__23186),
            .I(N__23182));
    InMux I__4391 (
            .O(N__23185),
            .I(N__23179));
    InMux I__4390 (
            .O(N__23182),
            .I(N__23176));
    LocalMux I__4389 (
            .O(N__23179),
            .I(\b2v_inst.cuentaZ0Z_4 ));
    LocalMux I__4388 (
            .O(N__23176),
            .I(\b2v_inst.cuentaZ0Z_4 ));
    InMux I__4387 (
            .O(N__23171),
            .I(N__23167));
    InMux I__4386 (
            .O(N__23170),
            .I(N__23164));
    LocalMux I__4385 (
            .O(N__23167),
            .I(\b2v_inst.un4_cuenta_cry_3_c_RNIDZ0Z578 ));
    LocalMux I__4384 (
            .O(N__23164),
            .I(\b2v_inst.un4_cuenta_cry_3_c_RNIDZ0Z578 ));
    InMux I__4383 (
            .O(N__23159),
            .I(\b2v_inst.un4_cuenta_cry_3 ));
    InMux I__4382 (
            .O(N__23156),
            .I(\b2v_inst.un4_cuenta_cry_4 ));
    InMux I__4381 (
            .O(N__23153),
            .I(N__23149));
    InMux I__4380 (
            .O(N__23152),
            .I(N__23146));
    LocalMux I__4379 (
            .O(N__23149),
            .I(N__23141));
    LocalMux I__4378 (
            .O(N__23146),
            .I(N__23141));
    Span4Mux_v I__4377 (
            .O(N__23141),
            .I(N__23138));
    Odrv4 I__4376 (
            .O(N__23138),
            .I(\b2v_inst.cuentaZ0Z_6 ));
    InMux I__4375 (
            .O(N__23135),
            .I(N__23132));
    LocalMux I__4374 (
            .O(N__23132),
            .I(N__23128));
    InMux I__4373 (
            .O(N__23131),
            .I(N__23125));
    Odrv12 I__4372 (
            .O(N__23128),
            .I(\b2v_inst.un4_cuenta_cry_5_c_RNIHBZ0Z98 ));
    LocalMux I__4371 (
            .O(N__23125),
            .I(\b2v_inst.un4_cuenta_cry_5_c_RNIHBZ0Z98 ));
    InMux I__4370 (
            .O(N__23120),
            .I(\b2v_inst.un4_cuenta_cry_5 ));
    CascadeMux I__4369 (
            .O(N__23117),
            .I(N__23113));
    InMux I__4368 (
            .O(N__23116),
            .I(N__23110));
    InMux I__4367 (
            .O(N__23113),
            .I(N__23107));
    LocalMux I__4366 (
            .O(N__23110),
            .I(N__23104));
    LocalMux I__4365 (
            .O(N__23107),
            .I(N__23099));
    Span4Mux_v I__4364 (
            .O(N__23104),
            .I(N__23099));
    Odrv4 I__4363 (
            .O(N__23099),
            .I(\b2v_inst.cuentaZ0Z_7 ));
    InMux I__4362 (
            .O(N__23096),
            .I(N__23093));
    LocalMux I__4361 (
            .O(N__23093),
            .I(N__23089));
    InMux I__4360 (
            .O(N__23092),
            .I(N__23086));
    Odrv12 I__4359 (
            .O(N__23089),
            .I(\b2v_inst.un4_cuenta_cry_6_c_RNIJEAZ0Z8 ));
    LocalMux I__4358 (
            .O(N__23086),
            .I(\b2v_inst.un4_cuenta_cry_6_c_RNIJEAZ0Z8 ));
    InMux I__4357 (
            .O(N__23081),
            .I(\b2v_inst.un4_cuenta_cry_6 ));
    InMux I__4356 (
            .O(N__23078),
            .I(N__23075));
    LocalMux I__4355 (
            .O(N__23075),
            .I(N__23071));
    InMux I__4354 (
            .O(N__23074),
            .I(N__23068));
    Span4Mux_v I__4353 (
            .O(N__23071),
            .I(N__23065));
    LocalMux I__4352 (
            .O(N__23068),
            .I(\b2v_inst.cuentaZ0Z_8 ));
    Odrv4 I__4351 (
            .O(N__23065),
            .I(\b2v_inst.cuentaZ0Z_8 ));
    InMux I__4350 (
            .O(N__23060),
            .I(N__23057));
    LocalMux I__4349 (
            .O(N__23057),
            .I(N__23052));
    InMux I__4348 (
            .O(N__23056),
            .I(N__23047));
    InMux I__4347 (
            .O(N__23055),
            .I(N__23047));
    Odrv12 I__4346 (
            .O(N__23052),
            .I(\b2v_inst.un4_cuenta_cry_7_c_RNILHBZ0Z8 ));
    LocalMux I__4345 (
            .O(N__23047),
            .I(\b2v_inst.un4_cuenta_cry_7_c_RNILHBZ0Z8 ));
    InMux I__4344 (
            .O(N__23042),
            .I(\b2v_inst.un4_cuenta_cry_7 ));
    CascadeMux I__4343 (
            .O(N__23039),
            .I(\b2v_inst9.data_to_send_10_0_0_0_3_cascade_ ));
    CascadeMux I__4342 (
            .O(N__23036),
            .I(N__23033));
    InMux I__4341 (
            .O(N__23033),
            .I(N__23030));
    LocalMux I__4340 (
            .O(N__23030),
            .I(\b2v_inst9.data_to_sendZ0Z_6 ));
    InMux I__4339 (
            .O(N__23027),
            .I(N__23024));
    LocalMux I__4338 (
            .O(N__23024),
            .I(\b2v_inst.un1_data_a_escribir_0_sqmuxa_3_i_i_a2_0 ));
    CascadeMux I__4337 (
            .O(N__23021),
            .I(\b2v_inst.N_655_cascade_ ));
    InMux I__4336 (
            .O(N__23018),
            .I(N__23011));
    InMux I__4335 (
            .O(N__23017),
            .I(N__23006));
    InMux I__4334 (
            .O(N__23016),
            .I(N__23006));
    CascadeMux I__4333 (
            .O(N__23015),
            .I(N__23001));
    CascadeMux I__4332 (
            .O(N__23014),
            .I(N__22997));
    LocalMux I__4331 (
            .O(N__23011),
            .I(N__22989));
    LocalMux I__4330 (
            .O(N__23006),
            .I(N__22986));
    InMux I__4329 (
            .O(N__23005),
            .I(N__22979));
    InMux I__4328 (
            .O(N__23004),
            .I(N__22979));
    InMux I__4327 (
            .O(N__23001),
            .I(N__22979));
    InMux I__4326 (
            .O(N__23000),
            .I(N__22972));
    InMux I__4325 (
            .O(N__22997),
            .I(N__22972));
    InMux I__4324 (
            .O(N__22996),
            .I(N__22972));
    CascadeMux I__4323 (
            .O(N__22995),
            .I(N__22969));
    InMux I__4322 (
            .O(N__22994),
            .I(N__22963));
    InMux I__4321 (
            .O(N__22993),
            .I(N__22963));
    InMux I__4320 (
            .O(N__22992),
            .I(N__22960));
    Span4Mux_h I__4319 (
            .O(N__22989),
            .I(N__22951));
    Span4Mux_h I__4318 (
            .O(N__22986),
            .I(N__22951));
    LocalMux I__4317 (
            .O(N__22979),
            .I(N__22951));
    LocalMux I__4316 (
            .O(N__22972),
            .I(N__22951));
    InMux I__4315 (
            .O(N__22969),
            .I(N__22946));
    InMux I__4314 (
            .O(N__22968),
            .I(N__22946));
    LocalMux I__4313 (
            .O(N__22963),
            .I(\b2v_inst.state18_li_0 ));
    LocalMux I__4312 (
            .O(N__22960),
            .I(\b2v_inst.state18_li_0 ));
    Odrv4 I__4311 (
            .O(N__22951),
            .I(\b2v_inst.state18_li_0 ));
    LocalMux I__4310 (
            .O(N__22946),
            .I(\b2v_inst.state18_li_0 ));
    InMux I__4309 (
            .O(N__22937),
            .I(N__22933));
    InMux I__4308 (
            .O(N__22936),
            .I(N__22930));
    LocalMux I__4307 (
            .O(N__22933),
            .I(\b2v_inst.cuenta_RNIR03AZ0Z_1 ));
    LocalMux I__4306 (
            .O(N__22930),
            .I(\b2v_inst.cuenta_RNIR03AZ0Z_1 ));
    CascadeMux I__4305 (
            .O(N__22925),
            .I(N__22920));
    CascadeMux I__4304 (
            .O(N__22924),
            .I(N__22917));
    CascadeMux I__4303 (
            .O(N__22923),
            .I(N__22912));
    InMux I__4302 (
            .O(N__22920),
            .I(N__22909));
    InMux I__4301 (
            .O(N__22917),
            .I(N__22904));
    InMux I__4300 (
            .O(N__22916),
            .I(N__22897));
    InMux I__4299 (
            .O(N__22915),
            .I(N__22897));
    InMux I__4298 (
            .O(N__22912),
            .I(N__22897));
    LocalMux I__4297 (
            .O(N__22909),
            .I(N__22894));
    InMux I__4296 (
            .O(N__22908),
            .I(N__22890));
    InMux I__4295 (
            .O(N__22907),
            .I(N__22887));
    LocalMux I__4294 (
            .O(N__22904),
            .I(N__22884));
    LocalMux I__4293 (
            .O(N__22897),
            .I(N__22881));
    Span4Mux_v I__4292 (
            .O(N__22894),
            .I(N__22878));
    InMux I__4291 (
            .O(N__22893),
            .I(N__22875));
    LocalMux I__4290 (
            .O(N__22890),
            .I(N__22872));
    LocalMux I__4289 (
            .O(N__22887),
            .I(N__22869));
    Span4Mux_v I__4288 (
            .O(N__22884),
            .I(N__22864));
    Span4Mux_h I__4287 (
            .O(N__22881),
            .I(N__22864));
    Span4Mux_h I__4286 (
            .O(N__22878),
            .I(N__22859));
    LocalMux I__4285 (
            .O(N__22875),
            .I(N__22856));
    Span12Mux_h I__4284 (
            .O(N__22872),
            .I(N__22853));
    Span4Mux_h I__4283 (
            .O(N__22869),
            .I(N__22848));
    Span4Mux_h I__4282 (
            .O(N__22864),
            .I(N__22848));
    InMux I__4281 (
            .O(N__22863),
            .I(N__22843));
    InMux I__4280 (
            .O(N__22862),
            .I(N__22843));
    Odrv4 I__4279 (
            .O(N__22859),
            .I(\b2v_inst1.r_SM_MainZ0Z_1 ));
    Odrv12 I__4278 (
            .O(N__22856),
            .I(\b2v_inst1.r_SM_MainZ0Z_1 ));
    Odrv12 I__4277 (
            .O(N__22853),
            .I(\b2v_inst1.r_SM_MainZ0Z_1 ));
    Odrv4 I__4276 (
            .O(N__22848),
            .I(\b2v_inst1.r_SM_MainZ0Z_1 ));
    LocalMux I__4275 (
            .O(N__22843),
            .I(\b2v_inst1.r_SM_MainZ0Z_1 ));
    InMux I__4274 (
            .O(N__22832),
            .I(N__22823));
    InMux I__4273 (
            .O(N__22831),
            .I(N__22820));
    InMux I__4272 (
            .O(N__22830),
            .I(N__22817));
    InMux I__4271 (
            .O(N__22829),
            .I(N__22813));
    InMux I__4270 (
            .O(N__22828),
            .I(N__22809));
    InMux I__4269 (
            .O(N__22827),
            .I(N__22804));
    InMux I__4268 (
            .O(N__22826),
            .I(N__22804));
    LocalMux I__4267 (
            .O(N__22823),
            .I(N__22801));
    LocalMux I__4266 (
            .O(N__22820),
            .I(N__22796));
    LocalMux I__4265 (
            .O(N__22817),
            .I(N__22796));
    InMux I__4264 (
            .O(N__22816),
            .I(N__22793));
    LocalMux I__4263 (
            .O(N__22813),
            .I(N__22790));
    InMux I__4262 (
            .O(N__22812),
            .I(N__22787));
    LocalMux I__4261 (
            .O(N__22809),
            .I(N__22782));
    LocalMux I__4260 (
            .O(N__22804),
            .I(N__22777));
    Span4Mux_h I__4259 (
            .O(N__22801),
            .I(N__22777));
    Span4Mux_v I__4258 (
            .O(N__22796),
            .I(N__22770));
    LocalMux I__4257 (
            .O(N__22793),
            .I(N__22770));
    Span4Mux_h I__4256 (
            .O(N__22790),
            .I(N__22770));
    LocalMux I__4255 (
            .O(N__22787),
            .I(N__22767));
    InMux I__4254 (
            .O(N__22786),
            .I(N__22762));
    InMux I__4253 (
            .O(N__22785),
            .I(N__22762));
    Span4Mux_h I__4252 (
            .O(N__22782),
            .I(N__22759));
    Span4Mux_h I__4251 (
            .O(N__22777),
            .I(N__22756));
    Span4Mux_h I__4250 (
            .O(N__22770),
            .I(N__22753));
    Span12Mux_h I__4249 (
            .O(N__22767),
            .I(N__22748));
    LocalMux I__4248 (
            .O(N__22762),
            .I(N__22748));
    Odrv4 I__4247 (
            .O(N__22759),
            .I(\b2v_inst1.r_RX_DataZ0 ));
    Odrv4 I__4246 (
            .O(N__22756),
            .I(\b2v_inst1.r_RX_DataZ0 ));
    Odrv4 I__4245 (
            .O(N__22753),
            .I(\b2v_inst1.r_RX_DataZ0 ));
    Odrv12 I__4244 (
            .O(N__22748),
            .I(\b2v_inst1.r_RX_DataZ0 ));
    InMux I__4243 (
            .O(N__22739),
            .I(N__22734));
    InMux I__4242 (
            .O(N__22738),
            .I(N__22728));
    InMux I__4241 (
            .O(N__22737),
            .I(N__22728));
    LocalMux I__4240 (
            .O(N__22734),
            .I(N__22725));
    CascadeMux I__4239 (
            .O(N__22733),
            .I(N__22721));
    LocalMux I__4238 (
            .O(N__22728),
            .I(N__22717));
    Span4Mux_h I__4237 (
            .O(N__22725),
            .I(N__22714));
    InMux I__4236 (
            .O(N__22724),
            .I(N__22710));
    InMux I__4235 (
            .O(N__22721),
            .I(N__22707));
    InMux I__4234 (
            .O(N__22720),
            .I(N__22704));
    Span4Mux_v I__4233 (
            .O(N__22717),
            .I(N__22701));
    Span4Mux_h I__4232 (
            .O(N__22714),
            .I(N__22698));
    InMux I__4231 (
            .O(N__22713),
            .I(N__22695));
    LocalMux I__4230 (
            .O(N__22710),
            .I(N__22690));
    LocalMux I__4229 (
            .O(N__22707),
            .I(N__22690));
    LocalMux I__4228 (
            .O(N__22704),
            .I(N__22685));
    Span4Mux_h I__4227 (
            .O(N__22701),
            .I(N__22685));
    Odrv4 I__4226 (
            .O(N__22698),
            .I(\b2v_inst1.r_SM_MainZ0Z_2 ));
    LocalMux I__4225 (
            .O(N__22695),
            .I(\b2v_inst1.r_SM_MainZ0Z_2 ));
    Odrv4 I__4224 (
            .O(N__22690),
            .I(\b2v_inst1.r_SM_MainZ0Z_2 ));
    Odrv4 I__4223 (
            .O(N__22685),
            .I(\b2v_inst1.r_SM_MainZ0Z_2 ));
    InMux I__4222 (
            .O(N__22676),
            .I(N__22673));
    LocalMux I__4221 (
            .O(N__22673),
            .I(N__22670));
    Span4Mux_v I__4220 (
            .O(N__22670),
            .I(N__22667));
    Span4Mux_h I__4219 (
            .O(N__22667),
            .I(N__22664));
    Odrv4 I__4218 (
            .O(N__22664),
            .I(\b2v_inst1.m13_i_2 ));
    CascadeMux I__4217 (
            .O(N__22661),
            .I(\b2v_inst1.N_95_cascade_ ));
    InMux I__4216 (
            .O(N__22658),
            .I(N__22655));
    LocalMux I__4215 (
            .O(N__22655),
            .I(N__22652));
    Span4Mux_v I__4214 (
            .O(N__22652),
            .I(N__22649));
    Span4Mux_h I__4213 (
            .O(N__22649),
            .I(N__22646));
    Odrv4 I__4212 (
            .O(N__22646),
            .I(\b2v_inst1.N_96 ));
    InMux I__4211 (
            .O(N__22643),
            .I(N__22639));
    InMux I__4210 (
            .O(N__22642),
            .I(N__22635));
    LocalMux I__4209 (
            .O(N__22639),
            .I(N__22631));
    InMux I__4208 (
            .O(N__22638),
            .I(N__22628));
    LocalMux I__4207 (
            .O(N__22635),
            .I(N__22621));
    InMux I__4206 (
            .O(N__22634),
            .I(N__22616));
    Span4Mux_v I__4205 (
            .O(N__22631),
            .I(N__22611));
    LocalMux I__4204 (
            .O(N__22628),
            .I(N__22611));
    InMux I__4203 (
            .O(N__22627),
            .I(N__22608));
    InMux I__4202 (
            .O(N__22626),
            .I(N__22601));
    InMux I__4201 (
            .O(N__22625),
            .I(N__22601));
    InMux I__4200 (
            .O(N__22624),
            .I(N__22601));
    Span4Mux_h I__4199 (
            .O(N__22621),
            .I(N__22598));
    InMux I__4198 (
            .O(N__22620),
            .I(N__22593));
    InMux I__4197 (
            .O(N__22619),
            .I(N__22593));
    LocalMux I__4196 (
            .O(N__22616),
            .I(N__22590));
    Span4Mux_v I__4195 (
            .O(N__22611),
            .I(N__22583));
    LocalMux I__4194 (
            .O(N__22608),
            .I(N__22583));
    LocalMux I__4193 (
            .O(N__22601),
            .I(N__22583));
    Span4Mux_h I__4192 (
            .O(N__22598),
            .I(N__22580));
    LocalMux I__4191 (
            .O(N__22593),
            .I(N__22577));
    Span4Mux_h I__4190 (
            .O(N__22590),
            .I(N__22574));
    Span4Mux_v I__4189 (
            .O(N__22583),
            .I(N__22570));
    Span4Mux_v I__4188 (
            .O(N__22580),
            .I(N__22567));
    Span4Mux_v I__4187 (
            .O(N__22577),
            .I(N__22564));
    Span4Mux_h I__4186 (
            .O(N__22574),
            .I(N__22561));
    InMux I__4185 (
            .O(N__22573),
            .I(N__22558));
    Span4Mux_h I__4184 (
            .O(N__22570),
            .I(N__22555));
    Odrv4 I__4183 (
            .O(N__22567),
            .I(\b2v_inst1.r_SM_MainZ0Z_0 ));
    Odrv4 I__4182 (
            .O(N__22564),
            .I(\b2v_inst1.r_SM_MainZ0Z_0 ));
    Odrv4 I__4181 (
            .O(N__22561),
            .I(\b2v_inst1.r_SM_MainZ0Z_0 ));
    LocalMux I__4180 (
            .O(N__22558),
            .I(\b2v_inst1.r_SM_MainZ0Z_0 ));
    Odrv4 I__4179 (
            .O(N__22555),
            .I(\b2v_inst1.r_SM_MainZ0Z_0 ));
    InMux I__4178 (
            .O(N__22544),
            .I(N__22541));
    LocalMux I__4177 (
            .O(N__22541),
            .I(N__22538));
    Span4Mux_v I__4176 (
            .O(N__22538),
            .I(N__22535));
    Odrv4 I__4175 (
            .O(N__22535),
            .I(\b2v_inst.dir_memZ0Z_5 ));
    CascadeMux I__4174 (
            .O(N__22532),
            .I(N__22528));
    InMux I__4173 (
            .O(N__22531),
            .I(N__22520));
    InMux I__4172 (
            .O(N__22528),
            .I(N__22515));
    InMux I__4171 (
            .O(N__22527),
            .I(N__22515));
    InMux I__4170 (
            .O(N__22526),
            .I(N__22512));
    InMux I__4169 (
            .O(N__22525),
            .I(N__22508));
    InMux I__4168 (
            .O(N__22524),
            .I(N__22505));
    InMux I__4167 (
            .O(N__22523),
            .I(N__22502));
    LocalMux I__4166 (
            .O(N__22520),
            .I(N__22494));
    LocalMux I__4165 (
            .O(N__22515),
            .I(N__22494));
    LocalMux I__4164 (
            .O(N__22512),
            .I(N__22491));
    InMux I__4163 (
            .O(N__22511),
            .I(N__22488));
    LocalMux I__4162 (
            .O(N__22508),
            .I(N__22481));
    LocalMux I__4161 (
            .O(N__22505),
            .I(N__22481));
    LocalMux I__4160 (
            .O(N__22502),
            .I(N__22481));
    InMux I__4159 (
            .O(N__22501),
            .I(N__22476));
    InMux I__4158 (
            .O(N__22500),
            .I(N__22476));
    InMux I__4157 (
            .O(N__22499),
            .I(N__22473));
    Odrv4 I__4156 (
            .O(N__22494),
            .I(\b2v_inst.N_450_i_1 ));
    Odrv4 I__4155 (
            .O(N__22491),
            .I(\b2v_inst.N_450_i_1 ));
    LocalMux I__4154 (
            .O(N__22488),
            .I(\b2v_inst.N_450_i_1 ));
    Odrv4 I__4153 (
            .O(N__22481),
            .I(\b2v_inst.N_450_i_1 ));
    LocalMux I__4152 (
            .O(N__22476),
            .I(\b2v_inst.N_450_i_1 ));
    LocalMux I__4151 (
            .O(N__22473),
            .I(\b2v_inst.N_450_i_1 ));
    CascadeMux I__4150 (
            .O(N__22460),
            .I(N__22457));
    InMux I__4149 (
            .O(N__22457),
            .I(N__22454));
    LocalMux I__4148 (
            .O(N__22454),
            .I(N__22451));
    Span4Mux_h I__4147 (
            .O(N__22451),
            .I(N__22448));
    Odrv4 I__4146 (
            .O(N__22448),
            .I(\b2v_inst.dir_mem_2Z0Z_5 ));
    CascadeMux I__4145 (
            .O(N__22445),
            .I(N__22440));
    InMux I__4144 (
            .O(N__22444),
            .I(N__22435));
    InMux I__4143 (
            .O(N__22443),
            .I(N__22432));
    InMux I__4142 (
            .O(N__22440),
            .I(N__22426));
    InMux I__4141 (
            .O(N__22439),
            .I(N__22421));
    InMux I__4140 (
            .O(N__22438),
            .I(N__22421));
    LocalMux I__4139 (
            .O(N__22435),
            .I(N__22415));
    LocalMux I__4138 (
            .O(N__22432),
            .I(N__22415));
    InMux I__4137 (
            .O(N__22431),
            .I(N__22410));
    InMux I__4136 (
            .O(N__22430),
            .I(N__22410));
    InMux I__4135 (
            .O(N__22429),
            .I(N__22407));
    LocalMux I__4134 (
            .O(N__22426),
            .I(N__22399));
    LocalMux I__4133 (
            .O(N__22421),
            .I(N__22399));
    InMux I__4132 (
            .O(N__22420),
            .I(N__22396));
    Span4Mux_v I__4131 (
            .O(N__22415),
            .I(N__22389));
    LocalMux I__4130 (
            .O(N__22410),
            .I(N__22389));
    LocalMux I__4129 (
            .O(N__22407),
            .I(N__22389));
    InMux I__4128 (
            .O(N__22406),
            .I(N__22386));
    InMux I__4127 (
            .O(N__22405),
            .I(N__22381));
    InMux I__4126 (
            .O(N__22404),
            .I(N__22381));
    Odrv4 I__4125 (
            .O(N__22399),
            .I(\b2v_inst.N_489 ));
    LocalMux I__4124 (
            .O(N__22396),
            .I(\b2v_inst.N_489 ));
    Odrv4 I__4123 (
            .O(N__22389),
            .I(\b2v_inst.N_489 ));
    LocalMux I__4122 (
            .O(N__22386),
            .I(\b2v_inst.N_489 ));
    LocalMux I__4121 (
            .O(N__22381),
            .I(\b2v_inst.N_489 ));
    CascadeMux I__4120 (
            .O(N__22370),
            .I(\b2v_inst9.data_to_send_10_0_0_0_5_cascade_ ));
    CascadeMux I__4119 (
            .O(N__22367),
            .I(N__22364));
    InMux I__4118 (
            .O(N__22364),
            .I(N__22361));
    LocalMux I__4117 (
            .O(N__22361),
            .I(\b2v_inst9.data_to_sendZ0Z_5 ));
    CascadeMux I__4116 (
            .O(N__22358),
            .I(N__22355));
    InMux I__4115 (
            .O(N__22355),
            .I(N__22352));
    LocalMux I__4114 (
            .O(N__22352),
            .I(N__22349));
    Odrv4 I__4113 (
            .O(N__22349),
            .I(\b2v_inst.dir_mem_2_RNO_0Z0Z_5 ));
    InMux I__4112 (
            .O(N__22346),
            .I(\b2v_inst.un2_dir_mem_2_cry_4 ));
    CascadeMux I__4111 (
            .O(N__22343),
            .I(N__22340));
    InMux I__4110 (
            .O(N__22340),
            .I(N__22337));
    LocalMux I__4109 (
            .O(N__22337),
            .I(N__22334));
    Odrv4 I__4108 (
            .O(N__22334),
            .I(\b2v_inst.dir_mem_2_RNO_0Z0Z_6 ));
    InMux I__4107 (
            .O(N__22331),
            .I(\b2v_inst.un2_dir_mem_2_cry_5 ));
    CascadeMux I__4106 (
            .O(N__22328),
            .I(N__22325));
    InMux I__4105 (
            .O(N__22325),
            .I(N__22322));
    LocalMux I__4104 (
            .O(N__22322),
            .I(N__22319));
    Odrv4 I__4103 (
            .O(N__22319),
            .I(\b2v_inst.dir_mem_2_RNO_0Z0Z_7 ));
    InMux I__4102 (
            .O(N__22316),
            .I(\b2v_inst.un2_dir_mem_2_cry_6 ));
    InMux I__4101 (
            .O(N__22313),
            .I(N__22310));
    LocalMux I__4100 (
            .O(N__22310),
            .I(N__22307));
    Odrv4 I__4099 (
            .O(N__22307),
            .I(\b2v_inst.dir_mem_2_RNO_0Z0Z_8 ));
    InMux I__4098 (
            .O(N__22304),
            .I(bfn_13_7_0_));
    CascadeMux I__4097 (
            .O(N__22301),
            .I(N__22298));
    InMux I__4096 (
            .O(N__22298),
            .I(N__22295));
    LocalMux I__4095 (
            .O(N__22295),
            .I(\b2v_inst.dir_mem_2_RNO_0Z0Z_9 ));
    InMux I__4094 (
            .O(N__22292),
            .I(\b2v_inst.un2_dir_mem_2_cry_8 ));
    InMux I__4093 (
            .O(N__22289),
            .I(\b2v_inst.un2_dir_mem_2_cry_9 ));
    CascadeMux I__4092 (
            .O(N__22286),
            .I(N__22283));
    InMux I__4091 (
            .O(N__22283),
            .I(N__22280));
    LocalMux I__4090 (
            .O(N__22280),
            .I(\b2v_inst.dir_mem_2_RNO_0Z0Z_10 ));
    InMux I__4089 (
            .O(N__22277),
            .I(N__22274));
    LocalMux I__4088 (
            .O(N__22274),
            .I(\b2v_inst1.r_RX_Data_RZ0 ));
    CascadeMux I__4087 (
            .O(N__22271),
            .I(N__22267));
    InMux I__4086 (
            .O(N__22270),
            .I(N__22259));
    InMux I__4085 (
            .O(N__22267),
            .I(N__22259));
    InMux I__4084 (
            .O(N__22266),
            .I(N__22259));
    LocalMux I__4083 (
            .O(N__22259),
            .I(N__22256));
    Sp12to4 I__4082 (
            .O(N__22256),
            .I(N__22253));
    Odrv12 I__4081 (
            .O(N__22253),
            .I(\b2v_inst.un9_indice_0_a2_2 ));
    CascadeMux I__4080 (
            .O(N__22250),
            .I(N__22245));
    InMux I__4079 (
            .O(N__22249),
            .I(N__22238));
    InMux I__4078 (
            .O(N__22248),
            .I(N__22238));
    InMux I__4077 (
            .O(N__22245),
            .I(N__22238));
    LocalMux I__4076 (
            .O(N__22238),
            .I(N__22234));
    InMux I__4075 (
            .O(N__22237),
            .I(N__22231));
    Span4Mux_h I__4074 (
            .O(N__22234),
            .I(N__22228));
    LocalMux I__4073 (
            .O(N__22231),
            .I(N__22225));
    Span4Mux_v I__4072 (
            .O(N__22228),
            .I(N__22222));
    Span4Mux_v I__4071 (
            .O(N__22225),
            .I(N__22217));
    Span4Mux_v I__4070 (
            .O(N__22222),
            .I(N__22217));
    Odrv4 I__4069 (
            .O(N__22217),
            .I(\b2v_inst.un9_indice_0_a2_3 ));
    InMux I__4068 (
            .O(N__22214),
            .I(N__22211));
    LocalMux I__4067 (
            .O(N__22211),
            .I(N__22208));
    Span4Mux_h I__4066 (
            .O(N__22208),
            .I(N__22205));
    Span4Mux_h I__4065 (
            .O(N__22205),
            .I(N__22202));
    Odrv4 I__4064 (
            .O(N__22202),
            .I(\b2v_inst.dir_mem_RNO_0Z0Z_5 ));
    CascadeMux I__4063 (
            .O(N__22199),
            .I(\b2v_inst.un9_indice_0_a2_2_cascade_ ));
    CEMux I__4062 (
            .O(N__22196),
            .I(N__22192));
    CEMux I__4061 (
            .O(N__22195),
            .I(N__22189));
    LocalMux I__4060 (
            .O(N__22192),
            .I(N__22183));
    LocalMux I__4059 (
            .O(N__22189),
            .I(N__22180));
    CEMux I__4058 (
            .O(N__22188),
            .I(N__22177));
    CEMux I__4057 (
            .O(N__22187),
            .I(N__22174));
    CEMux I__4056 (
            .O(N__22186),
            .I(N__22171));
    Span4Mux_v I__4055 (
            .O(N__22183),
            .I(N__22166));
    Span4Mux_v I__4054 (
            .O(N__22180),
            .I(N__22163));
    LocalMux I__4053 (
            .O(N__22177),
            .I(N__22160));
    LocalMux I__4052 (
            .O(N__22174),
            .I(N__22157));
    LocalMux I__4051 (
            .O(N__22171),
            .I(N__22154));
    CEMux I__4050 (
            .O(N__22170),
            .I(N__22151));
    CascadeMux I__4049 (
            .O(N__22169),
            .I(N__22146));
    Span4Mux_h I__4048 (
            .O(N__22166),
            .I(N__22139));
    Span4Mux_h I__4047 (
            .O(N__22163),
            .I(N__22139));
    Span4Mux_h I__4046 (
            .O(N__22160),
            .I(N__22139));
    Span4Mux_v I__4045 (
            .O(N__22157),
            .I(N__22136));
    Span4Mux_h I__4044 (
            .O(N__22154),
            .I(N__22131));
    LocalMux I__4043 (
            .O(N__22151),
            .I(N__22131));
    InMux I__4042 (
            .O(N__22150),
            .I(N__22128));
    InMux I__4041 (
            .O(N__22149),
            .I(N__22125));
    InMux I__4040 (
            .O(N__22146),
            .I(N__22122));
    Odrv4 I__4039 (
            .O(N__22139),
            .I(\b2v_inst.stateZ0Z_28 ));
    Odrv4 I__4038 (
            .O(N__22136),
            .I(\b2v_inst.stateZ0Z_28 ));
    Odrv4 I__4037 (
            .O(N__22131),
            .I(\b2v_inst.stateZ0Z_28 ));
    LocalMux I__4036 (
            .O(N__22128),
            .I(\b2v_inst.stateZ0Z_28 ));
    LocalMux I__4035 (
            .O(N__22125),
            .I(\b2v_inst.stateZ0Z_28 ));
    LocalMux I__4034 (
            .O(N__22122),
            .I(\b2v_inst.stateZ0Z_28 ));
    InMux I__4033 (
            .O(N__22109),
            .I(N__22097));
    InMux I__4032 (
            .O(N__22108),
            .I(N__22097));
    InMux I__4031 (
            .O(N__22107),
            .I(N__22097));
    InMux I__4030 (
            .O(N__22106),
            .I(N__22097));
    LocalMux I__4029 (
            .O(N__22097),
            .I(N__22092));
    InMux I__4028 (
            .O(N__22096),
            .I(N__22089));
    InMux I__4027 (
            .O(N__22095),
            .I(N__22082));
    Sp12to4 I__4026 (
            .O(N__22092),
            .I(N__22077));
    LocalMux I__4025 (
            .O(N__22089),
            .I(N__22077));
    InMux I__4024 (
            .O(N__22088),
            .I(N__22070));
    InMux I__4023 (
            .O(N__22087),
            .I(N__22070));
    InMux I__4022 (
            .O(N__22086),
            .I(N__22070));
    InMux I__4021 (
            .O(N__22085),
            .I(N__22067));
    LocalMux I__4020 (
            .O(N__22082),
            .I(\b2v_inst.N_432_1 ));
    Odrv12 I__4019 (
            .O(N__22077),
            .I(\b2v_inst.N_432_1 ));
    LocalMux I__4018 (
            .O(N__22070),
            .I(\b2v_inst.N_432_1 ));
    LocalMux I__4017 (
            .O(N__22067),
            .I(\b2v_inst.N_432_1 ));
    CEMux I__4016 (
            .O(N__22058),
            .I(N__22053));
    CEMux I__4015 (
            .O(N__22057),
            .I(N__22050));
    CEMux I__4014 (
            .O(N__22056),
            .I(N__22047));
    LocalMux I__4013 (
            .O(N__22053),
            .I(N__22043));
    LocalMux I__4012 (
            .O(N__22050),
            .I(N__22040));
    LocalMux I__4011 (
            .O(N__22047),
            .I(N__22037));
    CEMux I__4010 (
            .O(N__22046),
            .I(N__22034));
    Span4Mux_h I__4009 (
            .O(N__22043),
            .I(N__22030));
    Span4Mux_h I__4008 (
            .O(N__22040),
            .I(N__22027));
    Span4Mux_h I__4007 (
            .O(N__22037),
            .I(N__22022));
    LocalMux I__4006 (
            .O(N__22034),
            .I(N__22022));
    CEMux I__4005 (
            .O(N__22033),
            .I(N__22019));
    Span4Mux_h I__4004 (
            .O(N__22030),
            .I(N__22016));
    Span4Mux_h I__4003 (
            .O(N__22027),
            .I(N__22011));
    Span4Mux_h I__4002 (
            .O(N__22022),
            .I(N__22011));
    LocalMux I__4001 (
            .O(N__22019),
            .I(N__22008));
    Odrv4 I__4000 (
            .O(N__22016),
            .I(\b2v_inst.N_442_i ));
    Odrv4 I__3999 (
            .O(N__22011),
            .I(\b2v_inst.N_442_i ));
    Odrv4 I__3998 (
            .O(N__22008),
            .I(\b2v_inst.N_442_i ));
    CascadeMux I__3997 (
            .O(N__22001),
            .I(N__21998));
    InMux I__3996 (
            .O(N__21998),
            .I(N__21995));
    LocalMux I__3995 (
            .O(N__21995),
            .I(N__21992));
    Span4Mux_h I__3994 (
            .O(N__21992),
            .I(N__21989));
    Odrv4 I__3993 (
            .O(N__21989),
            .I(\b2v_inst.un2_dir_mem_2_cry_0_THRU_CO ));
    InMux I__3992 (
            .O(N__21986),
            .I(\b2v_inst.un2_dir_mem_2_cry_0 ));
    CascadeMux I__3991 (
            .O(N__21983),
            .I(N__21980));
    InMux I__3990 (
            .O(N__21980),
            .I(N__21977));
    LocalMux I__3989 (
            .O(N__21977),
            .I(N__21974));
    Span4Mux_h I__3988 (
            .O(N__21974),
            .I(N__21971));
    Odrv4 I__3987 (
            .O(N__21971),
            .I(\b2v_inst.dir_mem_2_RNO_0Z0Z_2 ));
    InMux I__3986 (
            .O(N__21968),
            .I(\b2v_inst.un2_dir_mem_2_cry_1 ));
    CascadeMux I__3985 (
            .O(N__21965),
            .I(N__21962));
    InMux I__3984 (
            .O(N__21962),
            .I(N__21959));
    LocalMux I__3983 (
            .O(N__21959),
            .I(N__21956));
    Odrv4 I__3982 (
            .O(N__21956),
            .I(\b2v_inst.dir_mem_2_RNO_0Z0Z_3 ));
    InMux I__3981 (
            .O(N__21953),
            .I(\b2v_inst.un2_dir_mem_2_cry_2 ));
    CascadeMux I__3980 (
            .O(N__21950),
            .I(N__21947));
    InMux I__3979 (
            .O(N__21947),
            .I(N__21944));
    LocalMux I__3978 (
            .O(N__21944),
            .I(N__21941));
    Odrv4 I__3977 (
            .O(N__21941),
            .I(\b2v_inst.dir_mem_2_RNO_0Z0Z_4 ));
    InMux I__3976 (
            .O(N__21938),
            .I(\b2v_inst.un2_dir_mem_2_cry_3 ));
    InMux I__3975 (
            .O(N__21935),
            .I(N__21932));
    LocalMux I__3974 (
            .O(N__21932),
            .I(N__21928));
    InMux I__3973 (
            .O(N__21931),
            .I(N__21925));
    Span4Mux_v I__3972 (
            .O(N__21928),
            .I(N__21920));
    LocalMux I__3971 (
            .O(N__21925),
            .I(N__21920));
    Odrv4 I__3970 (
            .O(N__21920),
            .I(\b2v_inst.state_ns_0_i_o2_8_23 ));
    InMux I__3969 (
            .O(N__21917),
            .I(N__21914));
    LocalMux I__3968 (
            .O(N__21914),
            .I(N__21911));
    Span4Mux_h I__3967 (
            .O(N__21911),
            .I(N__21908));
    Span4Mux_v I__3966 (
            .O(N__21908),
            .I(N__21905));
    Span4Mux_h I__3965 (
            .O(N__21905),
            .I(N__21902));
    Odrv4 I__3964 (
            .O(N__21902),
            .I(N_550_i));
    InMux I__3963 (
            .O(N__21899),
            .I(N__21896));
    LocalMux I__3962 (
            .O(N__21896),
            .I(\b2v_inst.state_fastZ0Z_32 ));
    InMux I__3961 (
            .O(N__21893),
            .I(N__21883));
    InMux I__3960 (
            .O(N__21892),
            .I(N__21883));
    CascadeMux I__3959 (
            .O(N__21891),
            .I(N__21879));
    InMux I__3958 (
            .O(N__21890),
            .I(N__21871));
    InMux I__3957 (
            .O(N__21889),
            .I(N__21871));
    InMux I__3956 (
            .O(N__21888),
            .I(N__21871));
    LocalMux I__3955 (
            .O(N__21883),
            .I(N__21868));
    InMux I__3954 (
            .O(N__21882),
            .I(N__21865));
    InMux I__3953 (
            .O(N__21879),
            .I(N__21860));
    InMux I__3952 (
            .O(N__21878),
            .I(N__21857));
    LocalMux I__3951 (
            .O(N__21871),
            .I(N__21854));
    Span4Mux_h I__3950 (
            .O(N__21868),
            .I(N__21851));
    LocalMux I__3949 (
            .O(N__21865),
            .I(N__21848));
    InMux I__3948 (
            .O(N__21864),
            .I(N__21845));
    InMux I__3947 (
            .O(N__21863),
            .I(N__21842));
    LocalMux I__3946 (
            .O(N__21860),
            .I(\b2v_inst.stateZ0Z_5 ));
    LocalMux I__3945 (
            .O(N__21857),
            .I(\b2v_inst.stateZ0Z_5 ));
    Odrv4 I__3944 (
            .O(N__21854),
            .I(\b2v_inst.stateZ0Z_5 ));
    Odrv4 I__3943 (
            .O(N__21851),
            .I(\b2v_inst.stateZ0Z_5 ));
    Odrv12 I__3942 (
            .O(N__21848),
            .I(\b2v_inst.stateZ0Z_5 ));
    LocalMux I__3941 (
            .O(N__21845),
            .I(\b2v_inst.stateZ0Z_5 ));
    LocalMux I__3940 (
            .O(N__21842),
            .I(\b2v_inst.stateZ0Z_5 ));
    InMux I__3939 (
            .O(N__21827),
            .I(N__21824));
    LocalMux I__3938 (
            .O(N__21824),
            .I(\b2v_inst.addr_ram_energia_ss0_0_i_o2_i_o2_0 ));
    InMux I__3937 (
            .O(N__21821),
            .I(N__21818));
    LocalMux I__3936 (
            .O(N__21818),
            .I(N__21815));
    Span12Mux_h I__3935 (
            .O(N__21815),
            .I(N__21812));
    Odrv12 I__3934 (
            .O(N__21812),
            .I(\b2v_inst.dir_mem_RNO_0Z0Z_6 ));
    InMux I__3933 (
            .O(N__21809),
            .I(N__21806));
    LocalMux I__3932 (
            .O(N__21806),
            .I(N__21803));
    Span4Mux_h I__3931 (
            .O(N__21803),
            .I(N__21800));
    Span4Mux_v I__3930 (
            .O(N__21800),
            .I(N__21797));
    Odrv4 I__3929 (
            .O(N__21797),
            .I(\b2v_inst.dir_memZ0Z_6 ));
    InMux I__3928 (
            .O(N__21794),
            .I(N__21791));
    LocalMux I__3927 (
            .O(N__21791),
            .I(N__21788));
    Span4Mux_v I__3926 (
            .O(N__21788),
            .I(N__21785));
    Span4Mux_h I__3925 (
            .O(N__21785),
            .I(N__21782));
    Odrv4 I__3924 (
            .O(N__21782),
            .I(\b2v_inst.dir_mem_RNO_0Z0Z_8 ));
    InMux I__3923 (
            .O(N__21779),
            .I(N__21776));
    LocalMux I__3922 (
            .O(N__21776),
            .I(N__21773));
    Span4Mux_v I__3921 (
            .O(N__21773),
            .I(N__21770));
    Span4Mux_v I__3920 (
            .O(N__21770),
            .I(N__21767));
    Odrv4 I__3919 (
            .O(N__21767),
            .I(\b2v_inst.dir_memZ0Z_8 ));
    CascadeMux I__3918 (
            .O(N__21764),
            .I(N__21761));
    InMux I__3917 (
            .O(N__21761),
            .I(N__21758));
    LocalMux I__3916 (
            .O(N__21758),
            .I(N__21755));
    Span4Mux_v I__3915 (
            .O(N__21755),
            .I(N__21752));
    Span4Mux_h I__3914 (
            .O(N__21752),
            .I(N__21749));
    Odrv4 I__3913 (
            .O(N__21749),
            .I(\b2v_inst.dir_mem_RNO_0Z0Z_9 ));
    InMux I__3912 (
            .O(N__21746),
            .I(N__21743));
    LocalMux I__3911 (
            .O(N__21743),
            .I(N__21740));
    Odrv12 I__3910 (
            .O(N__21740),
            .I(\b2v_inst.dir_memZ0Z_9 ));
    InMux I__3909 (
            .O(N__21737),
            .I(N__21734));
    LocalMux I__3908 (
            .O(N__21734),
            .I(N__21731));
    Span4Mux_v I__3907 (
            .O(N__21731),
            .I(N__21728));
    Sp12to4 I__3906 (
            .O(N__21728),
            .I(N__21725));
    Span12Mux_h I__3905 (
            .O(N__21725),
            .I(N__21722));
    Odrv12 I__3904 (
            .O(N__21722),
            .I(swit_c_4));
    InMux I__3903 (
            .O(N__21719),
            .I(N__21714));
    InMux I__3902 (
            .O(N__21718),
            .I(N__21711));
    InMux I__3901 (
            .O(N__21717),
            .I(N__21701));
    LocalMux I__3900 (
            .O(N__21714),
            .I(N__21698));
    LocalMux I__3899 (
            .O(N__21711),
            .I(N__21695));
    InMux I__3898 (
            .O(N__21710),
            .I(N__21692));
    InMux I__3897 (
            .O(N__21709),
            .I(N__21687));
    InMux I__3896 (
            .O(N__21708),
            .I(N__21687));
    InMux I__3895 (
            .O(N__21707),
            .I(N__21678));
    InMux I__3894 (
            .O(N__21706),
            .I(N__21678));
    InMux I__3893 (
            .O(N__21705),
            .I(N__21678));
    InMux I__3892 (
            .O(N__21704),
            .I(N__21678));
    LocalMux I__3891 (
            .O(N__21701),
            .I(\b2v_inst.N_494 ));
    Odrv12 I__3890 (
            .O(N__21698),
            .I(\b2v_inst.N_494 ));
    Odrv4 I__3889 (
            .O(N__21695),
            .I(\b2v_inst.N_494 ));
    LocalMux I__3888 (
            .O(N__21692),
            .I(\b2v_inst.N_494 ));
    LocalMux I__3887 (
            .O(N__21687),
            .I(\b2v_inst.N_494 ));
    LocalMux I__3886 (
            .O(N__21678),
            .I(\b2v_inst.N_494 ));
    InMux I__3885 (
            .O(N__21665),
            .I(N__21655));
    InMux I__3884 (
            .O(N__21664),
            .I(N__21655));
    InMux I__3883 (
            .O(N__21663),
            .I(N__21655));
    InMux I__3882 (
            .O(N__21662),
            .I(N__21651));
    LocalMux I__3881 (
            .O(N__21655),
            .I(N__21648));
    InMux I__3880 (
            .O(N__21654),
            .I(N__21645));
    LocalMux I__3879 (
            .O(N__21651),
            .I(N__21642));
    Span4Mux_h I__3878 (
            .O(N__21648),
            .I(N__21637));
    LocalMux I__3877 (
            .O(N__21645),
            .I(N__21637));
    Span12Mux_h I__3876 (
            .O(N__21642),
            .I(N__21628));
    Span4Mux_v I__3875 (
            .O(N__21637),
            .I(N__21625));
    InMux I__3874 (
            .O(N__21636),
            .I(N__21622));
    InMux I__3873 (
            .O(N__21635),
            .I(N__21619));
    InMux I__3872 (
            .O(N__21634),
            .I(N__21610));
    InMux I__3871 (
            .O(N__21633),
            .I(N__21610));
    InMux I__3870 (
            .O(N__21632),
            .I(N__21610));
    InMux I__3869 (
            .O(N__21631),
            .I(N__21610));
    Odrv12 I__3868 (
            .O(N__21628),
            .I(\b2v_inst.N_247 ));
    Odrv4 I__3867 (
            .O(N__21625),
            .I(\b2v_inst.N_247 ));
    LocalMux I__3866 (
            .O(N__21622),
            .I(\b2v_inst.N_247 ));
    LocalMux I__3865 (
            .O(N__21619),
            .I(\b2v_inst.N_247 ));
    LocalMux I__3864 (
            .O(N__21610),
            .I(\b2v_inst.N_247 ));
    CascadeMux I__3863 (
            .O(N__21599),
            .I(\b2v_inst.addr_ram_energia_m0_4_cascade_ ));
    CascadeMux I__3862 (
            .O(N__21596),
            .I(N__21592));
    CascadeMux I__3861 (
            .O(N__21595),
            .I(N__21589));
    CascadeBuf I__3860 (
            .O(N__21592),
            .I(N__21586));
    CascadeBuf I__3859 (
            .O(N__21589),
            .I(N__21583));
    CascadeMux I__3858 (
            .O(N__21586),
            .I(N__21580));
    CascadeMux I__3857 (
            .O(N__21583),
            .I(N__21577));
    CascadeBuf I__3856 (
            .O(N__21580),
            .I(N__21574));
    CascadeBuf I__3855 (
            .O(N__21577),
            .I(N__21571));
    CascadeMux I__3854 (
            .O(N__21574),
            .I(N__21568));
    CascadeMux I__3853 (
            .O(N__21571),
            .I(N__21565));
    CascadeBuf I__3852 (
            .O(N__21568),
            .I(N__21562));
    CascadeBuf I__3851 (
            .O(N__21565),
            .I(N__21559));
    CascadeMux I__3850 (
            .O(N__21562),
            .I(N__21556));
    CascadeMux I__3849 (
            .O(N__21559),
            .I(N__21553));
    CascadeBuf I__3848 (
            .O(N__21556),
            .I(N__21550));
    CascadeBuf I__3847 (
            .O(N__21553),
            .I(N__21547));
    CascadeMux I__3846 (
            .O(N__21550),
            .I(N__21544));
    CascadeMux I__3845 (
            .O(N__21547),
            .I(N__21541));
    CascadeBuf I__3844 (
            .O(N__21544),
            .I(N__21538));
    CascadeBuf I__3843 (
            .O(N__21541),
            .I(N__21535));
    CascadeMux I__3842 (
            .O(N__21538),
            .I(N__21532));
    CascadeMux I__3841 (
            .O(N__21535),
            .I(N__21529));
    CascadeBuf I__3840 (
            .O(N__21532),
            .I(N__21526));
    CascadeBuf I__3839 (
            .O(N__21529),
            .I(N__21523));
    CascadeMux I__3838 (
            .O(N__21526),
            .I(N__21520));
    CascadeMux I__3837 (
            .O(N__21523),
            .I(N__21517));
    InMux I__3836 (
            .O(N__21520),
            .I(N__21514));
    InMux I__3835 (
            .O(N__21517),
            .I(N__21511));
    LocalMux I__3834 (
            .O(N__21514),
            .I(N__21506));
    LocalMux I__3833 (
            .O(N__21511),
            .I(N__21506));
    Span4Mux_v I__3832 (
            .O(N__21506),
            .I(N__21503));
    Span4Mux_h I__3831 (
            .O(N__21503),
            .I(N__21500));
    Span4Mux_h I__3830 (
            .O(N__21500),
            .I(N__21497));
    Odrv4 I__3829 (
            .O(N__21497),
            .I(SYNTHESIZED_WIRE_12_4));
    InMux I__3828 (
            .O(N__21494),
            .I(N__21491));
    LocalMux I__3827 (
            .O(N__21491),
            .I(N__21488));
    Span4Mux_h I__3826 (
            .O(N__21488),
            .I(N__21485));
    Span4Mux_v I__3825 (
            .O(N__21485),
            .I(N__21482));
    Span4Mux_v I__3824 (
            .O(N__21482),
            .I(N__21479));
    Odrv4 I__3823 (
            .O(N__21479),
            .I(uart_rx_i_c));
    CascadeMux I__3822 (
            .O(N__21476),
            .I(\b2v_inst.state18_li_0_cascade_ ));
    CEMux I__3821 (
            .O(N__21473),
            .I(N__21470));
    LocalMux I__3820 (
            .O(N__21470),
            .I(N__21464));
    CEMux I__3819 (
            .O(N__21469),
            .I(N__21461));
    CEMux I__3818 (
            .O(N__21468),
            .I(N__21458));
    CEMux I__3817 (
            .O(N__21467),
            .I(N__21450));
    Span4Mux_v I__3816 (
            .O(N__21464),
            .I(N__21440));
    LocalMux I__3815 (
            .O(N__21461),
            .I(N__21440));
    LocalMux I__3814 (
            .O(N__21458),
            .I(N__21440));
    CEMux I__3813 (
            .O(N__21457),
            .I(N__21437));
    CEMux I__3812 (
            .O(N__21456),
            .I(N__21434));
    CEMux I__3811 (
            .O(N__21455),
            .I(N__21431));
    CEMux I__3810 (
            .O(N__21454),
            .I(N__21428));
    CEMux I__3809 (
            .O(N__21453),
            .I(N__21423));
    LocalMux I__3808 (
            .O(N__21450),
            .I(N__21420));
    CEMux I__3807 (
            .O(N__21449),
            .I(N__21417));
    CEMux I__3806 (
            .O(N__21448),
            .I(N__21414));
    CEMux I__3805 (
            .O(N__21447),
            .I(N__21411));
    Span4Mux_v I__3804 (
            .O(N__21440),
            .I(N__21403));
    LocalMux I__3803 (
            .O(N__21437),
            .I(N__21403));
    LocalMux I__3802 (
            .O(N__21434),
            .I(N__21403));
    LocalMux I__3801 (
            .O(N__21431),
            .I(N__21398));
    LocalMux I__3800 (
            .O(N__21428),
            .I(N__21398));
    CEMux I__3799 (
            .O(N__21427),
            .I(N__21395));
    CEMux I__3798 (
            .O(N__21426),
            .I(N__21392));
    LocalMux I__3797 (
            .O(N__21423),
            .I(N__21388));
    Span4Mux_v I__3796 (
            .O(N__21420),
            .I(N__21381));
    LocalMux I__3795 (
            .O(N__21417),
            .I(N__21381));
    LocalMux I__3794 (
            .O(N__21414),
            .I(N__21381));
    LocalMux I__3793 (
            .O(N__21411),
            .I(N__21378));
    CEMux I__3792 (
            .O(N__21410),
            .I(N__21375));
    Span4Mux_v I__3791 (
            .O(N__21403),
            .I(N__21368));
    Span4Mux_v I__3790 (
            .O(N__21398),
            .I(N__21368));
    LocalMux I__3789 (
            .O(N__21395),
            .I(N__21368));
    LocalMux I__3788 (
            .O(N__21392),
            .I(N__21365));
    CEMux I__3787 (
            .O(N__21391),
            .I(N__21362));
    Span4Mux_h I__3786 (
            .O(N__21388),
            .I(N__21359));
    Span4Mux_v I__3785 (
            .O(N__21381),
            .I(N__21352));
    Span4Mux_v I__3784 (
            .O(N__21378),
            .I(N__21352));
    LocalMux I__3783 (
            .O(N__21375),
            .I(N__21352));
    Span4Mux_v I__3782 (
            .O(N__21368),
            .I(N__21349));
    Span4Mux_v I__3781 (
            .O(N__21365),
            .I(N__21344));
    LocalMux I__3780 (
            .O(N__21362),
            .I(N__21344));
    Span4Mux_h I__3779 (
            .O(N__21359),
            .I(N__21341));
    Span4Mux_h I__3778 (
            .O(N__21352),
            .I(N__21338));
    Span4Mux_h I__3777 (
            .O(N__21349),
            .I(N__21335));
    Span4Mux_h I__3776 (
            .O(N__21344),
            .I(N__21332));
    Span4Mux_v I__3775 (
            .O(N__21341),
            .I(N__21327));
    Span4Mux_h I__3774 (
            .O(N__21338),
            .I(N__21327));
    Span4Mux_h I__3773 (
            .O(N__21335),
            .I(N__21324));
    Span4Mux_h I__3772 (
            .O(N__21332),
            .I(N__21319));
    Span4Mux_h I__3771 (
            .O(N__21327),
            .I(N__21319));
    Odrv4 I__3770 (
            .O(N__21324),
            .I(N_130_i));
    Odrv4 I__3769 (
            .O(N__21319),
            .I(N_130_i));
    InMux I__3768 (
            .O(N__21314),
            .I(N__21309));
    InMux I__3767 (
            .O(N__21313),
            .I(N__21304));
    InMux I__3766 (
            .O(N__21312),
            .I(N__21304));
    LocalMux I__3765 (
            .O(N__21309),
            .I(N__21299));
    LocalMux I__3764 (
            .O(N__21304),
            .I(N__21296));
    CascadeMux I__3763 (
            .O(N__21303),
            .I(N__21293));
    CascadeMux I__3762 (
            .O(N__21302),
            .I(N__21290));
    Span4Mux_h I__3761 (
            .O(N__21299),
            .I(N__21287));
    Span4Mux_h I__3760 (
            .O(N__21296),
            .I(N__21284));
    InMux I__3759 (
            .O(N__21293),
            .I(N__21281));
    InMux I__3758 (
            .O(N__21290),
            .I(N__21278));
    Odrv4 I__3757 (
            .O(N__21287),
            .I(\b2v_inst.N_512 ));
    Odrv4 I__3756 (
            .O(N__21284),
            .I(\b2v_inst.N_512 ));
    LocalMux I__3755 (
            .O(N__21281),
            .I(\b2v_inst.N_512 ));
    LocalMux I__3754 (
            .O(N__21278),
            .I(\b2v_inst.N_512 ));
    InMux I__3753 (
            .O(N__21269),
            .I(N__21266));
    LocalMux I__3752 (
            .O(N__21266),
            .I(N__21262));
    CascadeMux I__3751 (
            .O(N__21265),
            .I(N__21259));
    Span4Mux_v I__3750 (
            .O(N__21262),
            .I(N__21255));
    InMux I__3749 (
            .O(N__21259),
            .I(N__21244));
    InMux I__3748 (
            .O(N__21258),
            .I(N__21244));
    Span4Mux_h I__3747 (
            .O(N__21255),
            .I(N__21241));
    InMux I__3746 (
            .O(N__21254),
            .I(N__21236));
    InMux I__3745 (
            .O(N__21253),
            .I(N__21236));
    InMux I__3744 (
            .O(N__21252),
            .I(N__21229));
    InMux I__3743 (
            .O(N__21251),
            .I(N__21229));
    InMux I__3742 (
            .O(N__21250),
            .I(N__21229));
    InMux I__3741 (
            .O(N__21249),
            .I(N__21226));
    LocalMux I__3740 (
            .O(N__21244),
            .I(N__21223));
    Span4Mux_h I__3739 (
            .O(N__21241),
            .I(N__21218));
    LocalMux I__3738 (
            .O(N__21236),
            .I(N__21218));
    LocalMux I__3737 (
            .O(N__21229),
            .I(\b2v_inst.stateZ0Z_30 ));
    LocalMux I__3736 (
            .O(N__21226),
            .I(\b2v_inst.stateZ0Z_30 ));
    Odrv4 I__3735 (
            .O(N__21223),
            .I(\b2v_inst.stateZ0Z_30 ));
    Odrv4 I__3734 (
            .O(N__21218),
            .I(\b2v_inst.stateZ0Z_30 ));
    CascadeMux I__3733 (
            .O(N__21209),
            .I(\b2v_inst.N_828_cascade_ ));
    InMux I__3732 (
            .O(N__21206),
            .I(N__21203));
    LocalMux I__3731 (
            .O(N__21203),
            .I(N__21200));
    Span4Mux_h I__3730 (
            .O(N__21200),
            .I(N__21197));
    Span4Mux_h I__3729 (
            .O(N__21197),
            .I(N__21194));
    Odrv4 I__3728 (
            .O(N__21194),
            .I(N_552_i));
    InMux I__3727 (
            .O(N__21191),
            .I(N__21185));
    InMux I__3726 (
            .O(N__21190),
            .I(N__21185));
    LocalMux I__3725 (
            .O(N__21185),
            .I(N__21182));
    Span4Mux_h I__3724 (
            .O(N__21182),
            .I(N__21178));
    InMux I__3723 (
            .O(N__21181),
            .I(N__21175));
    Odrv4 I__3722 (
            .O(N__21178),
            .I(\b2v_inst1.N_119 ));
    LocalMux I__3721 (
            .O(N__21175),
            .I(\b2v_inst1.N_119 ));
    CascadeMux I__3720 (
            .O(N__21170),
            .I(\b2v_inst1.r_Clk_Count_6_iv_0_a3_1_1_1_cascade_ ));
    InMux I__3719 (
            .O(N__21167),
            .I(N__21160));
    InMux I__3718 (
            .O(N__21166),
            .I(N__21160));
    InMux I__3717 (
            .O(N__21165),
            .I(N__21157));
    LocalMux I__3716 (
            .O(N__21160),
            .I(N__21154));
    LocalMux I__3715 (
            .O(N__21157),
            .I(N__21151));
    Span4Mux_v I__3714 (
            .O(N__21154),
            .I(N__21147));
    Span4Mux_h I__3713 (
            .O(N__21151),
            .I(N__21142));
    InMux I__3712 (
            .O(N__21150),
            .I(N__21139));
    Span4Mux_h I__3711 (
            .O(N__21147),
            .I(N__21136));
    InMux I__3710 (
            .O(N__21146),
            .I(N__21131));
    InMux I__3709 (
            .O(N__21145),
            .I(N__21131));
    Odrv4 I__3708 (
            .O(N__21142),
            .I(\b2v_inst1.N_43 ));
    LocalMux I__3707 (
            .O(N__21139),
            .I(\b2v_inst1.N_43 ));
    Odrv4 I__3706 (
            .O(N__21136),
            .I(\b2v_inst1.N_43 ));
    LocalMux I__3705 (
            .O(N__21131),
            .I(\b2v_inst1.N_43 ));
    CascadeMux I__3704 (
            .O(N__21122),
            .I(\b2v_inst1.r_Clk_Count_6_iv_0_0_1_cascade_ ));
    InMux I__3703 (
            .O(N__21119),
            .I(N__21116));
    LocalMux I__3702 (
            .O(N__21116),
            .I(N__21113));
    Span4Mux_h I__3701 (
            .O(N__21113),
            .I(N__21105));
    InMux I__3700 (
            .O(N__21112),
            .I(N__21102));
    InMux I__3699 (
            .O(N__21111),
            .I(N__21097));
    InMux I__3698 (
            .O(N__21110),
            .I(N__21097));
    InMux I__3697 (
            .O(N__21109),
            .I(N__21092));
    InMux I__3696 (
            .O(N__21108),
            .I(N__21092));
    Odrv4 I__3695 (
            .O(N__21105),
            .I(\b2v_inst1.r_Clk_CountZ0Z_0 ));
    LocalMux I__3694 (
            .O(N__21102),
            .I(\b2v_inst1.r_Clk_CountZ0Z_0 ));
    LocalMux I__3693 (
            .O(N__21097),
            .I(\b2v_inst1.r_Clk_CountZ0Z_0 ));
    LocalMux I__3692 (
            .O(N__21092),
            .I(\b2v_inst1.r_Clk_CountZ0Z_0 ));
    CascadeMux I__3691 (
            .O(N__21083),
            .I(N__21079));
    InMux I__3690 (
            .O(N__21082),
            .I(N__21073));
    InMux I__3689 (
            .O(N__21079),
            .I(N__21068));
    InMux I__3688 (
            .O(N__21078),
            .I(N__21068));
    InMux I__3687 (
            .O(N__21077),
            .I(N__21064));
    CascadeMux I__3686 (
            .O(N__21076),
            .I(N__21061));
    LocalMux I__3685 (
            .O(N__21073),
            .I(N__21058));
    LocalMux I__3684 (
            .O(N__21068),
            .I(N__21055));
    InMux I__3683 (
            .O(N__21067),
            .I(N__21052));
    LocalMux I__3682 (
            .O(N__21064),
            .I(N__21049));
    InMux I__3681 (
            .O(N__21061),
            .I(N__21046));
    Span4Mux_h I__3680 (
            .O(N__21058),
            .I(N__21043));
    Span4Mux_h I__3679 (
            .O(N__21055),
            .I(N__21040));
    LocalMux I__3678 (
            .O(N__21052),
            .I(N__21035));
    Span4Mux_h I__3677 (
            .O(N__21049),
            .I(N__21035));
    LocalMux I__3676 (
            .O(N__21046),
            .I(\b2v_inst1.r_Clk_CountZ0Z_1 ));
    Odrv4 I__3675 (
            .O(N__21043),
            .I(\b2v_inst1.r_Clk_CountZ0Z_1 ));
    Odrv4 I__3674 (
            .O(N__21040),
            .I(\b2v_inst1.r_Clk_CountZ0Z_1 ));
    Odrv4 I__3673 (
            .O(N__21035),
            .I(\b2v_inst1.r_Clk_CountZ0Z_1 ));
    CascadeMux I__3672 (
            .O(N__21026),
            .I(\b2v_inst.N_653_cascade_ ));
    CascadeMux I__3671 (
            .O(N__21023),
            .I(N__21019));
    InMux I__3670 (
            .O(N__21022),
            .I(N__21011));
    InMux I__3669 (
            .O(N__21019),
            .I(N__21011));
    InMux I__3668 (
            .O(N__21018),
            .I(N__21011));
    LocalMux I__3667 (
            .O(N__21011),
            .I(\b2v_inst.stateZ0Z_17 ));
    InMux I__3666 (
            .O(N__21008),
            .I(N__21005));
    LocalMux I__3665 (
            .O(N__21005),
            .I(\b2v_inst.state_ns_i_a2_1_15 ));
    CascadeMux I__3664 (
            .O(N__21002),
            .I(\b2v_inst.cuenta_RNIKUJVZ0Z_0_cascade_ ));
    CascadeMux I__3663 (
            .O(N__20999),
            .I(\b2v_inst.un20_cuentalto10_5_cascade_ ));
    InMux I__3662 (
            .O(N__20996),
            .I(N__20993));
    LocalMux I__3661 (
            .O(N__20993),
            .I(\b2v_inst.un20_cuentalto10_sx ));
    CascadeMux I__3660 (
            .O(N__20990),
            .I(\b2v_inst.un20_cuentalto10_sx_cascade_ ));
    InMux I__3659 (
            .O(N__20987),
            .I(N__20983));
    InMux I__3658 (
            .O(N__20986),
            .I(N__20980));
    LocalMux I__3657 (
            .O(N__20983),
            .I(\b2v_inst.N_829 ));
    LocalMux I__3656 (
            .O(N__20980),
            .I(\b2v_inst.N_829 ));
    CascadeMux I__3655 (
            .O(N__20975),
            .I(\b2v_inst.un1_state_23_i_a2_0_a2_0_a2_0_cascade_ ));
    InMux I__3654 (
            .O(N__20972),
            .I(N__20969));
    LocalMux I__3653 (
            .O(N__20969),
            .I(N__20965));
    InMux I__3652 (
            .O(N__20968),
            .I(N__20961));
    Span4Mux_h I__3651 (
            .O(N__20965),
            .I(N__20958));
    InMux I__3650 (
            .O(N__20964),
            .I(N__20955));
    LocalMux I__3649 (
            .O(N__20961),
            .I(\b2v_inst.stateZ0Z_22 ));
    Odrv4 I__3648 (
            .O(N__20958),
            .I(\b2v_inst.stateZ0Z_22 ));
    LocalMux I__3647 (
            .O(N__20955),
            .I(\b2v_inst.stateZ0Z_22 ));
    InMux I__3646 (
            .O(N__20948),
            .I(N__20943));
    InMux I__3645 (
            .O(N__20947),
            .I(N__20939));
    InMux I__3644 (
            .O(N__20946),
            .I(N__20936));
    LocalMux I__3643 (
            .O(N__20943),
            .I(N__20933));
    InMux I__3642 (
            .O(N__20942),
            .I(N__20930));
    LocalMux I__3641 (
            .O(N__20939),
            .I(N__20927));
    LocalMux I__3640 (
            .O(N__20936),
            .I(\b2v_inst.stateZ0Z_26 ));
    Odrv4 I__3639 (
            .O(N__20933),
            .I(\b2v_inst.stateZ0Z_26 ));
    LocalMux I__3638 (
            .O(N__20930),
            .I(\b2v_inst.stateZ0Z_26 ));
    Odrv4 I__3637 (
            .O(N__20927),
            .I(\b2v_inst.stateZ0Z_26 ));
    InMux I__3636 (
            .O(N__20918),
            .I(N__20915));
    LocalMux I__3635 (
            .O(N__20915),
            .I(\b2v_inst.un2_cuentalto10_i_a2_6 ));
    InMux I__3634 (
            .O(N__20912),
            .I(N__20909));
    LocalMux I__3633 (
            .O(N__20909),
            .I(N__20906));
    Span4Mux_v I__3632 (
            .O(N__20906),
            .I(N__20903));
    Span4Mux_h I__3631 (
            .O(N__20903),
            .I(N__20899));
    InMux I__3630 (
            .O(N__20902),
            .I(N__20896));
    Odrv4 I__3629 (
            .O(N__20899),
            .I(\b2v_inst1.m16_0_o2 ));
    LocalMux I__3628 (
            .O(N__20896),
            .I(\b2v_inst1.m16_0_o2 ));
    CascadeMux I__3627 (
            .O(N__20891),
            .I(\b2v_inst1.m16_0_a3_0_cascade_ ));
    InMux I__3626 (
            .O(N__20888),
            .I(N__20885));
    LocalMux I__3625 (
            .O(N__20885),
            .I(N__20882));
    Span4Mux_h I__3624 (
            .O(N__20882),
            .I(N__20879));
    Odrv4 I__3623 (
            .O(N__20879),
            .I(\b2v_inst.dir_mem_1Z0Z_9 ));
    CascadeMux I__3622 (
            .O(N__20876),
            .I(N__20873));
    InMux I__3621 (
            .O(N__20873),
            .I(N__20870));
    LocalMux I__3620 (
            .O(N__20870),
            .I(N__20867));
    Span4Mux_v I__3619 (
            .O(N__20867),
            .I(N__20864));
    Span4Mux_h I__3618 (
            .O(N__20864),
            .I(N__20861));
    Odrv4 I__3617 (
            .O(N__20861),
            .I(\b2v_inst.dir_mem_3Z0Z_9 ));
    InMux I__3616 (
            .O(N__20858),
            .I(N__20855));
    LocalMux I__3615 (
            .O(N__20855),
            .I(N__20852));
    Span4Mux_h I__3614 (
            .O(N__20852),
            .I(N__20849));
    Span4Mux_h I__3613 (
            .O(N__20849),
            .I(N__20846));
    Odrv4 I__3612 (
            .O(N__20846),
            .I(N_554_i));
    InMux I__3611 (
            .O(N__20843),
            .I(N__20840));
    LocalMux I__3610 (
            .O(N__20840),
            .I(N__20837));
    Span4Mux_v I__3609 (
            .O(N__20837),
            .I(N__20834));
    Span4Mux_h I__3608 (
            .O(N__20834),
            .I(N__20831));
    Odrv4 I__3607 (
            .O(N__20831),
            .I(\b2v_inst.dir_mem_2Z0Z_2 ));
    CascadeMux I__3606 (
            .O(N__20828),
            .I(N__20825));
    InMux I__3605 (
            .O(N__20825),
            .I(N__20822));
    LocalMux I__3604 (
            .O(N__20822),
            .I(N__20819));
    Odrv12 I__3603 (
            .O(N__20819),
            .I(\b2v_inst.dir_memZ0Z_2 ));
    CascadeMux I__3602 (
            .O(N__20816),
            .I(N__20813));
    InMux I__3601 (
            .O(N__20813),
            .I(N__20810));
    LocalMux I__3600 (
            .O(N__20810),
            .I(N__20807));
    Odrv4 I__3599 (
            .O(N__20807),
            .I(\b2v_inst.dir_mem_2Z0Z_9 ));
    InMux I__3598 (
            .O(N__20804),
            .I(N__20801));
    LocalMux I__3597 (
            .O(N__20801),
            .I(\b2v_inst.dir_mem_1Z0Z_2 ));
    CascadeMux I__3596 (
            .O(N__20798),
            .I(N__20795));
    InMux I__3595 (
            .O(N__20795),
            .I(N__20792));
    LocalMux I__3594 (
            .O(N__20792),
            .I(N__20789));
    Odrv12 I__3593 (
            .O(N__20789),
            .I(\b2v_inst.dir_mem_3Z0Z_2 ));
    CascadeMux I__3592 (
            .O(N__20786),
            .I(\b2v_inst.N_829_cascade_ ));
    InMux I__3591 (
            .O(N__20783),
            .I(N__20780));
    LocalMux I__3590 (
            .O(N__20780),
            .I(N__20776));
    CascadeMux I__3589 (
            .O(N__20779),
            .I(N__20773));
    Span4Mux_v I__3588 (
            .O(N__20776),
            .I(N__20770));
    InMux I__3587 (
            .O(N__20773),
            .I(N__20767));
    Span4Mux_h I__3586 (
            .O(N__20770),
            .I(N__20764));
    LocalMux I__3585 (
            .O(N__20767),
            .I(N__20761));
    Odrv4 I__3584 (
            .O(N__20764),
            .I(\b2v_inst.dir_mem_215lto7 ));
    Odrv4 I__3583 (
            .O(N__20761),
            .I(\b2v_inst.dir_mem_215lto7 ));
    InMux I__3582 (
            .O(N__20756),
            .I(N__20753));
    LocalMux I__3581 (
            .O(N__20753),
            .I(N__20750));
    Span4Mux_v I__3580 (
            .O(N__20750),
            .I(N__20747));
    Span4Mux_h I__3579 (
            .O(N__20747),
            .I(N__20744));
    Odrv4 I__3578 (
            .O(N__20744),
            .I(\b2v_inst.dir_mem_2Z0Z_7 ));
    InMux I__3577 (
            .O(N__20741),
            .I(N__20738));
    LocalMux I__3576 (
            .O(N__20738),
            .I(N__20735));
    Span4Mux_v I__3575 (
            .O(N__20735),
            .I(N__20731));
    InMux I__3574 (
            .O(N__20734),
            .I(N__20728));
    Odrv4 I__3573 (
            .O(N__20731),
            .I(\b2v_inst.un8_dir_mem_2_cry_6_c_RNIINQZ0Z5 ));
    LocalMux I__3572 (
            .O(N__20728),
            .I(\b2v_inst.un8_dir_mem_2_cry_6_c_RNIINQZ0Z5 ));
    CascadeMux I__3571 (
            .O(N__20723),
            .I(N__20720));
    InMux I__3570 (
            .O(N__20720),
            .I(N__20717));
    LocalMux I__3569 (
            .O(N__20717),
            .I(N__20714));
    Span4Mux_v I__3568 (
            .O(N__20714),
            .I(N__20711));
    Odrv4 I__3567 (
            .O(N__20711),
            .I(\b2v_inst.dir_mem_2Z0Z_8 ));
    InMux I__3566 (
            .O(N__20708),
            .I(N__20705));
    LocalMux I__3565 (
            .O(N__20705),
            .I(N__20702));
    Span4Mux_h I__3564 (
            .O(N__20702),
            .I(N__20698));
    InMux I__3563 (
            .O(N__20701),
            .I(N__20695));
    Odrv4 I__3562 (
            .O(N__20698),
            .I(\b2v_inst.un8_dir_mem_2_cry_7_c_RNIKQRZ0Z5 ));
    LocalMux I__3561 (
            .O(N__20695),
            .I(\b2v_inst.un8_dir_mem_2_cry_7_c_RNIKQRZ0Z5 ));
    CascadeMux I__3560 (
            .O(N__20690),
            .I(N__20686));
    InMux I__3559 (
            .O(N__20689),
            .I(N__20672));
    InMux I__3558 (
            .O(N__20686),
            .I(N__20672));
    InMux I__3557 (
            .O(N__20685),
            .I(N__20672));
    InMux I__3556 (
            .O(N__20684),
            .I(N__20659));
    InMux I__3555 (
            .O(N__20683),
            .I(N__20659));
    InMux I__3554 (
            .O(N__20682),
            .I(N__20659));
    InMux I__3553 (
            .O(N__20681),
            .I(N__20659));
    InMux I__3552 (
            .O(N__20680),
            .I(N__20659));
    InMux I__3551 (
            .O(N__20679),
            .I(N__20659));
    LocalMux I__3550 (
            .O(N__20672),
            .I(N__20656));
    LocalMux I__3549 (
            .O(N__20659),
            .I(N__20653));
    Odrv12 I__3548 (
            .O(N__20656),
            .I(\b2v_inst.dir_mem_215lto11_0 ));
    Odrv4 I__3547 (
            .O(N__20653),
            .I(\b2v_inst.dir_mem_215lto11_0 ));
    InMux I__3546 (
            .O(N__20648),
            .I(N__20627));
    InMux I__3545 (
            .O(N__20647),
            .I(N__20627));
    InMux I__3544 (
            .O(N__20646),
            .I(N__20627));
    InMux I__3543 (
            .O(N__20645),
            .I(N__20627));
    InMux I__3542 (
            .O(N__20644),
            .I(N__20627));
    InMux I__3541 (
            .O(N__20643),
            .I(N__20614));
    InMux I__3540 (
            .O(N__20642),
            .I(N__20614));
    InMux I__3539 (
            .O(N__20641),
            .I(N__20614));
    InMux I__3538 (
            .O(N__20640),
            .I(N__20614));
    InMux I__3537 (
            .O(N__20639),
            .I(N__20614));
    InMux I__3536 (
            .O(N__20638),
            .I(N__20614));
    LocalMux I__3535 (
            .O(N__20627),
            .I(N__20611));
    LocalMux I__3534 (
            .O(N__20614),
            .I(\b2v_inst.dir_mem_215lt11 ));
    Odrv4 I__3533 (
            .O(N__20611),
            .I(\b2v_inst.dir_mem_215lt11 ));
    CEMux I__3532 (
            .O(N__20606),
            .I(N__20603));
    LocalMux I__3531 (
            .O(N__20603),
            .I(N__20599));
    CEMux I__3530 (
            .O(N__20602),
            .I(N__20596));
    Odrv4 I__3529 (
            .O(N__20599),
            .I(\b2v_inst.N_463_i ));
    LocalMux I__3528 (
            .O(N__20596),
            .I(\b2v_inst.N_463_i ));
    InMux I__3527 (
            .O(N__20591),
            .I(N__20588));
    LocalMux I__3526 (
            .O(N__20588),
            .I(N__20585));
    Odrv12 I__3525 (
            .O(N__20585),
            .I(\b2v_inst.indice_4_i_a2_0_7_3_1 ));
    InMux I__3524 (
            .O(N__20582),
            .I(N__20579));
    LocalMux I__3523 (
            .O(N__20579),
            .I(\b2v_inst.N_432_1_tz ));
    InMux I__3522 (
            .O(N__20576),
            .I(N__20573));
    LocalMux I__3521 (
            .O(N__20573),
            .I(N__20570));
    Span4Mux_h I__3520 (
            .O(N__20570),
            .I(N__20567));
    Span4Mux_h I__3519 (
            .O(N__20567),
            .I(N__20564));
    Odrv4 I__3518 (
            .O(N__20564),
            .I(N_556_i));
    InMux I__3517 (
            .O(N__20561),
            .I(N__20558));
    LocalMux I__3516 (
            .O(N__20558),
            .I(\b2v_inst.indice_4_i_a2_0_7_2_1 ));
    InMux I__3515 (
            .O(N__20555),
            .I(N__20552));
    LocalMux I__3514 (
            .O(N__20552),
            .I(N__20549));
    Span4Mux_h I__3513 (
            .O(N__20549),
            .I(N__20546));
    Span4Mux_v I__3512 (
            .O(N__20546),
            .I(N__20543));
    Span4Mux_h I__3511 (
            .O(N__20543),
            .I(N__20540));
    Odrv4 I__3510 (
            .O(N__20540),
            .I(N_117_i));
    CascadeMux I__3509 (
            .O(N__20537),
            .I(\b2v_inst.addr_ram_energia_m0_3_cascade_ ));
    CascadeMux I__3508 (
            .O(N__20534),
            .I(N__20530));
    CascadeMux I__3507 (
            .O(N__20533),
            .I(N__20527));
    CascadeBuf I__3506 (
            .O(N__20530),
            .I(N__20524));
    CascadeBuf I__3505 (
            .O(N__20527),
            .I(N__20521));
    CascadeMux I__3504 (
            .O(N__20524),
            .I(N__20518));
    CascadeMux I__3503 (
            .O(N__20521),
            .I(N__20515));
    CascadeBuf I__3502 (
            .O(N__20518),
            .I(N__20512));
    CascadeBuf I__3501 (
            .O(N__20515),
            .I(N__20509));
    CascadeMux I__3500 (
            .O(N__20512),
            .I(N__20506));
    CascadeMux I__3499 (
            .O(N__20509),
            .I(N__20503));
    CascadeBuf I__3498 (
            .O(N__20506),
            .I(N__20500));
    CascadeBuf I__3497 (
            .O(N__20503),
            .I(N__20497));
    CascadeMux I__3496 (
            .O(N__20500),
            .I(N__20494));
    CascadeMux I__3495 (
            .O(N__20497),
            .I(N__20491));
    CascadeBuf I__3494 (
            .O(N__20494),
            .I(N__20488));
    CascadeBuf I__3493 (
            .O(N__20491),
            .I(N__20485));
    CascadeMux I__3492 (
            .O(N__20488),
            .I(N__20482));
    CascadeMux I__3491 (
            .O(N__20485),
            .I(N__20479));
    CascadeBuf I__3490 (
            .O(N__20482),
            .I(N__20476));
    CascadeBuf I__3489 (
            .O(N__20479),
            .I(N__20473));
    CascadeMux I__3488 (
            .O(N__20476),
            .I(N__20470));
    CascadeMux I__3487 (
            .O(N__20473),
            .I(N__20467));
    CascadeBuf I__3486 (
            .O(N__20470),
            .I(N__20464));
    CascadeBuf I__3485 (
            .O(N__20467),
            .I(N__20461));
    CascadeMux I__3484 (
            .O(N__20464),
            .I(N__20458));
    CascadeMux I__3483 (
            .O(N__20461),
            .I(N__20455));
    InMux I__3482 (
            .O(N__20458),
            .I(N__20452));
    InMux I__3481 (
            .O(N__20455),
            .I(N__20449));
    LocalMux I__3480 (
            .O(N__20452),
            .I(N__20444));
    LocalMux I__3479 (
            .O(N__20449),
            .I(N__20444));
    Span4Mux_v I__3478 (
            .O(N__20444),
            .I(N__20441));
    Span4Mux_h I__3477 (
            .O(N__20441),
            .I(N__20438));
    Span4Mux_h I__3476 (
            .O(N__20438),
            .I(N__20435));
    Odrv4 I__3475 (
            .O(N__20435),
            .I(SYNTHESIZED_WIRE_12_3));
    IoInMux I__3474 (
            .O(N__20432),
            .I(N__20429));
    LocalMux I__3473 (
            .O(N__20429),
            .I(N__20426));
    Span4Mux_s3_h I__3472 (
            .O(N__20426),
            .I(N__20422));
    InMux I__3471 (
            .O(N__20425),
            .I(N__20419));
    Span4Mux_v I__3470 (
            .O(N__20422),
            .I(N__20416));
    LocalMux I__3469 (
            .O(N__20419),
            .I(N__20413));
    Span4Mux_h I__3468 (
            .O(N__20416),
            .I(N__20410));
    Span4Mux_h I__3467 (
            .O(N__20413),
            .I(N__20407));
    Sp12to4 I__3466 (
            .O(N__20410),
            .I(N__20404));
    Span4Mux_h I__3465 (
            .O(N__20407),
            .I(N__20401));
    Odrv12 I__3464 (
            .O(N__20404),
            .I(leds_c_6));
    Odrv4 I__3463 (
            .O(N__20401),
            .I(leds_c_6));
    InMux I__3462 (
            .O(N__20396),
            .I(N__20393));
    LocalMux I__3461 (
            .O(N__20393),
            .I(N__20390));
    Sp12to4 I__3460 (
            .O(N__20390),
            .I(N__20387));
    Odrv12 I__3459 (
            .O(N__20387),
            .I(swit_c_0));
    CascadeMux I__3458 (
            .O(N__20384),
            .I(N__20381));
    InMux I__3457 (
            .O(N__20381),
            .I(N__20378));
    LocalMux I__3456 (
            .O(N__20378),
            .I(N__20375));
    Odrv12 I__3455 (
            .O(N__20375),
            .I(\b2v_inst.addr_ram_energia_m0_0 ));
    InMux I__3454 (
            .O(N__20372),
            .I(N__20369));
    LocalMux I__3453 (
            .O(N__20369),
            .I(N__20366));
    Span4Mux_v I__3452 (
            .O(N__20366),
            .I(N__20363));
    Sp12to4 I__3451 (
            .O(N__20363),
            .I(N__20360));
    Odrv12 I__3450 (
            .O(N__20360),
            .I(N_120_i));
    CascadeMux I__3449 (
            .O(N__20357),
            .I(\b2v_inst.N_432_1_cascade_ ));
    InMux I__3448 (
            .O(N__20354),
            .I(N__20351));
    LocalMux I__3447 (
            .O(N__20351),
            .I(N__20346));
    InMux I__3446 (
            .O(N__20350),
            .I(N__20341));
    InMux I__3445 (
            .O(N__20349),
            .I(N__20341));
    Span4Mux_h I__3444 (
            .O(N__20346),
            .I(N__20338));
    LocalMux I__3443 (
            .O(N__20341),
            .I(N__20334));
    Span4Mux_h I__3442 (
            .O(N__20338),
            .I(N__20331));
    InMux I__3441 (
            .O(N__20337),
            .I(N__20328));
    Odrv4 I__3440 (
            .O(N__20334),
            .I(\b2v_inst.un1_indice_cry_9_c_RNILAJPZ0 ));
    Odrv4 I__3439 (
            .O(N__20331),
            .I(\b2v_inst.un1_indice_cry_9_c_RNILAJPZ0 ));
    LocalMux I__3438 (
            .O(N__20328),
            .I(\b2v_inst.un1_indice_cry_9_c_RNILAJPZ0 ));
    InMux I__3437 (
            .O(N__20321),
            .I(N__20317));
    InMux I__3436 (
            .O(N__20320),
            .I(N__20314));
    LocalMux I__3435 (
            .O(N__20317),
            .I(N__20311));
    LocalMux I__3434 (
            .O(N__20314),
            .I(N__20307));
    Span4Mux_h I__3433 (
            .O(N__20311),
            .I(N__20304));
    InMux I__3432 (
            .O(N__20310),
            .I(N__20301));
    Span4Mux_h I__3431 (
            .O(N__20307),
            .I(N__20298));
    Span4Mux_h I__3430 (
            .O(N__20304),
            .I(N__20293));
    LocalMux I__3429 (
            .O(N__20301),
            .I(N__20293));
    Odrv4 I__3428 (
            .O(N__20298),
            .I(\b2v_inst.un1_indice_cry_7_c_RNIAFQGZ0 ));
    Odrv4 I__3427 (
            .O(N__20293),
            .I(\b2v_inst.un1_indice_cry_7_c_RNIAFQGZ0 ));
    CascadeMux I__3426 (
            .O(N__20288),
            .I(N__20285));
    InMux I__3425 (
            .O(N__20285),
            .I(N__20282));
    LocalMux I__3424 (
            .O(N__20282),
            .I(N__20279));
    Span4Mux_h I__3423 (
            .O(N__20279),
            .I(N__20276));
    Span4Mux_v I__3422 (
            .O(N__20276),
            .I(N__20273));
    Odrv4 I__3421 (
            .O(N__20273),
            .I(\b2v_inst.dir_mem_2Z0Z_0 ));
    CascadeMux I__3420 (
            .O(N__20270),
            .I(N__20266));
    InMux I__3419 (
            .O(N__20269),
            .I(N__20261));
    InMux I__3418 (
            .O(N__20266),
            .I(N__20261));
    LocalMux I__3417 (
            .O(N__20261),
            .I(N__20257));
    InMux I__3416 (
            .O(N__20260),
            .I(N__20254));
    Odrv4 I__3415 (
            .O(N__20257),
            .I(\b2v_inst.un8_dir_mem_2_cry_9_THRU_CO ));
    LocalMux I__3414 (
            .O(N__20254),
            .I(\b2v_inst.un8_dir_mem_2_cry_9_THRU_CO ));
    InMux I__3413 (
            .O(N__20249),
            .I(N__20245));
    InMux I__3412 (
            .O(N__20248),
            .I(N__20242));
    LocalMux I__3411 (
            .O(N__20245),
            .I(N__20236));
    LocalMux I__3410 (
            .O(N__20242),
            .I(N__20236));
    InMux I__3409 (
            .O(N__20241),
            .I(N__20233));
    Odrv4 I__3408 (
            .O(N__20236),
            .I(\b2v_inst.un8_dir_mem_2_cry_8_c_RNITIJEZ0 ));
    LocalMux I__3407 (
            .O(N__20233),
            .I(\b2v_inst.un8_dir_mem_2_cry_8_c_RNITIJEZ0 ));
    CascadeMux I__3406 (
            .O(N__20228),
            .I(N__20225));
    InMux I__3405 (
            .O(N__20225),
            .I(N__20222));
    LocalMux I__3404 (
            .O(N__20222),
            .I(N__20219));
    Span4Mux_v I__3403 (
            .O(N__20219),
            .I(N__20216));
    Odrv4 I__3402 (
            .O(N__20216),
            .I(\b2v_inst.dir_mem_2Z0Z_10 ));
    InMux I__3401 (
            .O(N__20213),
            .I(N__20205));
    InMux I__3400 (
            .O(N__20212),
            .I(N__20205));
    InMux I__3399 (
            .O(N__20211),
            .I(N__20200));
    InMux I__3398 (
            .O(N__20210),
            .I(N__20200));
    LocalMux I__3397 (
            .O(N__20205),
            .I(\b2v_inst.N_477 ));
    LocalMux I__3396 (
            .O(N__20200),
            .I(\b2v_inst.N_477 ));
    InMux I__3395 (
            .O(N__20195),
            .I(N__20192));
    LocalMux I__3394 (
            .O(N__20192),
            .I(N__20189));
    Span4Mux_v I__3393 (
            .O(N__20189),
            .I(N__20186));
    Span4Mux_v I__3392 (
            .O(N__20186),
            .I(N__20183));
    Span4Mux_v I__3391 (
            .O(N__20183),
            .I(N__20180));
    Sp12to4 I__3390 (
            .O(N__20180),
            .I(N__20177));
    Span12Mux_h I__3389 (
            .O(N__20177),
            .I(N__20174));
    Odrv12 I__3388 (
            .O(N__20174),
            .I(swit_c_1));
    CascadeMux I__3387 (
            .O(N__20171),
            .I(\b2v_inst.N_494_cascade_ ));
    CascadeMux I__3386 (
            .O(N__20168),
            .I(N__20165));
    InMux I__3385 (
            .O(N__20165),
            .I(N__20162));
    LocalMux I__3384 (
            .O(N__20162),
            .I(N__20159));
    Span4Mux_v I__3383 (
            .O(N__20159),
            .I(N__20156));
    Span4Mux_h I__3382 (
            .O(N__20156),
            .I(N__20153));
    Odrv4 I__3381 (
            .O(N__20153),
            .I(\b2v_inst.addr_ram_energia_m0_1 ));
    CascadeMux I__3380 (
            .O(N__20150),
            .I(N__20146));
    CascadeMux I__3379 (
            .O(N__20149),
            .I(N__20143));
    CascadeBuf I__3378 (
            .O(N__20146),
            .I(N__20140));
    CascadeBuf I__3377 (
            .O(N__20143),
            .I(N__20137));
    CascadeMux I__3376 (
            .O(N__20140),
            .I(N__20134));
    CascadeMux I__3375 (
            .O(N__20137),
            .I(N__20131));
    CascadeBuf I__3374 (
            .O(N__20134),
            .I(N__20128));
    CascadeBuf I__3373 (
            .O(N__20131),
            .I(N__20125));
    CascadeMux I__3372 (
            .O(N__20128),
            .I(N__20122));
    CascadeMux I__3371 (
            .O(N__20125),
            .I(N__20119));
    CascadeBuf I__3370 (
            .O(N__20122),
            .I(N__20116));
    CascadeBuf I__3369 (
            .O(N__20119),
            .I(N__20113));
    CascadeMux I__3368 (
            .O(N__20116),
            .I(N__20110));
    CascadeMux I__3367 (
            .O(N__20113),
            .I(N__20107));
    CascadeBuf I__3366 (
            .O(N__20110),
            .I(N__20104));
    CascadeBuf I__3365 (
            .O(N__20107),
            .I(N__20101));
    CascadeMux I__3364 (
            .O(N__20104),
            .I(N__20098));
    CascadeMux I__3363 (
            .O(N__20101),
            .I(N__20095));
    CascadeBuf I__3362 (
            .O(N__20098),
            .I(N__20092));
    CascadeBuf I__3361 (
            .O(N__20095),
            .I(N__20089));
    CascadeMux I__3360 (
            .O(N__20092),
            .I(N__20086));
    CascadeMux I__3359 (
            .O(N__20089),
            .I(N__20083));
    CascadeBuf I__3358 (
            .O(N__20086),
            .I(N__20080));
    CascadeBuf I__3357 (
            .O(N__20083),
            .I(N__20077));
    CascadeMux I__3356 (
            .O(N__20080),
            .I(N__20074));
    CascadeMux I__3355 (
            .O(N__20077),
            .I(N__20071));
    InMux I__3354 (
            .O(N__20074),
            .I(N__20068));
    InMux I__3353 (
            .O(N__20071),
            .I(N__20065));
    LocalMux I__3352 (
            .O(N__20068),
            .I(N__20062));
    LocalMux I__3351 (
            .O(N__20065),
            .I(N__20059));
    Span4Mux_v I__3350 (
            .O(N__20062),
            .I(N__20056));
    Span4Mux_v I__3349 (
            .O(N__20059),
            .I(N__20053));
    Span4Mux_h I__3348 (
            .O(N__20056),
            .I(N__20048));
    Span4Mux_h I__3347 (
            .O(N__20053),
            .I(N__20048));
    Span4Mux_h I__3346 (
            .O(N__20048),
            .I(N__20045));
    Odrv4 I__3345 (
            .O(N__20045),
            .I(SYNTHESIZED_WIRE_12_10));
    InMux I__3344 (
            .O(N__20042),
            .I(N__20039));
    LocalMux I__3343 (
            .O(N__20039),
            .I(N__20036));
    Span4Mux_h I__3342 (
            .O(N__20036),
            .I(N__20033));
    Sp12to4 I__3341 (
            .O(N__20033),
            .I(N__20030));
    Span12Mux_v I__3340 (
            .O(N__20030),
            .I(N__20027));
    Span12Mux_h I__3339 (
            .O(N__20027),
            .I(N__20024));
    Odrv12 I__3338 (
            .O(N__20024),
            .I(swit_c_2));
    CascadeMux I__3337 (
            .O(N__20021),
            .I(\b2v_inst.addr_ram_energia_m0_2_cascade_ ));
    CascadeMux I__3336 (
            .O(N__20018),
            .I(N__20014));
    CascadeMux I__3335 (
            .O(N__20017),
            .I(N__20011));
    CascadeBuf I__3334 (
            .O(N__20014),
            .I(N__20008));
    CascadeBuf I__3333 (
            .O(N__20011),
            .I(N__20005));
    CascadeMux I__3332 (
            .O(N__20008),
            .I(N__20002));
    CascadeMux I__3331 (
            .O(N__20005),
            .I(N__19999));
    CascadeBuf I__3330 (
            .O(N__20002),
            .I(N__19996));
    CascadeBuf I__3329 (
            .O(N__19999),
            .I(N__19993));
    CascadeMux I__3328 (
            .O(N__19996),
            .I(N__19990));
    CascadeMux I__3327 (
            .O(N__19993),
            .I(N__19987));
    CascadeBuf I__3326 (
            .O(N__19990),
            .I(N__19984));
    CascadeBuf I__3325 (
            .O(N__19987),
            .I(N__19981));
    CascadeMux I__3324 (
            .O(N__19984),
            .I(N__19978));
    CascadeMux I__3323 (
            .O(N__19981),
            .I(N__19975));
    CascadeBuf I__3322 (
            .O(N__19978),
            .I(N__19972));
    CascadeBuf I__3321 (
            .O(N__19975),
            .I(N__19969));
    CascadeMux I__3320 (
            .O(N__19972),
            .I(N__19966));
    CascadeMux I__3319 (
            .O(N__19969),
            .I(N__19963));
    CascadeBuf I__3318 (
            .O(N__19966),
            .I(N__19960));
    CascadeBuf I__3317 (
            .O(N__19963),
            .I(N__19957));
    CascadeMux I__3316 (
            .O(N__19960),
            .I(N__19954));
    CascadeMux I__3315 (
            .O(N__19957),
            .I(N__19951));
    CascadeBuf I__3314 (
            .O(N__19954),
            .I(N__19948));
    CascadeBuf I__3313 (
            .O(N__19951),
            .I(N__19945));
    CascadeMux I__3312 (
            .O(N__19948),
            .I(N__19942));
    CascadeMux I__3311 (
            .O(N__19945),
            .I(N__19939));
    InMux I__3310 (
            .O(N__19942),
            .I(N__19936));
    InMux I__3309 (
            .O(N__19939),
            .I(N__19933));
    LocalMux I__3308 (
            .O(N__19936),
            .I(N__19928));
    LocalMux I__3307 (
            .O(N__19933),
            .I(N__19928));
    Span4Mux_v I__3306 (
            .O(N__19928),
            .I(N__19925));
    Span4Mux_h I__3305 (
            .O(N__19925),
            .I(N__19922));
    Span4Mux_h I__3304 (
            .O(N__19922),
            .I(N__19919));
    Odrv4 I__3303 (
            .O(N__19919),
            .I(SYNTHESIZED_WIRE_12_2));
    InMux I__3302 (
            .O(N__19916),
            .I(N__19913));
    LocalMux I__3301 (
            .O(N__19913),
            .I(N__19910));
    Span12Mux_h I__3300 (
            .O(N__19910),
            .I(N__19907));
    Odrv12 I__3299 (
            .O(N__19907),
            .I(swit_c_5));
    CascadeMux I__3298 (
            .O(N__19904),
            .I(\b2v_inst.addr_ram_energia_m0_5_cascade_ ));
    CascadeMux I__3297 (
            .O(N__19901),
            .I(N__19897));
    CascadeMux I__3296 (
            .O(N__19900),
            .I(N__19894));
    CascadeBuf I__3295 (
            .O(N__19897),
            .I(N__19891));
    CascadeBuf I__3294 (
            .O(N__19894),
            .I(N__19888));
    CascadeMux I__3293 (
            .O(N__19891),
            .I(N__19885));
    CascadeMux I__3292 (
            .O(N__19888),
            .I(N__19882));
    CascadeBuf I__3291 (
            .O(N__19885),
            .I(N__19879));
    CascadeBuf I__3290 (
            .O(N__19882),
            .I(N__19876));
    CascadeMux I__3289 (
            .O(N__19879),
            .I(N__19873));
    CascadeMux I__3288 (
            .O(N__19876),
            .I(N__19870));
    CascadeBuf I__3287 (
            .O(N__19873),
            .I(N__19867));
    CascadeBuf I__3286 (
            .O(N__19870),
            .I(N__19864));
    CascadeMux I__3285 (
            .O(N__19867),
            .I(N__19861));
    CascadeMux I__3284 (
            .O(N__19864),
            .I(N__19858));
    CascadeBuf I__3283 (
            .O(N__19861),
            .I(N__19855));
    CascadeBuf I__3282 (
            .O(N__19858),
            .I(N__19852));
    CascadeMux I__3281 (
            .O(N__19855),
            .I(N__19849));
    CascadeMux I__3280 (
            .O(N__19852),
            .I(N__19846));
    CascadeBuf I__3279 (
            .O(N__19849),
            .I(N__19843));
    CascadeBuf I__3278 (
            .O(N__19846),
            .I(N__19840));
    CascadeMux I__3277 (
            .O(N__19843),
            .I(N__19837));
    CascadeMux I__3276 (
            .O(N__19840),
            .I(N__19834));
    CascadeBuf I__3275 (
            .O(N__19837),
            .I(N__19831));
    CascadeBuf I__3274 (
            .O(N__19834),
            .I(N__19828));
    CascadeMux I__3273 (
            .O(N__19831),
            .I(N__19825));
    CascadeMux I__3272 (
            .O(N__19828),
            .I(N__19822));
    InMux I__3271 (
            .O(N__19825),
            .I(N__19819));
    InMux I__3270 (
            .O(N__19822),
            .I(N__19816));
    LocalMux I__3269 (
            .O(N__19819),
            .I(N__19811));
    LocalMux I__3268 (
            .O(N__19816),
            .I(N__19811));
    Span4Mux_v I__3267 (
            .O(N__19811),
            .I(N__19808));
    Span4Mux_h I__3266 (
            .O(N__19808),
            .I(N__19805));
    Span4Mux_h I__3265 (
            .O(N__19805),
            .I(N__19802));
    Odrv4 I__3264 (
            .O(N__19802),
            .I(SYNTHESIZED_WIRE_12_5));
    InMux I__3263 (
            .O(N__19799),
            .I(N__19796));
    LocalMux I__3262 (
            .O(N__19796),
            .I(N__19793));
    Span4Mux_v I__3261 (
            .O(N__19793),
            .I(N__19790));
    Sp12to4 I__3260 (
            .O(N__19790),
            .I(N__19787));
    Span12Mux_v I__3259 (
            .O(N__19787),
            .I(N__19784));
    Span12Mux_h I__3258 (
            .O(N__19784),
            .I(N__19781));
    Odrv12 I__3257 (
            .O(N__19781),
            .I(swit_c_10));
    InMux I__3256 (
            .O(N__19778),
            .I(N__19775));
    LocalMux I__3255 (
            .O(N__19775),
            .I(\b2v_inst.addr_ram_energia_m0_10 ));
    InMux I__3254 (
            .O(N__19772),
            .I(N__19769));
    LocalMux I__3253 (
            .O(N__19769),
            .I(N__19766));
    Span4Mux_h I__3252 (
            .O(N__19766),
            .I(N__19763));
    Sp12to4 I__3251 (
            .O(N__19763),
            .I(N__19760));
    Odrv12 I__3250 (
            .O(N__19760),
            .I(swit_c_3));
    CascadeMux I__3249 (
            .O(N__19757),
            .I(\b2v_inst.N_514_cascade_ ));
    InMux I__3248 (
            .O(N__19754),
            .I(N__19751));
    LocalMux I__3247 (
            .O(N__19751),
            .I(N__19748));
    Span4Mux_h I__3246 (
            .O(N__19748),
            .I(N__19745));
    Span4Mux_v I__3245 (
            .O(N__19745),
            .I(N__19742));
    Span4Mux_h I__3244 (
            .O(N__19742),
            .I(N__19739));
    Span4Mux_h I__3243 (
            .O(N__19739),
            .I(N__19736));
    Odrv4 I__3242 (
            .O(N__19736),
            .I(N_116_i));
    InMux I__3241 (
            .O(N__19733),
            .I(N__19730));
    LocalMux I__3240 (
            .O(N__19730),
            .I(N__19725));
    InMux I__3239 (
            .O(N__19729),
            .I(N__19720));
    InMux I__3238 (
            .O(N__19728),
            .I(N__19720));
    Odrv4 I__3237 (
            .O(N__19725),
            .I(\b2v_inst.stateZ0Z_16 ));
    LocalMux I__3236 (
            .O(N__19720),
            .I(\b2v_inst.stateZ0Z_16 ));
    InMux I__3235 (
            .O(N__19715),
            .I(N__19712));
    LocalMux I__3234 (
            .O(N__19712),
            .I(N__19709));
    Span4Mux_h I__3233 (
            .O(N__19709),
            .I(N__19706));
    Span4Mux_h I__3232 (
            .O(N__19706),
            .I(N__19703));
    Odrv4 I__3231 (
            .O(N__19703),
            .I(N_548_i));
    CascadeMux I__3230 (
            .O(N__19700),
            .I(N__19697));
    InMux I__3229 (
            .O(N__19697),
            .I(N__19694));
    LocalMux I__3228 (
            .O(N__19694),
            .I(N__19688));
    CascadeMux I__3227 (
            .O(N__19693),
            .I(N__19685));
    CascadeMux I__3226 (
            .O(N__19692),
            .I(N__19682));
    InMux I__3225 (
            .O(N__19691),
            .I(N__19679));
    Span4Mux_v I__3224 (
            .O(N__19688),
            .I(N__19676));
    InMux I__3223 (
            .O(N__19685),
            .I(N__19671));
    InMux I__3222 (
            .O(N__19682),
            .I(N__19671));
    LocalMux I__3221 (
            .O(N__19679),
            .I(\b2v_inst.stateZ0Z_0 ));
    Odrv4 I__3220 (
            .O(N__19676),
            .I(\b2v_inst.stateZ0Z_0 ));
    LocalMux I__3219 (
            .O(N__19671),
            .I(\b2v_inst.stateZ0Z_0 ));
    CascadeMux I__3218 (
            .O(N__19664),
            .I(\b2v_inst.N_692_cascade_ ));
    CascadeMux I__3217 (
            .O(N__19661),
            .I(\b2v_inst.addr_ram_iv_i_0_0_3_cascade_ ));
    CascadeMux I__3216 (
            .O(N__19658),
            .I(N__19655));
    CascadeBuf I__3215 (
            .O(N__19655),
            .I(N__19652));
    CascadeMux I__3214 (
            .O(N__19652),
            .I(N__19648));
    CascadeMux I__3213 (
            .O(N__19651),
            .I(N__19645));
    CascadeBuf I__3212 (
            .O(N__19648),
            .I(N__19642));
    CascadeBuf I__3211 (
            .O(N__19645),
            .I(N__19639));
    CascadeMux I__3210 (
            .O(N__19642),
            .I(N__19636));
    CascadeMux I__3209 (
            .O(N__19639),
            .I(N__19633));
    CascadeBuf I__3208 (
            .O(N__19636),
            .I(N__19630));
    CascadeBuf I__3207 (
            .O(N__19633),
            .I(N__19627));
    CascadeMux I__3206 (
            .O(N__19630),
            .I(N__19624));
    CascadeMux I__3205 (
            .O(N__19627),
            .I(N__19621));
    CascadeBuf I__3204 (
            .O(N__19624),
            .I(N__19618));
    CascadeBuf I__3203 (
            .O(N__19621),
            .I(N__19615));
    CascadeMux I__3202 (
            .O(N__19618),
            .I(N__19612));
    CascadeMux I__3201 (
            .O(N__19615),
            .I(N__19609));
    CascadeBuf I__3200 (
            .O(N__19612),
            .I(N__19606));
    CascadeBuf I__3199 (
            .O(N__19609),
            .I(N__19603));
    CascadeMux I__3198 (
            .O(N__19606),
            .I(N__19600));
    CascadeMux I__3197 (
            .O(N__19603),
            .I(N__19597));
    InMux I__3196 (
            .O(N__19600),
            .I(N__19594));
    CascadeBuf I__3195 (
            .O(N__19597),
            .I(N__19591));
    LocalMux I__3194 (
            .O(N__19594),
            .I(N__19588));
    CascadeMux I__3193 (
            .O(N__19591),
            .I(N__19585));
    Span4Mux_v I__3192 (
            .O(N__19588),
            .I(N__19582));
    InMux I__3191 (
            .O(N__19585),
            .I(N__19579));
    Span4Mux_h I__3190 (
            .O(N__19582),
            .I(N__19576));
    LocalMux I__3189 (
            .O(N__19579),
            .I(N__19573));
    Span4Mux_h I__3188 (
            .O(N__19576),
            .I(N__19570));
    Odrv12 I__3187 (
            .O(N__19573),
            .I(indice_RNIIU233_3));
    Odrv4 I__3186 (
            .O(N__19570),
            .I(indice_RNIIU233_3));
    InMux I__3185 (
            .O(N__19565),
            .I(N__19562));
    LocalMux I__3184 (
            .O(N__19562),
            .I(N__19559));
    Span4Mux_h I__3183 (
            .O(N__19559),
            .I(N__19556));
    Span4Mux_v I__3182 (
            .O(N__19556),
            .I(N__19553));
    Odrv4 I__3181 (
            .O(N__19553),
            .I(\b2v_inst.dir_mem_3Z0Z_3 ));
    InMux I__3180 (
            .O(N__19550),
            .I(N__19547));
    LocalMux I__3179 (
            .O(N__19547),
            .I(N__19544));
    Span4Mux_v I__3178 (
            .O(N__19544),
            .I(N__19541));
    Odrv4 I__3177 (
            .O(N__19541),
            .I(\b2v_inst.dir_mem_1Z0Z_3 ));
    InMux I__3176 (
            .O(N__19538),
            .I(N__19535));
    LocalMux I__3175 (
            .O(N__19535),
            .I(\b2v_inst.addr_ram_iv_i_0_1_3 ));
    InMux I__3174 (
            .O(N__19532),
            .I(N__19529));
    LocalMux I__3173 (
            .O(N__19529),
            .I(\b2v_inst.dir_memZ0Z_0 ));
    InMux I__3172 (
            .O(N__19526),
            .I(N__19522));
    InMux I__3171 (
            .O(N__19525),
            .I(N__19519));
    LocalMux I__3170 (
            .O(N__19522),
            .I(N__19516));
    LocalMux I__3169 (
            .O(N__19519),
            .I(N__19511));
    Span4Mux_v I__3168 (
            .O(N__19516),
            .I(N__19511));
    Odrv4 I__3167 (
            .O(N__19511),
            .I(\b2v_inst.N_618_6 ));
    InMux I__3166 (
            .O(N__19508),
            .I(N__19505));
    LocalMux I__3165 (
            .O(N__19505),
            .I(N__19502));
    Odrv4 I__3164 (
            .O(N__19502),
            .I(\b2v_inst.dir_mem_1Z0Z_7 ));
    InMux I__3163 (
            .O(N__19499),
            .I(N__19496));
    LocalMux I__3162 (
            .O(N__19496),
            .I(N__19493));
    Span4Mux_v I__3161 (
            .O(N__19493),
            .I(N__19490));
    Span4Mux_h I__3160 (
            .O(N__19490),
            .I(N__19487));
    Odrv4 I__3159 (
            .O(N__19487),
            .I(\b2v_inst.dir_mem_3Z0Z_7 ));
    CascadeMux I__3158 (
            .O(N__19484),
            .I(\b2v_inst.N_488_cascade_ ));
    InMux I__3157 (
            .O(N__19481),
            .I(N__19478));
    LocalMux I__3156 (
            .O(N__19478),
            .I(\b2v_inst.addr_ram_iv_i_0_0_7 ));
    CascadeMux I__3155 (
            .O(N__19475),
            .I(\b2v_inst.addr_ram_iv_i_0_1_7_cascade_ ));
    CascadeMux I__3154 (
            .O(N__19472),
            .I(N__19468));
    CascadeMux I__3153 (
            .O(N__19471),
            .I(N__19465));
    CascadeBuf I__3152 (
            .O(N__19468),
            .I(N__19462));
    CascadeBuf I__3151 (
            .O(N__19465),
            .I(N__19459));
    CascadeMux I__3150 (
            .O(N__19462),
            .I(N__19456));
    CascadeMux I__3149 (
            .O(N__19459),
            .I(N__19453));
    CascadeBuf I__3148 (
            .O(N__19456),
            .I(N__19450));
    CascadeBuf I__3147 (
            .O(N__19453),
            .I(N__19447));
    CascadeMux I__3146 (
            .O(N__19450),
            .I(N__19444));
    CascadeMux I__3145 (
            .O(N__19447),
            .I(N__19441));
    CascadeBuf I__3144 (
            .O(N__19444),
            .I(N__19438));
    CascadeBuf I__3143 (
            .O(N__19441),
            .I(N__19435));
    CascadeMux I__3142 (
            .O(N__19438),
            .I(N__19432));
    CascadeMux I__3141 (
            .O(N__19435),
            .I(N__19429));
    CascadeBuf I__3140 (
            .O(N__19432),
            .I(N__19426));
    CascadeBuf I__3139 (
            .O(N__19429),
            .I(N__19423));
    CascadeMux I__3138 (
            .O(N__19426),
            .I(N__19420));
    CascadeMux I__3137 (
            .O(N__19423),
            .I(N__19417));
    CascadeBuf I__3136 (
            .O(N__19420),
            .I(N__19414));
    CascadeBuf I__3135 (
            .O(N__19417),
            .I(N__19411));
    CascadeMux I__3134 (
            .O(N__19414),
            .I(N__19408));
    CascadeMux I__3133 (
            .O(N__19411),
            .I(N__19405));
    InMux I__3132 (
            .O(N__19408),
            .I(N__19402));
    InMux I__3131 (
            .O(N__19405),
            .I(N__19399));
    LocalMux I__3130 (
            .O(N__19402),
            .I(N__19394));
    LocalMux I__3129 (
            .O(N__19399),
            .I(N__19394));
    Span12Mux_v I__3128 (
            .O(N__19394),
            .I(N__19391));
    Odrv12 I__3127 (
            .O(N__19391),
            .I(indice_RNI6J333_7));
    InMux I__3126 (
            .O(N__19388),
            .I(N__19385));
    LocalMux I__3125 (
            .O(N__19385),
            .I(N__19382));
    Span4Mux_v I__3124 (
            .O(N__19382),
            .I(N__19379));
    Odrv4 I__3123 (
            .O(N__19379),
            .I(\b2v_inst.state_RNO_0Z0Z_29 ));
    InMux I__3122 (
            .O(N__19376),
            .I(N__19373));
    LocalMux I__3121 (
            .O(N__19373),
            .I(N__19370));
    Span4Mux_v I__3120 (
            .O(N__19370),
            .I(N__19367));
    Odrv4 I__3119 (
            .O(N__19367),
            .I(\b2v_inst.dir_mem_1Z0Z_0 ));
    CascadeMux I__3118 (
            .O(N__19364),
            .I(N__19361));
    InMux I__3117 (
            .O(N__19361),
            .I(N__19358));
    LocalMux I__3116 (
            .O(N__19358),
            .I(N__19355));
    Span4Mux_v I__3115 (
            .O(N__19355),
            .I(N__19352));
    Span4Mux_h I__3114 (
            .O(N__19352),
            .I(N__19349));
    Odrv4 I__3113 (
            .O(N__19349),
            .I(\b2v_inst.dir_mem_3Z0Z_0 ));
    InMux I__3112 (
            .O(N__19346),
            .I(N__19343));
    LocalMux I__3111 (
            .O(N__19343),
            .I(N__19340));
    Span4Mux_v I__3110 (
            .O(N__19340),
            .I(N__19337));
    Odrv4 I__3109 (
            .O(N__19337),
            .I(\b2v_inst.dir_mem_2Z0Z_3 ));
    InMux I__3108 (
            .O(N__19334),
            .I(N__19331));
    LocalMux I__3107 (
            .O(N__19331),
            .I(N__19328));
    Span4Mux_v I__3106 (
            .O(N__19328),
            .I(N__19325));
    Odrv4 I__3105 (
            .O(N__19325),
            .I(\b2v_inst.dir_memZ0Z_3 ));
    InMux I__3104 (
            .O(N__19322),
            .I(N__19319));
    LocalMux I__3103 (
            .O(N__19319),
            .I(N__19316));
    Span4Mux_h I__3102 (
            .O(N__19316),
            .I(N__19313));
    Odrv4 I__3101 (
            .O(N__19313),
            .I(\b2v_inst.dir_mem_3Z0Z_1 ));
    InMux I__3100 (
            .O(N__19310),
            .I(N__19307));
    LocalMux I__3099 (
            .O(N__19307),
            .I(N__19304));
    Odrv4 I__3098 (
            .O(N__19304),
            .I(\b2v_inst.dir_memZ0Z_1 ));
    CascadeMux I__3097 (
            .O(N__19301),
            .I(N__19298));
    InMux I__3096 (
            .O(N__19298),
            .I(N__19295));
    LocalMux I__3095 (
            .O(N__19295),
            .I(N__19292));
    Span4Mux_v I__3094 (
            .O(N__19292),
            .I(N__19289));
    Odrv4 I__3093 (
            .O(N__19289),
            .I(\b2v_inst.dir_mem_2Z0Z_1 ));
    InMux I__3092 (
            .O(N__19286),
            .I(N__19283));
    LocalMux I__3091 (
            .O(N__19283),
            .I(N__19279));
    InMux I__3090 (
            .O(N__19282),
            .I(N__19276));
    Span4Mux_h I__3089 (
            .O(N__19279),
            .I(N__19270));
    LocalMux I__3088 (
            .O(N__19276),
            .I(N__19270));
    CascadeMux I__3087 (
            .O(N__19275),
            .I(N__19267));
    Span4Mux_h I__3086 (
            .O(N__19270),
            .I(N__19264));
    InMux I__3085 (
            .O(N__19267),
            .I(N__19261));
    Odrv4 I__3084 (
            .O(N__19264),
            .I(\b2v_inst.un8_dir_mem_1_cry_0_c_RNI4SNCZ0 ));
    LocalMux I__3083 (
            .O(N__19261),
            .I(\b2v_inst.un8_dir_mem_1_cry_0_c_RNI4SNCZ0 ));
    InMux I__3082 (
            .O(N__19256),
            .I(N__19253));
    LocalMux I__3081 (
            .O(N__19253),
            .I(\b2v_inst.dir_mem_1Z0Z_1 ));
    InMux I__3080 (
            .O(N__19250),
            .I(N__19236));
    InMux I__3079 (
            .O(N__19249),
            .I(N__19236));
    InMux I__3078 (
            .O(N__19248),
            .I(N__19229));
    InMux I__3077 (
            .O(N__19247),
            .I(N__19229));
    InMux I__3076 (
            .O(N__19246),
            .I(N__19229));
    InMux I__3075 (
            .O(N__19245),
            .I(N__19218));
    InMux I__3074 (
            .O(N__19244),
            .I(N__19218));
    InMux I__3073 (
            .O(N__19243),
            .I(N__19218));
    InMux I__3072 (
            .O(N__19242),
            .I(N__19218));
    InMux I__3071 (
            .O(N__19241),
            .I(N__19218));
    LocalMux I__3070 (
            .O(N__19236),
            .I(\b2v_inst.dir_mem_115lt11 ));
    LocalMux I__3069 (
            .O(N__19229),
            .I(\b2v_inst.dir_mem_115lt11 ));
    LocalMux I__3068 (
            .O(N__19218),
            .I(\b2v_inst.dir_mem_115lt11 ));
    InMux I__3067 (
            .O(N__19211),
            .I(N__19207));
    InMux I__3066 (
            .O(N__19210),
            .I(N__19204));
    LocalMux I__3065 (
            .O(N__19207),
            .I(N__19201));
    LocalMux I__3064 (
            .O(N__19204),
            .I(N__19195));
    Span4Mux_v I__3063 (
            .O(N__19201),
            .I(N__19195));
    CascadeMux I__3062 (
            .O(N__19200),
            .I(N__19192));
    Span4Mux_h I__3061 (
            .O(N__19195),
            .I(N__19189));
    InMux I__3060 (
            .O(N__19192),
            .I(N__19186));
    Odrv4 I__3059 (
            .O(N__19189),
            .I(\b2v_inst.indice_RNILHHBZ0Z_2 ));
    LocalMux I__3058 (
            .O(N__19186),
            .I(\b2v_inst.indice_RNILHHBZ0Z_2 ));
    CascadeMux I__3057 (
            .O(N__19181),
            .I(N__19175));
    CascadeMux I__3056 (
            .O(N__19180),
            .I(N__19172));
    CascadeMux I__3055 (
            .O(N__19179),
            .I(N__19169));
    InMux I__3054 (
            .O(N__19178),
            .I(N__19159));
    InMux I__3053 (
            .O(N__19175),
            .I(N__19159));
    InMux I__3052 (
            .O(N__19172),
            .I(N__19156));
    InMux I__3051 (
            .O(N__19169),
            .I(N__19151));
    InMux I__3050 (
            .O(N__19168),
            .I(N__19151));
    InMux I__3049 (
            .O(N__19167),
            .I(N__19142));
    InMux I__3048 (
            .O(N__19166),
            .I(N__19142));
    InMux I__3047 (
            .O(N__19165),
            .I(N__19142));
    InMux I__3046 (
            .O(N__19164),
            .I(N__19142));
    LocalMux I__3045 (
            .O(N__19159),
            .I(N__19139));
    LocalMux I__3044 (
            .O(N__19156),
            .I(\b2v_inst.dir_mem_115lto11_0 ));
    LocalMux I__3043 (
            .O(N__19151),
            .I(\b2v_inst.dir_mem_115lto11_0 ));
    LocalMux I__3042 (
            .O(N__19142),
            .I(\b2v_inst.dir_mem_115lto11_0 ));
    Odrv12 I__3041 (
            .O(N__19139),
            .I(\b2v_inst.dir_mem_115lto11_0 ));
    InMux I__3040 (
            .O(N__19130),
            .I(N__19127));
    LocalMux I__3039 (
            .O(N__19127),
            .I(N__19124));
    Span12Mux_h I__3038 (
            .O(N__19124),
            .I(N__19120));
    InMux I__3037 (
            .O(N__19123),
            .I(N__19117));
    Odrv12 I__3036 (
            .O(N__19120),
            .I(\b2v_inst.un8_dir_mem_1_cry_1_c_RNI6VOCZ0 ));
    LocalMux I__3035 (
            .O(N__19117),
            .I(\b2v_inst.un8_dir_mem_1_cry_1_c_RNI6VOCZ0 ));
    CEMux I__3034 (
            .O(N__19112),
            .I(N__19108));
    CEMux I__3033 (
            .O(N__19111),
            .I(N__19105));
    LocalMux I__3032 (
            .O(N__19108),
            .I(N__19101));
    LocalMux I__3031 (
            .O(N__19105),
            .I(N__19098));
    CEMux I__3030 (
            .O(N__19104),
            .I(N__19095));
    Span4Mux_v I__3029 (
            .O(N__19101),
            .I(N__19092));
    Span4Mux_h I__3028 (
            .O(N__19098),
            .I(N__19089));
    LocalMux I__3027 (
            .O(N__19095),
            .I(N__19086));
    Odrv4 I__3026 (
            .O(N__19092),
            .I(\b2v_inst.N_363_i ));
    Odrv4 I__3025 (
            .O(N__19089),
            .I(\b2v_inst.N_363_i ));
    Odrv4 I__3024 (
            .O(N__19086),
            .I(\b2v_inst.N_363_i ));
    InMux I__3023 (
            .O(N__19079),
            .I(N__19076));
    LocalMux I__3022 (
            .O(N__19076),
            .I(N__19073));
    Odrv4 I__3021 (
            .O(N__19073),
            .I(\b2v_inst.dir_mem_2Z0Z_6 ));
    CascadeMux I__3020 (
            .O(N__19070),
            .I(\b2v_inst.N_489_cascade_ ));
    InMux I__3019 (
            .O(N__19067),
            .I(N__19064));
    LocalMux I__3018 (
            .O(N__19064),
            .I(N__19061));
    Span4Mux_h I__3017 (
            .O(N__19061),
            .I(N__19056));
    InMux I__3016 (
            .O(N__19060),
            .I(N__19053));
    InMux I__3015 (
            .O(N__19059),
            .I(N__19050));
    Odrv4 I__3014 (
            .O(N__19056),
            .I(\b2v_inst.un8_dir_mem_2_cry_1_c_RNI88LLZ0 ));
    LocalMux I__3013 (
            .O(N__19053),
            .I(\b2v_inst.un8_dir_mem_2_cry_1_c_RNI88LLZ0 ));
    LocalMux I__3012 (
            .O(N__19050),
            .I(\b2v_inst.un8_dir_mem_2_cry_1_c_RNI88LLZ0 ));
    InMux I__3011 (
            .O(N__19043),
            .I(N__19040));
    LocalMux I__3010 (
            .O(N__19040),
            .I(N__19037));
    Span4Mux_h I__3009 (
            .O(N__19037),
            .I(N__19032));
    InMux I__3008 (
            .O(N__19036),
            .I(N__19029));
    InMux I__3007 (
            .O(N__19035),
            .I(N__19026));
    Odrv4 I__3006 (
            .O(N__19032),
            .I(\b2v_inst.un8_dir_mem_2_cry_2_c_RNIABMLZ0 ));
    LocalMux I__3005 (
            .O(N__19029),
            .I(\b2v_inst.un8_dir_mem_2_cry_2_c_RNIABMLZ0 ));
    LocalMux I__3004 (
            .O(N__19026),
            .I(\b2v_inst.un8_dir_mem_2_cry_2_c_RNIABMLZ0 ));
    CascadeMux I__3003 (
            .O(N__19019),
            .I(N__19016));
    InMux I__3002 (
            .O(N__19016),
            .I(N__19013));
    LocalMux I__3001 (
            .O(N__19013),
            .I(N__19010));
    Span4Mux_v I__3000 (
            .O(N__19010),
            .I(N__19007));
    Odrv4 I__2999 (
            .O(N__19007),
            .I(\b2v_inst.dir_mem_2Z0Z_4 ));
    InMux I__2998 (
            .O(N__19004),
            .I(N__19001));
    LocalMux I__2997 (
            .O(N__19001),
            .I(N__18998));
    Span4Mux_h I__2996 (
            .O(N__18998),
            .I(N__18994));
    InMux I__2995 (
            .O(N__18997),
            .I(N__18991));
    Odrv4 I__2994 (
            .O(N__18994),
            .I(\b2v_inst.un8_dir_mem_2_cry_3_c_RNICENLZ0 ));
    LocalMux I__2993 (
            .O(N__18991),
            .I(\b2v_inst.un8_dir_mem_2_cry_3_c_RNICENLZ0 ));
    InMux I__2992 (
            .O(N__18986),
            .I(N__18983));
    LocalMux I__2991 (
            .O(N__18983),
            .I(N__18980));
    Span4Mux_v I__2990 (
            .O(N__18980),
            .I(N__18976));
    InMux I__2989 (
            .O(N__18979),
            .I(N__18973));
    Odrv4 I__2988 (
            .O(N__18976),
            .I(\b2v_inst.un8_dir_mem_2_cry_4_c_RNIEHOLZ0 ));
    LocalMux I__2987 (
            .O(N__18973),
            .I(\b2v_inst.un8_dir_mem_2_cry_4_c_RNIEHOLZ0 ));
    InMux I__2986 (
            .O(N__18968),
            .I(N__18961));
    InMux I__2985 (
            .O(N__18967),
            .I(N__18961));
    InMux I__2984 (
            .O(N__18966),
            .I(N__18958));
    LocalMux I__2983 (
            .O(N__18961),
            .I(N__18953));
    LocalMux I__2982 (
            .O(N__18958),
            .I(N__18953));
    Odrv12 I__2981 (
            .O(N__18953),
            .I(\b2v_inst.un8_dir_mem_1_cry_10_THRU_CO ));
    InMux I__2980 (
            .O(N__18950),
            .I(N__18943));
    InMux I__2979 (
            .O(N__18949),
            .I(N__18943));
    InMux I__2978 (
            .O(N__18948),
            .I(N__18940));
    LocalMux I__2977 (
            .O(N__18943),
            .I(N__18935));
    LocalMux I__2976 (
            .O(N__18940),
            .I(N__18935));
    Odrv12 I__2975 (
            .O(N__18935),
            .I(\b2v_inst.un8_dir_mem_1_cry_9_c_RNITCOLZ0 ));
    InMux I__2974 (
            .O(N__18932),
            .I(N__18929));
    LocalMux I__2973 (
            .O(N__18929),
            .I(\b2v_inst.dir_mem_1Z0Z_8 ));
    CascadeMux I__2972 (
            .O(N__18926),
            .I(N__18923));
    InMux I__2971 (
            .O(N__18923),
            .I(N__18920));
    LocalMux I__2970 (
            .O(N__18920),
            .I(N__18917));
    Odrv4 I__2969 (
            .O(N__18917),
            .I(\b2v_inst.dir_mem_3Z0Z_8 ));
    InMux I__2968 (
            .O(N__18914),
            .I(N__18911));
    LocalMux I__2967 (
            .O(N__18911),
            .I(N__18908));
    Span4Mux_h I__2966 (
            .O(N__18908),
            .I(N__18905));
    Sp12to4 I__2965 (
            .O(N__18905),
            .I(N__18902));
    Span12Mux_v I__2964 (
            .O(N__18902),
            .I(N__18899));
    Span12Mux_h I__2963 (
            .O(N__18899),
            .I(N__18896));
    Odrv12 I__2962 (
            .O(N__18896),
            .I(swit_c_7));
    CascadeMux I__2961 (
            .O(N__18893),
            .I(N__18890));
    InMux I__2960 (
            .O(N__18890),
            .I(N__18887));
    LocalMux I__2959 (
            .O(N__18887),
            .I(N__18884));
    Span4Mux_h I__2958 (
            .O(N__18884),
            .I(N__18881));
    Span4Mux_h I__2957 (
            .O(N__18881),
            .I(N__18878));
    Odrv4 I__2956 (
            .O(N__18878),
            .I(\b2v_inst.addr_ram_energia_m0_7 ));
    IoInMux I__2955 (
            .O(N__18875),
            .I(N__18871));
    InMux I__2954 (
            .O(N__18874),
            .I(N__18868));
    LocalMux I__2953 (
            .O(N__18871),
            .I(N__18865));
    LocalMux I__2952 (
            .O(N__18868),
            .I(N__18862));
    Span4Mux_s3_h I__2951 (
            .O(N__18865),
            .I(N__18859));
    Span4Mux_v I__2950 (
            .O(N__18862),
            .I(N__18856));
    Span4Mux_h I__2949 (
            .O(N__18859),
            .I(N__18853));
    Span4Mux_h I__2948 (
            .O(N__18856),
            .I(N__18850));
    Odrv4 I__2947 (
            .O(N__18853),
            .I(leds_c_12));
    Odrv4 I__2946 (
            .O(N__18850),
            .I(leds_c_12));
    InMux I__2945 (
            .O(N__18845),
            .I(N__18842));
    LocalMux I__2944 (
            .O(N__18842),
            .I(N__18838));
    InMux I__2943 (
            .O(N__18841),
            .I(N__18835));
    Span4Mux_v I__2942 (
            .O(N__18838),
            .I(N__18831));
    LocalMux I__2941 (
            .O(N__18835),
            .I(N__18828));
    InMux I__2940 (
            .O(N__18834),
            .I(N__18825));
    Span4Mux_h I__2939 (
            .O(N__18831),
            .I(N__18820));
    Span4Mux_v I__2938 (
            .O(N__18828),
            .I(N__18820));
    LocalMux I__2937 (
            .O(N__18825),
            .I(N__18817));
    Odrv4 I__2936 (
            .O(N__18820),
            .I(\b2v_inst.un1_indice_cry_4_c_RNI46NGZ0 ));
    Odrv4 I__2935 (
            .O(N__18817),
            .I(\b2v_inst.un1_indice_cry_4_c_RNI46NGZ0 ));
    InMux I__2934 (
            .O(N__18812),
            .I(N__18809));
    LocalMux I__2933 (
            .O(N__18809),
            .I(N__18805));
    InMux I__2932 (
            .O(N__18808),
            .I(N__18802));
    Span4Mux_v I__2931 (
            .O(N__18805),
            .I(N__18797));
    LocalMux I__2930 (
            .O(N__18802),
            .I(N__18797));
    Span4Mux_h I__2929 (
            .O(N__18797),
            .I(N__18793));
    InMux I__2928 (
            .O(N__18796),
            .I(N__18790));
    Odrv4 I__2927 (
            .O(N__18793),
            .I(\b2v_inst.un1_indice_cry_8_c_RNICIRGZ0 ));
    LocalMux I__2926 (
            .O(N__18790),
            .I(\b2v_inst.un1_indice_cry_8_c_RNICIRGZ0 ));
    InMux I__2925 (
            .O(N__18785),
            .I(N__18781));
    InMux I__2924 (
            .O(N__18784),
            .I(N__18777));
    LocalMux I__2923 (
            .O(N__18781),
            .I(N__18774));
    CascadeMux I__2922 (
            .O(N__18780),
            .I(N__18771));
    LocalMux I__2921 (
            .O(N__18777),
            .I(N__18768));
    Span4Mux_h I__2920 (
            .O(N__18774),
            .I(N__18765));
    InMux I__2919 (
            .O(N__18771),
            .I(N__18762));
    Span4Mux_h I__2918 (
            .O(N__18768),
            .I(N__18759));
    Span4Mux_h I__2917 (
            .O(N__18765),
            .I(N__18754));
    LocalMux I__2916 (
            .O(N__18762),
            .I(N__18754));
    Odrv4 I__2915 (
            .O(N__18759),
            .I(\b2v_inst.dir_mem_316lto7 ));
    Odrv4 I__2914 (
            .O(N__18754),
            .I(\b2v_inst.dir_mem_316lto7 ));
    InMux I__2913 (
            .O(N__18749),
            .I(N__18746));
    LocalMux I__2912 (
            .O(N__18746),
            .I(N__18743));
    Span4Mux_h I__2911 (
            .O(N__18743),
            .I(N__18740));
    Sp12to4 I__2910 (
            .O(N__18740),
            .I(N__18737));
    Span12Mux_v I__2909 (
            .O(N__18737),
            .I(N__18734));
    Span12Mux_h I__2908 (
            .O(N__18734),
            .I(N__18731));
    Odrv12 I__2907 (
            .O(N__18731),
            .I(swit_c_6));
    CascadeMux I__2906 (
            .O(N__18728),
            .I(\b2v_inst.addr_ram_energia_m0_6_cascade_ ));
    CascadeMux I__2905 (
            .O(N__18725),
            .I(N__18721));
    CascadeMux I__2904 (
            .O(N__18724),
            .I(N__18718));
    CascadeBuf I__2903 (
            .O(N__18721),
            .I(N__18715));
    CascadeBuf I__2902 (
            .O(N__18718),
            .I(N__18712));
    CascadeMux I__2901 (
            .O(N__18715),
            .I(N__18709));
    CascadeMux I__2900 (
            .O(N__18712),
            .I(N__18706));
    CascadeBuf I__2899 (
            .O(N__18709),
            .I(N__18703));
    CascadeBuf I__2898 (
            .O(N__18706),
            .I(N__18700));
    CascadeMux I__2897 (
            .O(N__18703),
            .I(N__18697));
    CascadeMux I__2896 (
            .O(N__18700),
            .I(N__18694));
    CascadeBuf I__2895 (
            .O(N__18697),
            .I(N__18691));
    CascadeBuf I__2894 (
            .O(N__18694),
            .I(N__18688));
    CascadeMux I__2893 (
            .O(N__18691),
            .I(N__18685));
    CascadeMux I__2892 (
            .O(N__18688),
            .I(N__18682));
    CascadeBuf I__2891 (
            .O(N__18685),
            .I(N__18679));
    CascadeBuf I__2890 (
            .O(N__18682),
            .I(N__18676));
    CascadeMux I__2889 (
            .O(N__18679),
            .I(N__18673));
    CascadeMux I__2888 (
            .O(N__18676),
            .I(N__18670));
    CascadeBuf I__2887 (
            .O(N__18673),
            .I(N__18667));
    CascadeBuf I__2886 (
            .O(N__18670),
            .I(N__18664));
    CascadeMux I__2885 (
            .O(N__18667),
            .I(N__18661));
    CascadeMux I__2884 (
            .O(N__18664),
            .I(N__18658));
    CascadeBuf I__2883 (
            .O(N__18661),
            .I(N__18655));
    CascadeBuf I__2882 (
            .O(N__18658),
            .I(N__18652));
    CascadeMux I__2881 (
            .O(N__18655),
            .I(N__18649));
    CascadeMux I__2880 (
            .O(N__18652),
            .I(N__18646));
    InMux I__2879 (
            .O(N__18649),
            .I(N__18643));
    InMux I__2878 (
            .O(N__18646),
            .I(N__18640));
    LocalMux I__2877 (
            .O(N__18643),
            .I(N__18635));
    LocalMux I__2876 (
            .O(N__18640),
            .I(N__18635));
    Span12Mux_s11_v I__2875 (
            .O(N__18635),
            .I(N__18632));
    Odrv12 I__2874 (
            .O(N__18632),
            .I(SYNTHESIZED_WIRE_12_6));
    InMux I__2873 (
            .O(N__18629),
            .I(N__18626));
    LocalMux I__2872 (
            .O(N__18626),
            .I(N__18623));
    Odrv4 I__2871 (
            .O(N__18623),
            .I(\b2v_inst.state_ns_0_i_a2_0_0_23 ));
    CascadeMux I__2870 (
            .O(N__18620),
            .I(\b2v_inst.state_ns_i_0_a2_11_o2_4_0_6_1_3_cascade_ ));
    InMux I__2869 (
            .O(N__18617),
            .I(N__18614));
    LocalMux I__2868 (
            .O(N__18614),
            .I(\b2v_inst.state_ns_i_0_a2_11_o2_4_0_1_3 ));
    InMux I__2867 (
            .O(N__18611),
            .I(N__18608));
    LocalMux I__2866 (
            .O(N__18608),
            .I(N__18605));
    Odrv12 I__2865 (
            .O(N__18605),
            .I(\b2v_inst.N_11 ));
    CascadeMux I__2864 (
            .O(N__18602),
            .I(\b2v_inst.N_4_i_i_1_cascade_ ));
    InMux I__2863 (
            .O(N__18599),
            .I(N__18596));
    LocalMux I__2862 (
            .O(N__18596),
            .I(\b2v_inst.g3_i_1 ));
    InMux I__2861 (
            .O(N__18593),
            .I(N__18590));
    LocalMux I__2860 (
            .O(N__18590),
            .I(N__18587));
    Span4Mux_v I__2859 (
            .O(N__18587),
            .I(N__18584));
    Sp12to4 I__2858 (
            .O(N__18584),
            .I(N__18581));
    Span12Mux_h I__2857 (
            .O(N__18581),
            .I(N__18578));
    Span12Mux_h I__2856 (
            .O(N__18578),
            .I(N__18575));
    Span12Mux_v I__2855 (
            .O(N__18575),
            .I(N__18572));
    Odrv12 I__2854 (
            .O(N__18572),
            .I(swit_c_8));
    InMux I__2853 (
            .O(N__18569),
            .I(N__18566));
    LocalMux I__2852 (
            .O(N__18566),
            .I(N__18563));
    Span12Mux_v I__2851 (
            .O(N__18563),
            .I(N__18560));
    Odrv12 I__2850 (
            .O(N__18560),
            .I(\b2v_inst.addr_ram_energia_m0_8 ));
    InMux I__2849 (
            .O(N__18557),
            .I(N__18554));
    LocalMux I__2848 (
            .O(N__18554),
            .I(\b2v_inst.state_ns_i_0_a2_11_o2_4_0_5_3 ));
    InMux I__2847 (
            .O(N__18551),
            .I(N__18548));
    LocalMux I__2846 (
            .O(N__18548),
            .I(\b2v_inst.state_RNO_2Z0Z_29 ));
    CascadeMux I__2845 (
            .O(N__18545),
            .I(\b2v_inst.state_ns_i_0_a2_11_o2_4_0_7_3_cascade_ ));
    InMux I__2844 (
            .O(N__18542),
            .I(N__18539));
    LocalMux I__2843 (
            .O(N__18539),
            .I(N__18536));
    Odrv4 I__2842 (
            .O(N__18536),
            .I(\b2v_inst.state_RNO_1Z0Z_29 ));
    InMux I__2841 (
            .O(N__18533),
            .I(N__18530));
    LocalMux I__2840 (
            .O(N__18530),
            .I(\b2v_inst.dir_energia_RNO_0Z0Z_0 ));
    CascadeMux I__2839 (
            .O(N__18527),
            .I(N__18524));
    InMux I__2838 (
            .O(N__18524),
            .I(N__18521));
    LocalMux I__2837 (
            .O(N__18521),
            .I(N__18518));
    Span4Mux_h I__2836 (
            .O(N__18518),
            .I(N__18515));
    Odrv4 I__2835 (
            .O(N__18515),
            .I(\b2v_inst.dir_mem_3Z0Z_5 ));
    CascadeMux I__2834 (
            .O(N__18512),
            .I(N__18509));
    InMux I__2833 (
            .O(N__18509),
            .I(N__18506));
    LocalMux I__2832 (
            .O(N__18506),
            .I(N__18503));
    Span4Mux_v I__2831 (
            .O(N__18503),
            .I(N__18500));
    Span4Mux_h I__2830 (
            .O(N__18500),
            .I(N__18497));
    Span4Mux_h I__2829 (
            .O(N__18497),
            .I(N__18494));
    Span4Mux_h I__2828 (
            .O(N__18494),
            .I(N__18491));
    Odrv4 I__2827 (
            .O(N__18491),
            .I(SYNTHESIZED_WIRE_1_5));
    InMux I__2826 (
            .O(N__18488),
            .I(N__18485));
    LocalMux I__2825 (
            .O(N__18485),
            .I(N__18482));
    Span4Mux_h I__2824 (
            .O(N__18482),
            .I(N__18479));
    Odrv4 I__2823 (
            .O(N__18479),
            .I(\b2v_inst.dir_memZ0Z_4 ));
    CascadeMux I__2822 (
            .O(N__18476),
            .I(\b2v_inst.addr_ram_iv_i_0_4_cascade_ ));
    CascadeMux I__2821 (
            .O(N__18473),
            .I(N__18470));
    CascadeBuf I__2820 (
            .O(N__18470),
            .I(N__18466));
    CascadeMux I__2819 (
            .O(N__18469),
            .I(N__18463));
    CascadeMux I__2818 (
            .O(N__18466),
            .I(N__18460));
    CascadeBuf I__2817 (
            .O(N__18463),
            .I(N__18457));
    CascadeBuf I__2816 (
            .O(N__18460),
            .I(N__18454));
    CascadeMux I__2815 (
            .O(N__18457),
            .I(N__18451));
    CascadeMux I__2814 (
            .O(N__18454),
            .I(N__18448));
    CascadeBuf I__2813 (
            .O(N__18451),
            .I(N__18445));
    CascadeBuf I__2812 (
            .O(N__18448),
            .I(N__18442));
    CascadeMux I__2811 (
            .O(N__18445),
            .I(N__18439));
    CascadeMux I__2810 (
            .O(N__18442),
            .I(N__18436));
    CascadeBuf I__2809 (
            .O(N__18439),
            .I(N__18433));
    CascadeBuf I__2808 (
            .O(N__18436),
            .I(N__18430));
    CascadeMux I__2807 (
            .O(N__18433),
            .I(N__18427));
    CascadeMux I__2806 (
            .O(N__18430),
            .I(N__18424));
    CascadeBuf I__2805 (
            .O(N__18427),
            .I(N__18421));
    CascadeBuf I__2804 (
            .O(N__18424),
            .I(N__18418));
    CascadeMux I__2803 (
            .O(N__18421),
            .I(N__18415));
    CascadeMux I__2802 (
            .O(N__18418),
            .I(N__18412));
    CascadeBuf I__2801 (
            .O(N__18415),
            .I(N__18409));
    InMux I__2800 (
            .O(N__18412),
            .I(N__18406));
    CascadeMux I__2799 (
            .O(N__18409),
            .I(N__18403));
    LocalMux I__2798 (
            .O(N__18406),
            .I(N__18400));
    InMux I__2797 (
            .O(N__18403),
            .I(N__18397));
    Span4Mux_h I__2796 (
            .O(N__18400),
            .I(N__18394));
    LocalMux I__2795 (
            .O(N__18397),
            .I(N__18391));
    Span4Mux_h I__2794 (
            .O(N__18394),
            .I(N__18388));
    Span12Mux_s11_h I__2793 (
            .O(N__18391),
            .I(N__18385));
    Span4Mux_h I__2792 (
            .O(N__18388),
            .I(N__18382));
    Odrv12 I__2791 (
            .O(N__18385),
            .I(indice_RNIN3333_4));
    Odrv4 I__2790 (
            .O(N__18382),
            .I(indice_RNIN3333_4));
    InMux I__2789 (
            .O(N__18377),
            .I(N__18374));
    LocalMux I__2788 (
            .O(N__18374),
            .I(N__18371));
    Odrv12 I__2787 (
            .O(N__18371),
            .I(\b2v_inst.dir_mem_1Z0Z_4 ));
    InMux I__2786 (
            .O(N__18368),
            .I(N__18365));
    LocalMux I__2785 (
            .O(N__18365),
            .I(\b2v_inst.addr_ram_iv_i_1_4 ));
    InMux I__2784 (
            .O(N__18362),
            .I(N__18358));
    InMux I__2783 (
            .O(N__18361),
            .I(N__18355));
    LocalMux I__2782 (
            .O(N__18358),
            .I(N__18352));
    LocalMux I__2781 (
            .O(N__18355),
            .I(N__18348));
    Span4Mux_v I__2780 (
            .O(N__18352),
            .I(N__18345));
    InMux I__2779 (
            .O(N__18351),
            .I(N__18342));
    Span4Mux_h I__2778 (
            .O(N__18348),
            .I(N__18335));
    Span4Mux_h I__2777 (
            .O(N__18345),
            .I(N__18335));
    LocalMux I__2776 (
            .O(N__18342),
            .I(N__18335));
    Odrv4 I__2775 (
            .O(N__18335),
            .I(\b2v_inst.un1_indice_cry_3_c_RNI23MGZ0 ));
    CascadeMux I__2774 (
            .O(N__18332),
            .I(N__18329));
    InMux I__2773 (
            .O(N__18329),
            .I(N__18326));
    LocalMux I__2772 (
            .O(N__18326),
            .I(N__18319));
    CascadeMux I__2771 (
            .O(N__18325),
            .I(N__18315));
    CascadeMux I__2770 (
            .O(N__18324),
            .I(N__18310));
    CascadeMux I__2769 (
            .O(N__18323),
            .I(N__18307));
    CascadeMux I__2768 (
            .O(N__18322),
            .I(N__18303));
    Span4Mux_h I__2767 (
            .O(N__18319),
            .I(N__18300));
    InMux I__2766 (
            .O(N__18318),
            .I(N__18295));
    InMux I__2765 (
            .O(N__18315),
            .I(N__18295));
    InMux I__2764 (
            .O(N__18314),
            .I(N__18288));
    InMux I__2763 (
            .O(N__18313),
            .I(N__18288));
    InMux I__2762 (
            .O(N__18310),
            .I(N__18288));
    InMux I__2761 (
            .O(N__18307),
            .I(N__18285));
    InMux I__2760 (
            .O(N__18306),
            .I(N__18280));
    InMux I__2759 (
            .O(N__18303),
            .I(N__18280));
    Odrv4 I__2758 (
            .O(N__18300),
            .I(\b2v_inst.dir_mem_316lto11_0 ));
    LocalMux I__2757 (
            .O(N__18295),
            .I(\b2v_inst.dir_mem_316lto11_0 ));
    LocalMux I__2756 (
            .O(N__18288),
            .I(\b2v_inst.dir_mem_316lto11_0 ));
    LocalMux I__2755 (
            .O(N__18285),
            .I(\b2v_inst.dir_mem_316lto11_0 ));
    LocalMux I__2754 (
            .O(N__18280),
            .I(\b2v_inst.dir_mem_316lto11_0 ));
    InMux I__2753 (
            .O(N__18269),
            .I(N__18266));
    LocalMux I__2752 (
            .O(N__18266),
            .I(N__18263));
    Span4Mux_v I__2751 (
            .O(N__18263),
            .I(N__18250));
    InMux I__2750 (
            .O(N__18262),
            .I(N__18247));
    InMux I__2749 (
            .O(N__18261),
            .I(N__18242));
    InMux I__2748 (
            .O(N__18260),
            .I(N__18242));
    InMux I__2747 (
            .O(N__18259),
            .I(N__18227));
    InMux I__2746 (
            .O(N__18258),
            .I(N__18227));
    InMux I__2745 (
            .O(N__18257),
            .I(N__18227));
    InMux I__2744 (
            .O(N__18256),
            .I(N__18227));
    InMux I__2743 (
            .O(N__18255),
            .I(N__18227));
    InMux I__2742 (
            .O(N__18254),
            .I(N__18227));
    InMux I__2741 (
            .O(N__18253),
            .I(N__18227));
    Odrv4 I__2740 (
            .O(N__18250),
            .I(\b2v_inst.dir_mem_316lt11 ));
    LocalMux I__2739 (
            .O(N__18247),
            .I(\b2v_inst.dir_mem_316lt11 ));
    LocalMux I__2738 (
            .O(N__18242),
            .I(\b2v_inst.dir_mem_316lt11 ));
    LocalMux I__2737 (
            .O(N__18227),
            .I(\b2v_inst.dir_mem_316lt11 ));
    CascadeMux I__2736 (
            .O(N__18218),
            .I(N__18215));
    InMux I__2735 (
            .O(N__18215),
            .I(N__18212));
    LocalMux I__2734 (
            .O(N__18212),
            .I(\b2v_inst.dir_mem_3Z0Z_4 ));
    CEMux I__2733 (
            .O(N__18209),
            .I(N__18205));
    CEMux I__2732 (
            .O(N__18208),
            .I(N__18200));
    LocalMux I__2731 (
            .O(N__18205),
            .I(N__18197));
    CEMux I__2730 (
            .O(N__18204),
            .I(N__18194));
    CEMux I__2729 (
            .O(N__18203),
            .I(N__18191));
    LocalMux I__2728 (
            .O(N__18200),
            .I(N__18188));
    Span4Mux_v I__2727 (
            .O(N__18197),
            .I(N__18183));
    LocalMux I__2726 (
            .O(N__18194),
            .I(N__18183));
    LocalMux I__2725 (
            .O(N__18191),
            .I(N__18180));
    Span4Mux_h I__2724 (
            .O(N__18188),
            .I(N__18177));
    Sp12to4 I__2723 (
            .O(N__18183),
            .I(N__18174));
    Odrv4 I__2722 (
            .O(N__18180),
            .I(\b2v_inst.N_362_i ));
    Odrv4 I__2721 (
            .O(N__18177),
            .I(\b2v_inst.N_362_i ));
    Odrv12 I__2720 (
            .O(N__18174),
            .I(\b2v_inst.N_362_i ));
    InMux I__2719 (
            .O(N__18167),
            .I(N__18161));
    InMux I__2718 (
            .O(N__18166),
            .I(N__18161));
    LocalMux I__2717 (
            .O(N__18161),
            .I(N__18158));
    Odrv12 I__2716 (
            .O(N__18158),
            .I(\b2v_inst.un8_dir_mem_1_cry_7_c_RNIIHVCZ0 ));
    CascadeMux I__2715 (
            .O(N__18155),
            .I(N__18152));
    InMux I__2714 (
            .O(N__18152),
            .I(N__18149));
    LocalMux I__2713 (
            .O(N__18149),
            .I(N__18146));
    Span4Mux_h I__2712 (
            .O(N__18146),
            .I(N__18143));
    Odrv4 I__2711 (
            .O(N__18143),
            .I(\b2v_inst.dir_mem_1_RNO_0Z0Z_8 ));
    InMux I__2710 (
            .O(N__18140),
            .I(N__18134));
    InMux I__2709 (
            .O(N__18139),
            .I(N__18134));
    LocalMux I__2708 (
            .O(N__18134),
            .I(N__18131));
    Odrv4 I__2707 (
            .O(N__18131),
            .I(\b2v_inst.un8_dir_mem_1_cry_8_c_RNIKK0DZ0 ));
    CascadeMux I__2706 (
            .O(N__18128),
            .I(N__18125));
    InMux I__2705 (
            .O(N__18125),
            .I(N__18122));
    LocalMux I__2704 (
            .O(N__18122),
            .I(N__18119));
    Span4Mux_h I__2703 (
            .O(N__18119),
            .I(N__18116));
    Odrv4 I__2702 (
            .O(N__18116),
            .I(\b2v_inst.dir_mem_1_RNO_0Z0Z_9 ));
    InMux I__2701 (
            .O(N__18113),
            .I(N__18109));
    InMux I__2700 (
            .O(N__18112),
            .I(N__18106));
    LocalMux I__2699 (
            .O(N__18109),
            .I(N__18103));
    LocalMux I__2698 (
            .O(N__18106),
            .I(N__18100));
    Span4Mux_v I__2697 (
            .O(N__18103),
            .I(N__18097));
    Span4Mux_v I__2696 (
            .O(N__18100),
            .I(N__18094));
    Odrv4 I__2695 (
            .O(N__18097),
            .I(\b2v_inst.un8_dir_mem_1_cry_4_c_RNIC8SCZ0 ));
    Odrv4 I__2694 (
            .O(N__18094),
            .I(\b2v_inst.un8_dir_mem_1_cry_4_c_RNIC8SCZ0 ));
    CascadeMux I__2693 (
            .O(N__18089),
            .I(N__18086));
    InMux I__2692 (
            .O(N__18086),
            .I(N__18083));
    LocalMux I__2691 (
            .O(N__18083),
            .I(N__18080));
    Span4Mux_h I__2690 (
            .O(N__18080),
            .I(N__18077));
    Odrv4 I__2689 (
            .O(N__18077),
            .I(\b2v_inst.dir_mem_1_RNO_0Z0Z_5 ));
    InMux I__2688 (
            .O(N__18074),
            .I(N__18071));
    LocalMux I__2687 (
            .O(N__18071),
            .I(N__18068));
    Odrv4 I__2686 (
            .O(N__18068),
            .I(\b2v_inst.dir_mem_1Z0Z_6 ));
    CascadeMux I__2685 (
            .O(N__18065),
            .I(N__18062));
    InMux I__2684 (
            .O(N__18062),
            .I(N__18059));
    LocalMux I__2683 (
            .O(N__18059),
            .I(N__18056));
    Span4Mux_v I__2682 (
            .O(N__18056),
            .I(N__18053));
    Odrv4 I__2681 (
            .O(N__18053),
            .I(\b2v_inst.dir_mem_3Z0Z_6 ));
    InMux I__2680 (
            .O(N__18050),
            .I(N__18047));
    LocalMux I__2679 (
            .O(N__18047),
            .I(N__18044));
    Odrv4 I__2678 (
            .O(N__18044),
            .I(\b2v_inst.dir_memZ0Z_7 ));
    CascadeMux I__2677 (
            .O(N__18041),
            .I(\b2v_inst.N_450_i_1_cascade_ ));
    InMux I__2676 (
            .O(N__18038),
            .I(N__18035));
    LocalMux I__2675 (
            .O(N__18035),
            .I(N__18032));
    Span4Mux_h I__2674 (
            .O(N__18032),
            .I(N__18029));
    Odrv4 I__2673 (
            .O(N__18029),
            .I(\b2v_inst.dir_memZ0Z_10 ));
    InMux I__2672 (
            .O(N__18026),
            .I(N__18023));
    LocalMux I__2671 (
            .O(N__18023),
            .I(N__18020));
    Odrv4 I__2670 (
            .O(N__18020),
            .I(\b2v_inst.dir_mem_1Z0Z_5 ));
    InMux I__2669 (
            .O(N__18017),
            .I(N__18014));
    LocalMux I__2668 (
            .O(N__18014),
            .I(N__18010));
    InMux I__2667 (
            .O(N__18013),
            .I(N__18007));
    Odrv4 I__2666 (
            .O(N__18010),
            .I(\b2v_inst.un8_dir_mem_1_cry_2_c_RNI82QCZ0 ));
    LocalMux I__2665 (
            .O(N__18007),
            .I(\b2v_inst.un8_dir_mem_1_cry_2_c_RNI82QCZ0 ));
    InMux I__2664 (
            .O(N__18002),
            .I(N__17999));
    LocalMux I__2663 (
            .O(N__17999),
            .I(N__17995));
    InMux I__2662 (
            .O(N__17998),
            .I(N__17992));
    Odrv4 I__2661 (
            .O(N__17995),
            .I(\b2v_inst.un8_dir_mem_1_cry_3_c_RNIA5RCZ0 ));
    LocalMux I__2660 (
            .O(N__17992),
            .I(\b2v_inst.un8_dir_mem_1_cry_3_c_RNIA5RCZ0 ));
    InMux I__2659 (
            .O(N__17987),
            .I(N__17983));
    InMux I__2658 (
            .O(N__17986),
            .I(N__17980));
    LocalMux I__2657 (
            .O(N__17983),
            .I(N__17977));
    LocalMux I__2656 (
            .O(N__17980),
            .I(N__17974));
    Span4Mux_h I__2655 (
            .O(N__17977),
            .I(N__17971));
    Odrv12 I__2654 (
            .O(N__17974),
            .I(\b2v_inst.un8_dir_mem_1_cry_5_c_RNIEBTCZ0 ));
    Odrv4 I__2653 (
            .O(N__17971),
            .I(\b2v_inst.un8_dir_mem_1_cry_5_c_RNIEBTCZ0 ));
    CascadeMux I__2652 (
            .O(N__17966),
            .I(N__17963));
    InMux I__2651 (
            .O(N__17963),
            .I(N__17960));
    LocalMux I__2650 (
            .O(N__17960),
            .I(N__17957));
    Sp12to4 I__2649 (
            .O(N__17957),
            .I(N__17954));
    Span12Mux_s10_v I__2648 (
            .O(N__17954),
            .I(N__17951));
    Odrv12 I__2647 (
            .O(N__17951),
            .I(\b2v_inst.dir_mem_1_RNO_0Z0Z_6 ));
    InMux I__2646 (
            .O(N__17948),
            .I(N__17945));
    LocalMux I__2645 (
            .O(N__17945),
            .I(\b2v_inst.dir_mem_215lt7 ));
    InMux I__2644 (
            .O(N__17942),
            .I(N__17939));
    LocalMux I__2643 (
            .O(N__17939),
            .I(\b2v_inst.dir_mem_115lt7 ));
    InMux I__2642 (
            .O(N__17936),
            .I(N__17933));
    LocalMux I__2641 (
            .O(N__17933),
            .I(N__17930));
    Span4Mux_h I__2640 (
            .O(N__17930),
            .I(N__17927));
    Odrv4 I__2639 (
            .O(N__17927),
            .I(\b2v_inst.dir_mem_1_RNO_0Z0Z_10 ));
    CascadeMux I__2638 (
            .O(N__17924),
            .I(\b2v_inst.dir_mem_115lt11_cascade_ ));
    CascadeMux I__2637 (
            .O(N__17921),
            .I(N__17917));
    InMux I__2636 (
            .O(N__17920),
            .I(N__17914));
    InMux I__2635 (
            .O(N__17917),
            .I(N__17911));
    LocalMux I__2634 (
            .O(N__17914),
            .I(N__17906));
    LocalMux I__2633 (
            .O(N__17911),
            .I(N__17906));
    Span4Mux_h I__2632 (
            .O(N__17906),
            .I(N__17903));
    Odrv4 I__2631 (
            .O(N__17903),
            .I(\b2v_inst.dir_mem_115lto7 ));
    CascadeMux I__2630 (
            .O(N__17900),
            .I(N__17897));
    InMux I__2629 (
            .O(N__17897),
            .I(N__17894));
    LocalMux I__2628 (
            .O(N__17894),
            .I(N__17891));
    Span4Mux_h I__2627 (
            .O(N__17891),
            .I(N__17888));
    Odrv4 I__2626 (
            .O(N__17888),
            .I(\b2v_inst.dir_mem_1_RNO_0Z0Z_7 ));
    CascadeMux I__2625 (
            .O(N__17885),
            .I(\b2v_inst.N_512_cascade_ ));
    InMux I__2624 (
            .O(N__17882),
            .I(N__17879));
    LocalMux I__2623 (
            .O(N__17879),
            .I(N__17876));
    Odrv4 I__2622 (
            .O(N__17876),
            .I(\b2v_inst.N_430_tz ));
    CascadeMux I__2621 (
            .O(N__17873),
            .I(\b2v_inst.g0_4_4_cascade_ ));
    InMux I__2620 (
            .O(N__17870),
            .I(N__17867));
    LocalMux I__2619 (
            .O(N__17867),
            .I(N__17864));
    Odrv12 I__2618 (
            .O(N__17864),
            .I(\b2v_inst.g3_0_0 ));
    CascadeMux I__2617 (
            .O(N__17861),
            .I(N__17858));
    InMux I__2616 (
            .O(N__17858),
            .I(N__17854));
    InMux I__2615 (
            .O(N__17857),
            .I(N__17851));
    LocalMux I__2614 (
            .O(N__17854),
            .I(N__17848));
    LocalMux I__2613 (
            .O(N__17851),
            .I(N__17843));
    Span4Mux_v I__2612 (
            .O(N__17848),
            .I(N__17843));
    Odrv4 I__2611 (
            .O(N__17843),
            .I(\b2v_inst.un4_pix_count_intlto18Z0Z_0 ));
    CascadeMux I__2610 (
            .O(N__17840),
            .I(\b2v_inst.g0_0_cascade_ ));
    InMux I__2609 (
            .O(N__17837),
            .I(N__17834));
    LocalMux I__2608 (
            .O(N__17834),
            .I(\b2v_inst.g3_0 ));
    InMux I__2607 (
            .O(N__17831),
            .I(N__17828));
    LocalMux I__2606 (
            .O(N__17828),
            .I(\b2v_inst.g0_4_5 ));
    IoInMux I__2605 (
            .O(N__17825),
            .I(N__17822));
    LocalMux I__2604 (
            .O(N__17822),
            .I(N__17818));
    InMux I__2603 (
            .O(N__17821),
            .I(N__17815));
    Span4Mux_s3_h I__2602 (
            .O(N__17818),
            .I(N__17812));
    LocalMux I__2601 (
            .O(N__17815),
            .I(N__17809));
    Span4Mux_h I__2600 (
            .O(N__17812),
            .I(N__17806));
    Span4Mux_h I__2599 (
            .O(N__17809),
            .I(N__17803));
    Span4Mux_v I__2598 (
            .O(N__17806),
            .I(N__17798));
    Span4Mux_h I__2597 (
            .O(N__17803),
            .I(N__17798));
    Odrv4 I__2596 (
            .O(N__17798),
            .I(leds_c_10));
    IoInMux I__2595 (
            .O(N__17795),
            .I(N__17792));
    LocalMux I__2594 (
            .O(N__17792),
            .I(N__17789));
    IoSpan4Mux I__2593 (
            .O(N__17789),
            .I(N__17786));
    Span4Mux_s2_v I__2592 (
            .O(N__17786),
            .I(N__17783));
    Span4Mux_h I__2591 (
            .O(N__17783),
            .I(N__17779));
    InMux I__2590 (
            .O(N__17782),
            .I(N__17776));
    Span4Mux_v I__2589 (
            .O(N__17779),
            .I(N__17773));
    LocalMux I__2588 (
            .O(N__17776),
            .I(N__17770));
    Odrv4 I__2587 (
            .O(N__17773),
            .I(leds_c_11));
    Odrv12 I__2586 (
            .O(N__17770),
            .I(leds_c_11));
    InMux I__2585 (
            .O(N__17765),
            .I(N__17761));
    IoInMux I__2584 (
            .O(N__17764),
            .I(N__17758));
    LocalMux I__2583 (
            .O(N__17761),
            .I(N__17755));
    LocalMux I__2582 (
            .O(N__17758),
            .I(N__17752));
    Span4Mux_h I__2581 (
            .O(N__17755),
            .I(N__17749));
    Span12Mux_s7_h I__2580 (
            .O(N__17752),
            .I(N__17746));
    Span4Mux_v I__2579 (
            .O(N__17749),
            .I(N__17743));
    Odrv12 I__2578 (
            .O(N__17746),
            .I(leds_c_7));
    Odrv4 I__2577 (
            .O(N__17743),
            .I(leds_c_7));
    InMux I__2576 (
            .O(N__17738),
            .I(N__17735));
    LocalMux I__2575 (
            .O(N__17735),
            .I(\b2v_inst.G_40_i_3 ));
    InMux I__2574 (
            .O(N__17732),
            .I(N__17724));
    InMux I__2573 (
            .O(N__17731),
            .I(N__17715));
    InMux I__2572 (
            .O(N__17730),
            .I(N__17715));
    InMux I__2571 (
            .O(N__17729),
            .I(N__17715));
    InMux I__2570 (
            .O(N__17728),
            .I(N__17710));
    CascadeMux I__2569 (
            .O(N__17727),
            .I(N__17706));
    LocalMux I__2568 (
            .O(N__17724),
            .I(N__17702));
    CascadeMux I__2567 (
            .O(N__17723),
            .I(N__17699));
    InMux I__2566 (
            .O(N__17722),
            .I(N__17696));
    LocalMux I__2565 (
            .O(N__17715),
            .I(N__17692));
    InMux I__2564 (
            .O(N__17714),
            .I(N__17689));
    InMux I__2563 (
            .O(N__17713),
            .I(N__17686));
    LocalMux I__2562 (
            .O(N__17710),
            .I(N__17682));
    InMux I__2561 (
            .O(N__17709),
            .I(N__17677));
    InMux I__2560 (
            .O(N__17706),
            .I(N__17677));
    InMux I__2559 (
            .O(N__17705),
            .I(N__17674));
    Span4Mux_v I__2558 (
            .O(N__17702),
            .I(N__17671));
    InMux I__2557 (
            .O(N__17699),
            .I(N__17668));
    LocalMux I__2556 (
            .O(N__17696),
            .I(N__17665));
    InMux I__2555 (
            .O(N__17695),
            .I(N__17662));
    Span4Mux_h I__2554 (
            .O(N__17692),
            .I(N__17659));
    LocalMux I__2553 (
            .O(N__17689),
            .I(N__17656));
    LocalMux I__2552 (
            .O(N__17686),
            .I(N__17653));
    InMux I__2551 (
            .O(N__17685),
            .I(N__17650));
    Span4Mux_h I__2550 (
            .O(N__17682),
            .I(N__17645));
    LocalMux I__2549 (
            .O(N__17677),
            .I(N__17645));
    LocalMux I__2548 (
            .O(N__17674),
            .I(N__17636));
    Span4Mux_h I__2547 (
            .O(N__17671),
            .I(N__17636));
    LocalMux I__2546 (
            .O(N__17668),
            .I(N__17636));
    Span4Mux_v I__2545 (
            .O(N__17665),
            .I(N__17636));
    LocalMux I__2544 (
            .O(N__17662),
            .I(SYNTHESIZED_WIRE_4_19));
    Odrv4 I__2543 (
            .O(N__17659),
            .I(SYNTHESIZED_WIRE_4_19));
    Odrv4 I__2542 (
            .O(N__17656),
            .I(SYNTHESIZED_WIRE_4_19));
    Odrv4 I__2541 (
            .O(N__17653),
            .I(SYNTHESIZED_WIRE_4_19));
    LocalMux I__2540 (
            .O(N__17650),
            .I(SYNTHESIZED_WIRE_4_19));
    Odrv4 I__2539 (
            .O(N__17645),
            .I(SYNTHESIZED_WIRE_4_19));
    Odrv4 I__2538 (
            .O(N__17636),
            .I(SYNTHESIZED_WIRE_4_19));
    InMux I__2537 (
            .O(N__17621),
            .I(N__17617));
    InMux I__2536 (
            .O(N__17620),
            .I(N__17614));
    LocalMux I__2535 (
            .O(N__17617),
            .I(N__17605));
    LocalMux I__2534 (
            .O(N__17614),
            .I(N__17605));
    InMux I__2533 (
            .O(N__17613),
            .I(N__17602));
    InMux I__2532 (
            .O(N__17612),
            .I(N__17599));
    InMux I__2531 (
            .O(N__17611),
            .I(N__17595));
    InMux I__2530 (
            .O(N__17610),
            .I(N__17589));
    Span4Mux_v I__2529 (
            .O(N__17605),
            .I(N__17584));
    LocalMux I__2528 (
            .O(N__17602),
            .I(N__17584));
    LocalMux I__2527 (
            .O(N__17599),
            .I(N__17581));
    InMux I__2526 (
            .O(N__17598),
            .I(N__17578));
    LocalMux I__2525 (
            .O(N__17595),
            .I(N__17575));
    InMux I__2524 (
            .O(N__17594),
            .I(N__17572));
    InMux I__2523 (
            .O(N__17593),
            .I(N__17569));
    InMux I__2522 (
            .O(N__17592),
            .I(N__17566));
    LocalMux I__2521 (
            .O(N__17589),
            .I(N__17562));
    Span4Mux_h I__2520 (
            .O(N__17584),
            .I(N__17559));
    Span4Mux_h I__2519 (
            .O(N__17581),
            .I(N__17552));
    LocalMux I__2518 (
            .O(N__17578),
            .I(N__17552));
    Span4Mux_v I__2517 (
            .O(N__17575),
            .I(N__17552));
    LocalMux I__2516 (
            .O(N__17572),
            .I(N__17549));
    LocalMux I__2515 (
            .O(N__17569),
            .I(N__17544));
    LocalMux I__2514 (
            .O(N__17566),
            .I(N__17544));
    InMux I__2513 (
            .O(N__17565),
            .I(N__17541));
    Span4Mux_h I__2512 (
            .O(N__17562),
            .I(N__17538));
    Odrv4 I__2511 (
            .O(N__17559),
            .I(SYNTHESIZED_WIRE_4_16));
    Odrv4 I__2510 (
            .O(N__17552),
            .I(SYNTHESIZED_WIRE_4_16));
    Odrv4 I__2509 (
            .O(N__17549),
            .I(SYNTHESIZED_WIRE_4_16));
    Odrv4 I__2508 (
            .O(N__17544),
            .I(SYNTHESIZED_WIRE_4_16));
    LocalMux I__2507 (
            .O(N__17541),
            .I(SYNTHESIZED_WIRE_4_16));
    Odrv4 I__2506 (
            .O(N__17538),
            .I(SYNTHESIZED_WIRE_4_16));
    InMux I__2505 (
            .O(N__17525),
            .I(N__17521));
    InMux I__2504 (
            .O(N__17524),
            .I(N__17518));
    LocalMux I__2503 (
            .O(N__17521),
            .I(\b2v_inst.N_5 ));
    LocalMux I__2502 (
            .O(N__17518),
            .I(\b2v_inst.N_5 ));
    CascadeMux I__2501 (
            .O(N__17513),
            .I(\b2v_inst.N_430_i_1_cascade_ ));
    InMux I__2500 (
            .O(N__17510),
            .I(N__17506));
    InMux I__2499 (
            .O(N__17509),
            .I(N__17503));
    LocalMux I__2498 (
            .O(N__17506),
            .I(N__17497));
    LocalMux I__2497 (
            .O(N__17503),
            .I(N__17494));
    InMux I__2496 (
            .O(N__17502),
            .I(N__17491));
    InMux I__2495 (
            .O(N__17501),
            .I(N__17485));
    InMux I__2494 (
            .O(N__17500),
            .I(N__17485));
    Span4Mux_v I__2493 (
            .O(N__17497),
            .I(N__17476));
    Span4Mux_v I__2492 (
            .O(N__17494),
            .I(N__17476));
    LocalMux I__2491 (
            .O(N__17491),
            .I(N__17476));
    InMux I__2490 (
            .O(N__17490),
            .I(N__17473));
    LocalMux I__2489 (
            .O(N__17485),
            .I(N__17470));
    InMux I__2488 (
            .O(N__17484),
            .I(N__17467));
    InMux I__2487 (
            .O(N__17483),
            .I(N__17464));
    Span4Mux_h I__2486 (
            .O(N__17476),
            .I(N__17461));
    LocalMux I__2485 (
            .O(N__17473),
            .I(N__17456));
    Span4Mux_v I__2484 (
            .O(N__17470),
            .I(N__17456));
    LocalMux I__2483 (
            .O(N__17467),
            .I(SYNTHESIZED_WIRE_4_18));
    LocalMux I__2482 (
            .O(N__17464),
            .I(SYNTHESIZED_WIRE_4_18));
    Odrv4 I__2481 (
            .O(N__17461),
            .I(SYNTHESIZED_WIRE_4_18));
    Odrv4 I__2480 (
            .O(N__17456),
            .I(SYNTHESIZED_WIRE_4_18));
    InMux I__2479 (
            .O(N__17447),
            .I(N__17441));
    InMux I__2478 (
            .O(N__17446),
            .I(N__17438));
    InMux I__2477 (
            .O(N__17445),
            .I(N__17433));
    InMux I__2476 (
            .O(N__17444),
            .I(N__17428));
    LocalMux I__2475 (
            .O(N__17441),
            .I(N__17423));
    LocalMux I__2474 (
            .O(N__17438),
            .I(N__17423));
    InMux I__2473 (
            .O(N__17437),
            .I(N__17420));
    InMux I__2472 (
            .O(N__17436),
            .I(N__17417));
    LocalMux I__2471 (
            .O(N__17433),
            .I(N__17414));
    InMux I__2470 (
            .O(N__17432),
            .I(N__17411));
    InMux I__2469 (
            .O(N__17431),
            .I(N__17408));
    LocalMux I__2468 (
            .O(N__17428),
            .I(N__17405));
    Span4Mux_v I__2467 (
            .O(N__17423),
            .I(N__17402));
    LocalMux I__2466 (
            .O(N__17420),
            .I(N__17397));
    LocalMux I__2465 (
            .O(N__17417),
            .I(N__17397));
    Span4Mux_h I__2464 (
            .O(N__17414),
            .I(N__17394));
    LocalMux I__2463 (
            .O(N__17411),
            .I(SYNTHESIZED_WIRE_4_17));
    LocalMux I__2462 (
            .O(N__17408),
            .I(SYNTHESIZED_WIRE_4_17));
    Odrv4 I__2461 (
            .O(N__17405),
            .I(SYNTHESIZED_WIRE_4_17));
    Odrv4 I__2460 (
            .O(N__17402),
            .I(SYNTHESIZED_WIRE_4_17));
    Odrv4 I__2459 (
            .O(N__17397),
            .I(SYNTHESIZED_WIRE_4_17));
    Odrv4 I__2458 (
            .O(N__17394),
            .I(SYNTHESIZED_WIRE_4_17));
    CascadeMux I__2457 (
            .O(N__17381),
            .I(N__17377));
    CascadeMux I__2456 (
            .O(N__17380),
            .I(N__17373));
    InMux I__2455 (
            .O(N__17377),
            .I(N__17370));
    InMux I__2454 (
            .O(N__17376),
            .I(N__17365));
    InMux I__2453 (
            .O(N__17373),
            .I(N__17365));
    LocalMux I__2452 (
            .O(N__17370),
            .I(\b2v_inst.g1Z0Z_0 ));
    LocalMux I__2451 (
            .O(N__17365),
            .I(\b2v_inst.g1Z0Z_0 ));
    InMux I__2450 (
            .O(N__17360),
            .I(N__17357));
    LocalMux I__2449 (
            .O(N__17357),
            .I(\b2v_inst.pix_count_anterior5 ));
    CascadeMux I__2448 (
            .O(N__17354),
            .I(\b2v_inst.state_ns_0_i_o2_6_23_cascade_ ));
    InMux I__2447 (
            .O(N__17351),
            .I(N__17348));
    LocalMux I__2446 (
            .O(N__17348),
            .I(\b2v_inst.state_ns_0_i_o2_7_23 ));
    CascadeMux I__2445 (
            .O(N__17345),
            .I(\b2v_inst.g0_6_cascade_ ));
    InMux I__2444 (
            .O(N__17342),
            .I(N__17339));
    LocalMux I__2443 (
            .O(N__17339),
            .I(\b2v_inst.o2 ));
    CascadeMux I__2442 (
            .O(N__17336),
            .I(\b2v_inst.G_40_i_6_cascade_ ));
    InMux I__2441 (
            .O(N__17333),
            .I(N__17330));
    LocalMux I__2440 (
            .O(N__17330),
            .I(\b2v_inst.state_ns_i_0_a2_11_a2_0_3_3 ));
    InMux I__2439 (
            .O(N__17327),
            .I(N__17324));
    LocalMux I__2438 (
            .O(N__17324),
            .I(\b2v_inst.N_618_5 ));
    InMux I__2437 (
            .O(N__17321),
            .I(N__17318));
    LocalMux I__2436 (
            .O(N__17318),
            .I(N__17315));
    Span4Mux_h I__2435 (
            .O(N__17315),
            .I(N__17311));
    InMux I__2434 (
            .O(N__17314),
            .I(N__17308));
    Odrv4 I__2433 (
            .O(N__17311),
            .I(\b2v_inst1.N_49 ));
    LocalMux I__2432 (
            .O(N__17308),
            .I(\b2v_inst1.N_49 ));
    InMux I__2431 (
            .O(N__17303),
            .I(N__17294));
    InMux I__2430 (
            .O(N__17302),
            .I(N__17294));
    InMux I__2429 (
            .O(N__17301),
            .I(N__17291));
    InMux I__2428 (
            .O(N__17300),
            .I(N__17286));
    InMux I__2427 (
            .O(N__17299),
            .I(N__17282));
    LocalMux I__2426 (
            .O(N__17294),
            .I(N__17279));
    LocalMux I__2425 (
            .O(N__17291),
            .I(N__17276));
    InMux I__2424 (
            .O(N__17290),
            .I(N__17273));
    InMux I__2423 (
            .O(N__17289),
            .I(N__17270));
    LocalMux I__2422 (
            .O(N__17286),
            .I(N__17267));
    InMux I__2421 (
            .O(N__17285),
            .I(N__17264));
    LocalMux I__2420 (
            .O(N__17282),
            .I(N__17261));
    Span4Mux_v I__2419 (
            .O(N__17279),
            .I(N__17254));
    Span4Mux_v I__2418 (
            .O(N__17276),
            .I(N__17254));
    LocalMux I__2417 (
            .O(N__17273),
            .I(N__17254));
    LocalMux I__2416 (
            .O(N__17270),
            .I(N__17247));
    Span4Mux_h I__2415 (
            .O(N__17267),
            .I(N__17247));
    LocalMux I__2414 (
            .O(N__17264),
            .I(N__17247));
    Span4Mux_v I__2413 (
            .O(N__17261),
            .I(N__17242));
    Span4Mux_h I__2412 (
            .O(N__17254),
            .I(N__17242));
    Span4Mux_v I__2411 (
            .O(N__17247),
            .I(N__17239));
    Odrv4 I__2410 (
            .O(N__17242),
            .I(\b2v_inst1.r_RX_Byte_1_sqmuxa ));
    Odrv4 I__2409 (
            .O(N__17239),
            .I(\b2v_inst1.r_RX_Byte_1_sqmuxa ));
    InMux I__2408 (
            .O(N__17234),
            .I(N__17231));
    LocalMux I__2407 (
            .O(N__17231),
            .I(\b2v_inst.N_618_3 ));
    InMux I__2406 (
            .O(N__17228),
            .I(N__17225));
    LocalMux I__2405 (
            .O(N__17225),
            .I(\b2v_inst.state_ns_i_0_a2_11_o2_4_0_3_3 ));
    CascadeMux I__2404 (
            .O(N__17222),
            .I(N__17218));
    InMux I__2403 (
            .O(N__17221),
            .I(N__17214));
    InMux I__2402 (
            .O(N__17218),
            .I(N__17209));
    InMux I__2401 (
            .O(N__17217),
            .I(N__17209));
    LocalMux I__2400 (
            .O(N__17214),
            .I(N__17206));
    LocalMux I__2399 (
            .O(N__17209),
            .I(\b2v_inst.un4_pix_count_intlto19_0_0 ));
    Odrv12 I__2398 (
            .O(N__17206),
            .I(\b2v_inst.un4_pix_count_intlto19_0_0 ));
    CascadeMux I__2397 (
            .O(N__17201),
            .I(N__17198));
    InMux I__2396 (
            .O(N__17198),
            .I(N__17195));
    LocalMux I__2395 (
            .O(N__17195),
            .I(\b2v_inst.G_40_i_2 ));
    IoInMux I__2394 (
            .O(N__17192),
            .I(N__17189));
    LocalMux I__2393 (
            .O(N__17189),
            .I(N__17186));
    IoSpan4Mux I__2392 (
            .O(N__17186),
            .I(N__17182));
    InMux I__2391 (
            .O(N__17185),
            .I(N__17179));
    Span4Mux_s3_v I__2390 (
            .O(N__17182),
            .I(N__17176));
    LocalMux I__2389 (
            .O(N__17179),
            .I(N__17173));
    Span4Mux_v I__2388 (
            .O(N__17176),
            .I(N__17170));
    Span4Mux_v I__2387 (
            .O(N__17173),
            .I(N__17167));
    Span4Mux_v I__2386 (
            .O(N__17170),
            .I(N__17164));
    Span4Mux_h I__2385 (
            .O(N__17167),
            .I(N__17161));
    Odrv4 I__2384 (
            .O(N__17164),
            .I(leds_c_4));
    Odrv4 I__2383 (
            .O(N__17161),
            .I(leds_c_4));
    IoInMux I__2382 (
            .O(N__17156),
            .I(N__17153));
    LocalMux I__2381 (
            .O(N__17153),
            .I(N__17150));
    Span4Mux_s3_v I__2380 (
            .O(N__17150),
            .I(N__17146));
    InMux I__2379 (
            .O(N__17149),
            .I(N__17143));
    Sp12to4 I__2378 (
            .O(N__17146),
            .I(N__17140));
    LocalMux I__2377 (
            .O(N__17143),
            .I(N__17137));
    Span12Mux_s11_h I__2376 (
            .O(N__17140),
            .I(N__17134));
    Span4Mux_h I__2375 (
            .O(N__17137),
            .I(N__17131));
    Span12Mux_v I__2374 (
            .O(N__17134),
            .I(N__17128));
    Span4Mux_v I__2373 (
            .O(N__17131),
            .I(N__17125));
    Odrv12 I__2372 (
            .O(N__17128),
            .I(leds_c_5));
    Odrv4 I__2371 (
            .O(N__17125),
            .I(leds_c_5));
    InMux I__2370 (
            .O(N__17120),
            .I(N__17117));
    LocalMux I__2369 (
            .O(N__17117),
            .I(\b2v_inst.dir_mem_115lt6_0 ));
    CascadeMux I__2368 (
            .O(N__17114),
            .I(\b2v_inst.g0_1_0_cascade_ ));
    InMux I__2367 (
            .O(N__17111),
            .I(N__17108));
    LocalMux I__2366 (
            .O(N__17108),
            .I(N__17105));
    Span4Mux_h I__2365 (
            .O(N__17105),
            .I(N__17101));
    InMux I__2364 (
            .O(N__17104),
            .I(N__17098));
    Span4Mux_h I__2363 (
            .O(N__17101),
            .I(N__17095));
    LocalMux I__2362 (
            .O(N__17098),
            .I(N__17092));
    Odrv4 I__2361 (
            .O(N__17095),
            .I(\b2v_inst.un7_pix_count_int_0_N_2_THRU_CO ));
    Odrv12 I__2360 (
            .O(N__17092),
            .I(\b2v_inst.un7_pix_count_int_0_N_2_THRU_CO ));
    InMux I__2359 (
            .O(N__17087),
            .I(\b2v_inst.un8_dir_mem_2_cry_4 ));
    InMux I__2358 (
            .O(N__17084),
            .I(\b2v_inst.un8_dir_mem_2_cry_5 ));
    InMux I__2357 (
            .O(N__17081),
            .I(\b2v_inst.un8_dir_mem_2_cry_6 ));
    InMux I__2356 (
            .O(N__17078),
            .I(\b2v_inst.un8_dir_mem_2_cry_7 ));
    InMux I__2355 (
            .O(N__17075),
            .I(bfn_9_6_0_));
    InMux I__2354 (
            .O(N__17072),
            .I(\b2v_inst.un8_dir_mem_2_cry_9 ));
    InMux I__2353 (
            .O(N__17069),
            .I(N__17066));
    LocalMux I__2352 (
            .O(N__17066),
            .I(\b2v_inst.dir_mem_215lt6_0 ));
    CascadeMux I__2351 (
            .O(N__17063),
            .I(\b2v_inst1.N_36_cascade_ ));
    CascadeMux I__2350 (
            .O(N__17060),
            .I(N__17057));
    InMux I__2349 (
            .O(N__17057),
            .I(N__17049));
    InMux I__2348 (
            .O(N__17056),
            .I(N__17049));
    CascadeMux I__2347 (
            .O(N__17055),
            .I(N__17043));
    InMux I__2346 (
            .O(N__17054),
            .I(N__17038));
    LocalMux I__2345 (
            .O(N__17049),
            .I(N__17035));
    InMux I__2344 (
            .O(N__17048),
            .I(N__17028));
    InMux I__2343 (
            .O(N__17047),
            .I(N__17028));
    InMux I__2342 (
            .O(N__17046),
            .I(N__17028));
    InMux I__2341 (
            .O(N__17043),
            .I(N__17021));
    InMux I__2340 (
            .O(N__17042),
            .I(N__17021));
    InMux I__2339 (
            .O(N__17041),
            .I(N__17021));
    LocalMux I__2338 (
            .O(N__17038),
            .I(\b2v_inst1.r_Bit_IndexZ0Z_1 ));
    Odrv12 I__2337 (
            .O(N__17035),
            .I(\b2v_inst1.r_Bit_IndexZ0Z_1 ));
    LocalMux I__2336 (
            .O(N__17028),
            .I(\b2v_inst1.r_Bit_IndexZ0Z_1 ));
    LocalMux I__2335 (
            .O(N__17021),
            .I(\b2v_inst1.r_Bit_IndexZ0Z_1 ));
    InMux I__2334 (
            .O(N__17012),
            .I(N__17006));
    InMux I__2333 (
            .O(N__17011),
            .I(N__17001));
    InMux I__2332 (
            .O(N__17010),
            .I(N__17001));
    InMux I__2331 (
            .O(N__17009),
            .I(N__16992));
    LocalMux I__2330 (
            .O(N__17006),
            .I(N__16987));
    LocalMux I__2329 (
            .O(N__17001),
            .I(N__16987));
    InMux I__2328 (
            .O(N__17000),
            .I(N__16982));
    InMux I__2327 (
            .O(N__16999),
            .I(N__16982));
    InMux I__2326 (
            .O(N__16998),
            .I(N__16973));
    InMux I__2325 (
            .O(N__16997),
            .I(N__16973));
    InMux I__2324 (
            .O(N__16996),
            .I(N__16973));
    InMux I__2323 (
            .O(N__16995),
            .I(N__16973));
    LocalMux I__2322 (
            .O(N__16992),
            .I(\b2v_inst1.r_Bit_IndexZ0Z_0 ));
    Odrv4 I__2321 (
            .O(N__16987),
            .I(\b2v_inst1.r_Bit_IndexZ0Z_0 ));
    LocalMux I__2320 (
            .O(N__16982),
            .I(\b2v_inst1.r_Bit_IndexZ0Z_0 ));
    LocalMux I__2319 (
            .O(N__16973),
            .I(\b2v_inst1.r_Bit_IndexZ0Z_0 ));
    InMux I__2318 (
            .O(N__16964),
            .I(N__16961));
    LocalMux I__2317 (
            .O(N__16961),
            .I(\b2v_inst1.N_50 ));
    CascadeMux I__2316 (
            .O(N__16958),
            .I(N__16955));
    InMux I__2315 (
            .O(N__16955),
            .I(N__16952));
    LocalMux I__2314 (
            .O(N__16952),
            .I(\b2v_inst1.r_RX_Bytece_0_5 ));
    InMux I__2313 (
            .O(N__16949),
            .I(N__16946));
    LocalMux I__2312 (
            .O(N__16946),
            .I(N__16943));
    Odrv12 I__2311 (
            .O(N__16943),
            .I(N_460_i));
    InMux I__2310 (
            .O(N__16940),
            .I(N__16937));
    LocalMux I__2309 (
            .O(N__16937),
            .I(N__16934));
    Span4Mux_v I__2308 (
            .O(N__16934),
            .I(N__16931));
    Odrv4 I__2307 (
            .O(N__16931),
            .I(N_459_i));
    InMux I__2306 (
            .O(N__16928),
            .I(\b2v_inst.un8_dir_mem_2_cry_1 ));
    InMux I__2305 (
            .O(N__16925),
            .I(\b2v_inst.un8_dir_mem_2_cry_2 ));
    InMux I__2304 (
            .O(N__16922),
            .I(\b2v_inst.un8_dir_mem_2_cry_3 ));
    InMux I__2303 (
            .O(N__16919),
            .I(N__16916));
    LocalMux I__2302 (
            .O(N__16916),
            .I(\b2v_inst1.r_RX_Bytece_0_6 ));
    CascadeMux I__2301 (
            .O(N__16913),
            .I(N__16910));
    InMux I__2300 (
            .O(N__16910),
            .I(N__16907));
    LocalMux I__2299 (
            .O(N__16907),
            .I(N__16898));
    InMux I__2298 (
            .O(N__16906),
            .I(N__16893));
    InMux I__2297 (
            .O(N__16905),
            .I(N__16893));
    InMux I__2296 (
            .O(N__16904),
            .I(N__16890));
    InMux I__2295 (
            .O(N__16903),
            .I(N__16887));
    InMux I__2294 (
            .O(N__16902),
            .I(N__16882));
    InMux I__2293 (
            .O(N__16901),
            .I(N__16882));
    Span4Mux_h I__2292 (
            .O(N__16898),
            .I(N__16879));
    LocalMux I__2291 (
            .O(N__16893),
            .I(N__16876));
    LocalMux I__2290 (
            .O(N__16890),
            .I(\b2v_inst1.r_Clk_CountZ0Z_2 ));
    LocalMux I__2289 (
            .O(N__16887),
            .I(\b2v_inst1.r_Clk_CountZ0Z_2 ));
    LocalMux I__2288 (
            .O(N__16882),
            .I(\b2v_inst1.r_Clk_CountZ0Z_2 ));
    Odrv4 I__2287 (
            .O(N__16879),
            .I(\b2v_inst1.r_Clk_CountZ0Z_2 ));
    Odrv4 I__2286 (
            .O(N__16876),
            .I(\b2v_inst1.r_Clk_CountZ0Z_2 ));
    CascadeMux I__2285 (
            .O(N__16865),
            .I(\b2v_inst1.m16_0_o2_cascade_ ));
    InMux I__2284 (
            .O(N__16862),
            .I(N__16859));
    LocalMux I__2283 (
            .O(N__16859),
            .I(N__16856));
    Odrv4 I__2282 (
            .O(N__16856),
            .I(\b2v_inst.g0_1_0_0 ));
    InMux I__2281 (
            .O(N__16853),
            .I(N__16849));
    CascadeMux I__2280 (
            .O(N__16852),
            .I(N__16844));
    LocalMux I__2279 (
            .O(N__16849),
            .I(N__16839));
    InMux I__2278 (
            .O(N__16848),
            .I(N__16836));
    InMux I__2277 (
            .O(N__16847),
            .I(N__16833));
    InMux I__2276 (
            .O(N__16844),
            .I(N__16828));
    InMux I__2275 (
            .O(N__16843),
            .I(N__16828));
    InMux I__2274 (
            .O(N__16842),
            .I(N__16825));
    Span4Mux_v I__2273 (
            .O(N__16839),
            .I(N__16816));
    LocalMux I__2272 (
            .O(N__16836),
            .I(N__16816));
    LocalMux I__2271 (
            .O(N__16833),
            .I(N__16813));
    LocalMux I__2270 (
            .O(N__16828),
            .I(N__16810));
    LocalMux I__2269 (
            .O(N__16825),
            .I(N__16807));
    InMux I__2268 (
            .O(N__16824),
            .I(N__16800));
    InMux I__2267 (
            .O(N__16823),
            .I(N__16800));
    InMux I__2266 (
            .O(N__16822),
            .I(N__16800));
    InMux I__2265 (
            .O(N__16821),
            .I(N__16797));
    Span4Mux_h I__2264 (
            .O(N__16816),
            .I(N__16794));
    Span4Mux_v I__2263 (
            .O(N__16813),
            .I(N__16789));
    Span4Mux_v I__2262 (
            .O(N__16810),
            .I(N__16789));
    Span4Mux_h I__2261 (
            .O(N__16807),
            .I(N__16784));
    LocalMux I__2260 (
            .O(N__16800),
            .I(N__16784));
    LocalMux I__2259 (
            .O(N__16797),
            .I(SYNTHESIZED_WIRE_4_7));
    Odrv4 I__2258 (
            .O(N__16794),
            .I(SYNTHESIZED_WIRE_4_7));
    Odrv4 I__2257 (
            .O(N__16789),
            .I(SYNTHESIZED_WIRE_4_7));
    Odrv4 I__2256 (
            .O(N__16784),
            .I(SYNTHESIZED_WIRE_4_7));
    CascadeMux I__2255 (
            .O(N__16775),
            .I(N__16772));
    InMux I__2254 (
            .O(N__16772),
            .I(N__16769));
    LocalMux I__2253 (
            .O(N__16769),
            .I(N__16766));
    Span4Mux_v I__2252 (
            .O(N__16766),
            .I(N__16763));
    Span4Mux_h I__2251 (
            .O(N__16763),
            .I(N__16760));
    Odrv4 I__2250 (
            .O(N__16760),
            .I(\b2v_inst.un4_pix_count_intlto6_d_1_2 ));
    InMux I__2249 (
            .O(N__16757),
            .I(N__16753));
    InMux I__2248 (
            .O(N__16756),
            .I(N__16749));
    LocalMux I__2247 (
            .O(N__16753),
            .I(N__16741));
    InMux I__2246 (
            .O(N__16752),
            .I(N__16738));
    LocalMux I__2245 (
            .O(N__16749),
            .I(N__16735));
    InMux I__2244 (
            .O(N__16748),
            .I(N__16728));
    InMux I__2243 (
            .O(N__16747),
            .I(N__16728));
    InMux I__2242 (
            .O(N__16746),
            .I(N__16728));
    InMux I__2241 (
            .O(N__16745),
            .I(N__16724));
    InMux I__2240 (
            .O(N__16744),
            .I(N__16721));
    Span4Mux_v I__2239 (
            .O(N__16741),
            .I(N__16716));
    LocalMux I__2238 (
            .O(N__16738),
            .I(N__16716));
    Span4Mux_v I__2237 (
            .O(N__16735),
            .I(N__16711));
    LocalMux I__2236 (
            .O(N__16728),
            .I(N__16711));
    InMux I__2235 (
            .O(N__16727),
            .I(N__16708));
    LocalMux I__2234 (
            .O(N__16724),
            .I(N__16703));
    LocalMux I__2233 (
            .O(N__16721),
            .I(N__16703));
    Span4Mux_v I__2232 (
            .O(N__16716),
            .I(N__16700));
    Span4Mux_h I__2231 (
            .O(N__16711),
            .I(N__16697));
    LocalMux I__2230 (
            .O(N__16708),
            .I(SYNTHESIZED_WIRE_4_4));
    Odrv4 I__2229 (
            .O(N__16703),
            .I(SYNTHESIZED_WIRE_4_4));
    Odrv4 I__2228 (
            .O(N__16700),
            .I(SYNTHESIZED_WIRE_4_4));
    Odrv4 I__2227 (
            .O(N__16697),
            .I(SYNTHESIZED_WIRE_4_4));
    InMux I__2226 (
            .O(N__16688),
            .I(N__16685));
    LocalMux I__2225 (
            .O(N__16685),
            .I(\b2v_inst.g1_0_0 ));
    InMux I__2224 (
            .O(N__16682),
            .I(N__16679));
    LocalMux I__2223 (
            .O(N__16679),
            .I(\b2v_inst.g1_0_0Z0Z_2 ));
    CascadeMux I__2222 (
            .O(N__16676),
            .I(N__16673));
    InMux I__2221 (
            .O(N__16673),
            .I(N__16670));
    LocalMux I__2220 (
            .O(N__16670),
            .I(\b2v_inst.g1_0_a4Z0Z_0 ));
    InMux I__2219 (
            .O(N__16667),
            .I(N__16664));
    LocalMux I__2218 (
            .O(N__16664),
            .I(N__16661));
    Sp12to4 I__2217 (
            .O(N__16661),
            .I(N__16658));
    Span12Mux_v I__2216 (
            .O(N__16658),
            .I(N__16655));
    Span12Mux_h I__2215 (
            .O(N__16655),
            .I(N__16652));
    Odrv12 I__2214 (
            .O(N__16652),
            .I(swit_c_9));
    InMux I__2213 (
            .O(N__16649),
            .I(N__16646));
    LocalMux I__2212 (
            .O(N__16646),
            .I(\b2v_inst.addr_ram_energia_m0_9 ));
    CascadeMux I__2211 (
            .O(N__16643),
            .I(\b2v_inst1.N_38_cascade_ ));
    InMux I__2210 (
            .O(N__16640),
            .I(N__16633));
    InMux I__2209 (
            .O(N__16639),
            .I(N__16633));
    InMux I__2208 (
            .O(N__16638),
            .I(N__16624));
    LocalMux I__2207 (
            .O(N__16633),
            .I(N__16621));
    InMux I__2206 (
            .O(N__16632),
            .I(N__16618));
    InMux I__2205 (
            .O(N__16631),
            .I(N__16615));
    InMux I__2204 (
            .O(N__16630),
            .I(N__16612));
    InMux I__2203 (
            .O(N__16629),
            .I(N__16609));
    InMux I__2202 (
            .O(N__16628),
            .I(N__16606));
    InMux I__2201 (
            .O(N__16627),
            .I(N__16603));
    LocalMux I__2200 (
            .O(N__16624),
            .I(N__16596));
    Span4Mux_v I__2199 (
            .O(N__16621),
            .I(N__16596));
    LocalMux I__2198 (
            .O(N__16618),
            .I(N__16596));
    LocalMux I__2197 (
            .O(N__16615),
            .I(\b2v_inst1.r_Bit_IndexZ0Z_2 ));
    LocalMux I__2196 (
            .O(N__16612),
            .I(\b2v_inst1.r_Bit_IndexZ0Z_2 ));
    LocalMux I__2195 (
            .O(N__16609),
            .I(\b2v_inst1.r_Bit_IndexZ0Z_2 ));
    LocalMux I__2194 (
            .O(N__16606),
            .I(\b2v_inst1.r_Bit_IndexZ0Z_2 ));
    LocalMux I__2193 (
            .O(N__16603),
            .I(\b2v_inst1.r_Bit_IndexZ0Z_2 ));
    Odrv4 I__2192 (
            .O(N__16596),
            .I(\b2v_inst1.r_Bit_IndexZ0Z_2 ));
    InMux I__2191 (
            .O(N__16583),
            .I(N__16580));
    LocalMux I__2190 (
            .O(N__16580),
            .I(\b2v_inst1.N_44 ));
    CascadeMux I__2189 (
            .O(N__16577),
            .I(\b2v_inst1.N_96_cascade_ ));
    InMux I__2188 (
            .O(N__16574),
            .I(N__16571));
    LocalMux I__2187 (
            .O(N__16571),
            .I(\b2v_inst.g0_0_i_a4Z0Z_0 ));
    InMux I__2186 (
            .O(N__16568),
            .I(N__16565));
    LocalMux I__2185 (
            .O(N__16565),
            .I(N__16562));
    Odrv4 I__2184 (
            .O(N__16562),
            .I(\b2v_inst.g0_0_iZ0Z_2 ));
    CascadeMux I__2183 (
            .O(N__16559),
            .I(N__16556));
    InMux I__2182 (
            .O(N__16556),
            .I(N__16553));
    LocalMux I__2181 (
            .O(N__16553),
            .I(N__16550));
    Span12Mux_h I__2180 (
            .O(N__16550),
            .I(N__16547));
    Odrv12 I__2179 (
            .O(N__16547),
            .I(\b2v_inst.g2Z0Z_1 ));
    CascadeMux I__2178 (
            .O(N__16544),
            .I(\b2v_inst1.N_58_i_cascade_ ));
    InMux I__2177 (
            .O(N__16541),
            .I(N__16537));
    InMux I__2176 (
            .O(N__16540),
            .I(N__16533));
    LocalMux I__2175 (
            .O(N__16537),
            .I(N__16530));
    InMux I__2174 (
            .O(N__16536),
            .I(N__16527));
    LocalMux I__2173 (
            .O(N__16533),
            .I(N__16524));
    Odrv12 I__2172 (
            .O(N__16530),
            .I(\b2v_inst1.un22_r_clk_count_ac0_3 ));
    LocalMux I__2171 (
            .O(N__16527),
            .I(\b2v_inst1.un22_r_clk_count_ac0_3 ));
    Odrv4 I__2170 (
            .O(N__16524),
            .I(\b2v_inst1.un22_r_clk_count_ac0_3 ));
    InMux I__2169 (
            .O(N__16517),
            .I(\b2v_inst.un3_dir_mem_cry_5 ));
    InMux I__2168 (
            .O(N__16514),
            .I(\b2v_inst.un3_dir_mem_cry_6 ));
    InMux I__2167 (
            .O(N__16511),
            .I(bfn_8_10_0_));
    InMux I__2166 (
            .O(N__16508),
            .I(\b2v_inst.un3_dir_mem_cry_8 ));
    InMux I__2165 (
            .O(N__16505),
            .I(\b2v_inst.un3_dir_mem_cry_9 ));
    InMux I__2164 (
            .O(N__16502),
            .I(N__16495));
    InMux I__2163 (
            .O(N__16501),
            .I(N__16491));
    InMux I__2162 (
            .O(N__16500),
            .I(N__16488));
    InMux I__2161 (
            .O(N__16499),
            .I(N__16485));
    InMux I__2160 (
            .O(N__16498),
            .I(N__16482));
    LocalMux I__2159 (
            .O(N__16495),
            .I(N__16479));
    InMux I__2158 (
            .O(N__16494),
            .I(N__16476));
    LocalMux I__2157 (
            .O(N__16491),
            .I(N__16470));
    LocalMux I__2156 (
            .O(N__16488),
            .I(N__16465));
    LocalMux I__2155 (
            .O(N__16485),
            .I(N__16465));
    LocalMux I__2154 (
            .O(N__16482),
            .I(N__16458));
    Span4Mux_h I__2153 (
            .O(N__16479),
            .I(N__16458));
    LocalMux I__2152 (
            .O(N__16476),
            .I(N__16458));
    InMux I__2151 (
            .O(N__16475),
            .I(N__16453));
    InMux I__2150 (
            .O(N__16474),
            .I(N__16453));
    InMux I__2149 (
            .O(N__16473),
            .I(N__16450));
    Span4Mux_v I__2148 (
            .O(N__16470),
            .I(N__16447));
    Span4Mux_v I__2147 (
            .O(N__16465),
            .I(N__16442));
    Span4Mux_v I__2146 (
            .O(N__16458),
            .I(N__16442));
    LocalMux I__2145 (
            .O(N__16453),
            .I(N__16439));
    LocalMux I__2144 (
            .O(N__16450),
            .I(SYNTHESIZED_WIRE_4_13));
    Odrv4 I__2143 (
            .O(N__16447),
            .I(SYNTHESIZED_WIRE_4_13));
    Odrv4 I__2142 (
            .O(N__16442),
            .I(SYNTHESIZED_WIRE_4_13));
    Odrv4 I__2141 (
            .O(N__16439),
            .I(SYNTHESIZED_WIRE_4_13));
    InMux I__2140 (
            .O(N__16430),
            .I(N__16426));
    InMux I__2139 (
            .O(N__16429),
            .I(N__16420));
    LocalMux I__2138 (
            .O(N__16426),
            .I(N__16417));
    InMux I__2137 (
            .O(N__16425),
            .I(N__16414));
    InMux I__2136 (
            .O(N__16424),
            .I(N__16411));
    InMux I__2135 (
            .O(N__16423),
            .I(N__16404));
    LocalMux I__2134 (
            .O(N__16420),
            .I(N__16399));
    Span4Mux_h I__2133 (
            .O(N__16417),
            .I(N__16399));
    LocalMux I__2132 (
            .O(N__16414),
            .I(N__16394));
    LocalMux I__2131 (
            .O(N__16411),
            .I(N__16394));
    InMux I__2130 (
            .O(N__16410),
            .I(N__16387));
    InMux I__2129 (
            .O(N__16409),
            .I(N__16387));
    InMux I__2128 (
            .O(N__16408),
            .I(N__16387));
    InMux I__2127 (
            .O(N__16407),
            .I(N__16384));
    LocalMux I__2126 (
            .O(N__16404),
            .I(N__16379));
    Span4Mux_v I__2125 (
            .O(N__16399),
            .I(N__16379));
    Span4Mux_h I__2124 (
            .O(N__16394),
            .I(N__16376));
    LocalMux I__2123 (
            .O(N__16387),
            .I(N__16373));
    LocalMux I__2122 (
            .O(N__16384),
            .I(SYNTHESIZED_WIRE_4_15));
    Odrv4 I__2121 (
            .O(N__16379),
            .I(SYNTHESIZED_WIRE_4_15));
    Odrv4 I__2120 (
            .O(N__16376),
            .I(SYNTHESIZED_WIRE_4_15));
    Odrv4 I__2119 (
            .O(N__16373),
            .I(SYNTHESIZED_WIRE_4_15));
    CascadeMux I__2118 (
            .O(N__16364),
            .I(N__16359));
    InMux I__2117 (
            .O(N__16363),
            .I(N__16355));
    InMux I__2116 (
            .O(N__16362),
            .I(N__16351));
    InMux I__2115 (
            .O(N__16359),
            .I(N__16347));
    InMux I__2114 (
            .O(N__16358),
            .I(N__16344));
    LocalMux I__2113 (
            .O(N__16355),
            .I(N__16341));
    InMux I__2112 (
            .O(N__16354),
            .I(N__16335));
    LocalMux I__2111 (
            .O(N__16351),
            .I(N__16332));
    InMux I__2110 (
            .O(N__16350),
            .I(N__16329));
    LocalMux I__2109 (
            .O(N__16347),
            .I(N__16326));
    LocalMux I__2108 (
            .O(N__16344),
            .I(N__16323));
    Span4Mux_h I__2107 (
            .O(N__16341),
            .I(N__16320));
    InMux I__2106 (
            .O(N__16340),
            .I(N__16313));
    InMux I__2105 (
            .O(N__16339),
            .I(N__16313));
    InMux I__2104 (
            .O(N__16338),
            .I(N__16313));
    LocalMux I__2103 (
            .O(N__16335),
            .I(N__16306));
    Span4Mux_v I__2102 (
            .O(N__16332),
            .I(N__16306));
    LocalMux I__2101 (
            .O(N__16329),
            .I(N__16306));
    Span4Mux_h I__2100 (
            .O(N__16326),
            .I(N__16301));
    Span4Mux_h I__2099 (
            .O(N__16323),
            .I(N__16301));
    Span4Mux_v I__2098 (
            .O(N__16320),
            .I(N__16296));
    LocalMux I__2097 (
            .O(N__16313),
            .I(N__16296));
    Odrv4 I__2096 (
            .O(N__16306),
            .I(SYNTHESIZED_WIRE_4_14));
    Odrv4 I__2095 (
            .O(N__16301),
            .I(SYNTHESIZED_WIRE_4_14));
    Odrv4 I__2094 (
            .O(N__16296),
            .I(SYNTHESIZED_WIRE_4_14));
    InMux I__2093 (
            .O(N__16289),
            .I(N__16286));
    LocalMux I__2092 (
            .O(N__16286),
            .I(\b2v_inst.state_RNO_25Z0Z_29 ));
    InMux I__2091 (
            .O(N__16283),
            .I(N__16280));
    LocalMux I__2090 (
            .O(N__16280),
            .I(N__16277));
    Odrv4 I__2089 (
            .O(N__16277),
            .I(\b2v_inst.g2_1_0 ));
    CascadeMux I__2088 (
            .O(N__16274),
            .I(\b2v_inst.m29_2_cascade_ ));
    InMux I__2087 (
            .O(N__16271),
            .I(N__16268));
    LocalMux I__2086 (
            .O(N__16268),
            .I(N__16263));
    InMux I__2085 (
            .O(N__16267),
            .I(N__16260));
    InMux I__2084 (
            .O(N__16266),
            .I(N__16257));
    Odrv12 I__2083 (
            .O(N__16263),
            .I(\b2v_inst.un4_pix_count_intlto10_1_d_0 ));
    LocalMux I__2082 (
            .O(N__16260),
            .I(\b2v_inst.un4_pix_count_intlto10_1_d_0 ));
    LocalMux I__2081 (
            .O(N__16257),
            .I(\b2v_inst.un4_pix_count_intlto10_1_d_0 ));
    CascadeMux I__2080 (
            .O(N__16250),
            .I(N__16247));
    InMux I__2079 (
            .O(N__16247),
            .I(N__16242));
    InMux I__2078 (
            .O(N__16246),
            .I(N__16239));
    InMux I__2077 (
            .O(N__16245),
            .I(N__16236));
    LocalMux I__2076 (
            .O(N__16242),
            .I(N__16233));
    LocalMux I__2075 (
            .O(N__16239),
            .I(N__16230));
    LocalMux I__2074 (
            .O(N__16236),
            .I(N__16225));
    Span4Mux_v I__2073 (
            .O(N__16233),
            .I(N__16225));
    Odrv12 I__2072 (
            .O(N__16230),
            .I(\b2v_inst.indice_RNIJFHBZ0Z_0 ));
    Odrv4 I__2071 (
            .O(N__16225),
            .I(\b2v_inst.indice_RNIJFHBZ0Z_0 ));
    InMux I__2070 (
            .O(N__16220),
            .I(N__16217));
    LocalMux I__2069 (
            .O(N__16217),
            .I(N__16212));
    InMux I__2068 (
            .O(N__16216),
            .I(N__16209));
    InMux I__2067 (
            .O(N__16215),
            .I(N__16206));
    Span4Mux_h I__2066 (
            .O(N__16212),
            .I(N__16203));
    LocalMux I__2065 (
            .O(N__16209),
            .I(N__16200));
    LocalMux I__2064 (
            .O(N__16206),
            .I(\b2v_inst.un1_indice_cry_5_c_RNI69OGZ0 ));
    Odrv4 I__2063 (
            .O(N__16203),
            .I(\b2v_inst.un1_indice_cry_5_c_RNI69OGZ0 ));
    Odrv4 I__2062 (
            .O(N__16200),
            .I(\b2v_inst.un1_indice_cry_5_c_RNI69OGZ0 ));
    CascadeMux I__2061 (
            .O(N__16193),
            .I(N__16190));
    InMux I__2060 (
            .O(N__16190),
            .I(N__16187));
    LocalMux I__2059 (
            .O(N__16187),
            .I(N__16184));
    Span4Mux_v I__2058 (
            .O(N__16184),
            .I(N__16181));
    Span4Mux_h I__2057 (
            .O(N__16181),
            .I(N__16178));
    Odrv4 I__2056 (
            .O(N__16178),
            .I(\b2v_inst.dir_mem_3_RNO_0Z0Z_6 ));
    InMux I__2055 (
            .O(N__16175),
            .I(\b2v_inst.un3_dir_mem_cry_1 ));
    InMux I__2054 (
            .O(N__16172),
            .I(\b2v_inst.un3_dir_mem_cry_2 ));
    InMux I__2053 (
            .O(N__16169),
            .I(\b2v_inst.un3_dir_mem_cry_3 ));
    InMux I__2052 (
            .O(N__16166),
            .I(\b2v_inst.un3_dir_mem_cry_4 ));
    InMux I__2051 (
            .O(N__16163),
            .I(\b2v_inst.un2_dir_mem_1_cry_8 ));
    CascadeMux I__2050 (
            .O(N__16160),
            .I(N__16156));
    InMux I__2049 (
            .O(N__16159),
            .I(N__16151));
    InMux I__2048 (
            .O(N__16156),
            .I(N__16151));
    LocalMux I__2047 (
            .O(N__16151),
            .I(N__16147));
    InMux I__2046 (
            .O(N__16150),
            .I(N__16144));
    Odrv4 I__2045 (
            .O(N__16147),
            .I(\b2v_inst.un1_indice_cry_10_THRU_CO ));
    LocalMux I__2044 (
            .O(N__16144),
            .I(\b2v_inst.un1_indice_cry_10_THRU_CO ));
    CascadeMux I__2043 (
            .O(N__16139),
            .I(N__16136));
    InMux I__2042 (
            .O(N__16136),
            .I(N__16133));
    LocalMux I__2041 (
            .O(N__16133),
            .I(N__16130));
    Span4Mux_h I__2040 (
            .O(N__16130),
            .I(N__16127));
    Span4Mux_h I__2039 (
            .O(N__16127),
            .I(N__16124));
    Odrv4 I__2038 (
            .O(N__16124),
            .I(\b2v_inst.dir_mem_3_RNO_0Z0Z_10 ));
    CascadeMux I__2037 (
            .O(N__16121),
            .I(N__16118));
    InMux I__2036 (
            .O(N__16118),
            .I(N__16115));
    LocalMux I__2035 (
            .O(N__16115),
            .I(N__16112));
    Span4Mux_v I__2034 (
            .O(N__16112),
            .I(N__16109));
    Odrv4 I__2033 (
            .O(N__16109),
            .I(\b2v_inst.dir_mem_3_RNO_0Z0Z_7 ));
    CascadeMux I__2032 (
            .O(N__16106),
            .I(N__16103));
    InMux I__2031 (
            .O(N__16103),
            .I(N__16100));
    LocalMux I__2030 (
            .O(N__16100),
            .I(N__16097));
    Span4Mux_v I__2029 (
            .O(N__16097),
            .I(N__16094));
    Odrv4 I__2028 (
            .O(N__16094),
            .I(\b2v_inst.dir_mem_3_RNO_0Z0Z_8 ));
    CascadeMux I__2027 (
            .O(N__16091),
            .I(N__16088));
    InMux I__2026 (
            .O(N__16088),
            .I(N__16085));
    LocalMux I__2025 (
            .O(N__16085),
            .I(N__16082));
    Span4Mux_h I__2024 (
            .O(N__16082),
            .I(N__16079));
    Odrv4 I__2023 (
            .O(N__16079),
            .I(\b2v_inst.dir_mem_3_RNO_0Z0Z_9 ));
    InMux I__2022 (
            .O(N__16076),
            .I(N__16073));
    LocalMux I__2021 (
            .O(N__16073),
            .I(N__16068));
    InMux I__2020 (
            .O(N__16072),
            .I(N__16065));
    InMux I__2019 (
            .O(N__16071),
            .I(N__16062));
    Span4Mux_h I__2018 (
            .O(N__16068),
            .I(N__16059));
    LocalMux I__2017 (
            .O(N__16065),
            .I(N__16056));
    LocalMux I__2016 (
            .O(N__16062),
            .I(\b2v_inst.un1_indice_cry_2_c_RNI00LGZ0 ));
    Odrv4 I__2015 (
            .O(N__16059),
            .I(\b2v_inst.un1_indice_cry_2_c_RNI00LGZ0 ));
    Odrv4 I__2014 (
            .O(N__16056),
            .I(\b2v_inst.un1_indice_cry_2_c_RNI00LGZ0 ));
    InMux I__2013 (
            .O(N__16049),
            .I(\b2v_inst.un2_dir_mem_1_cry_3 ));
    InMux I__2012 (
            .O(N__16046),
            .I(\b2v_inst.un2_dir_mem_1_cry_4 ));
    InMux I__2011 (
            .O(N__16043),
            .I(\b2v_inst.un2_dir_mem_1_cry_5 ));
    InMux I__2010 (
            .O(N__16040),
            .I(\b2v_inst.un2_dir_mem_1_cry_6 ));
    InMux I__2009 (
            .O(N__16037),
            .I(bfn_8_6_0_));
    CascadeMux I__2008 (
            .O(N__16034),
            .I(N__16031));
    InMux I__2007 (
            .O(N__16031),
            .I(N__16028));
    LocalMux I__2006 (
            .O(N__16028),
            .I(\b2v_inst.N_8 ));
    InMux I__2005 (
            .O(N__16025),
            .I(N__16022));
    LocalMux I__2004 (
            .O(N__16022),
            .I(\b2v_inst1.N_42 ));
    InMux I__2003 (
            .O(N__16019),
            .I(N__16016));
    LocalMux I__2002 (
            .O(N__16016),
            .I(N__16012));
    InMux I__2001 (
            .O(N__16015),
            .I(N__16009));
    Odrv4 I__2000 (
            .O(N__16012),
            .I(\b2v_inst1.r_SM_Main_d_4 ));
    LocalMux I__1999 (
            .O(N__16009),
            .I(\b2v_inst1.r_SM_Main_d_4 ));
    InMux I__1998 (
            .O(N__16004),
            .I(N__15999));
    InMux I__1997 (
            .O(N__16003),
            .I(N__15994));
    InMux I__1996 (
            .O(N__16002),
            .I(N__15994));
    LocalMux I__1995 (
            .O(N__15999),
            .I(N__15989));
    LocalMux I__1994 (
            .O(N__15994),
            .I(N__15989));
    Odrv4 I__1993 (
            .O(N__15989),
            .I(\b2v_inst1.N_47 ));
    CascadeMux I__1992 (
            .O(N__15986),
            .I(\b2v_inst1.r_SM_Main_d_4_cascade_ ));
    InMux I__1991 (
            .O(N__15983),
            .I(N__15980));
    LocalMux I__1990 (
            .O(N__15980),
            .I(\b2v_inst1.N_51 ));
    CascadeMux I__1989 (
            .O(N__15977),
            .I(N__15973));
    CascadeMux I__1988 (
            .O(N__15976),
            .I(N__15970));
    CascadeBuf I__1987 (
            .O(N__15973),
            .I(N__15967));
    CascadeBuf I__1986 (
            .O(N__15970),
            .I(N__15964));
    CascadeMux I__1985 (
            .O(N__15967),
            .I(N__15961));
    CascadeMux I__1984 (
            .O(N__15964),
            .I(N__15958));
    CascadeBuf I__1983 (
            .O(N__15961),
            .I(N__15955));
    CascadeBuf I__1982 (
            .O(N__15958),
            .I(N__15952));
    CascadeMux I__1981 (
            .O(N__15955),
            .I(N__15949));
    CascadeMux I__1980 (
            .O(N__15952),
            .I(N__15946));
    CascadeBuf I__1979 (
            .O(N__15949),
            .I(N__15943));
    CascadeBuf I__1978 (
            .O(N__15946),
            .I(N__15940));
    CascadeMux I__1977 (
            .O(N__15943),
            .I(N__15937));
    CascadeMux I__1976 (
            .O(N__15940),
            .I(N__15934));
    CascadeBuf I__1975 (
            .O(N__15937),
            .I(N__15931));
    CascadeBuf I__1974 (
            .O(N__15934),
            .I(N__15928));
    CascadeMux I__1973 (
            .O(N__15931),
            .I(N__15925));
    CascadeMux I__1972 (
            .O(N__15928),
            .I(N__15922));
    CascadeBuf I__1971 (
            .O(N__15925),
            .I(N__15919));
    CascadeBuf I__1970 (
            .O(N__15922),
            .I(N__15916));
    CascadeMux I__1969 (
            .O(N__15919),
            .I(N__15913));
    CascadeMux I__1968 (
            .O(N__15916),
            .I(N__15910));
    CascadeBuf I__1967 (
            .O(N__15913),
            .I(N__15907));
    CascadeBuf I__1966 (
            .O(N__15910),
            .I(N__15904));
    CascadeMux I__1965 (
            .O(N__15907),
            .I(N__15901));
    CascadeMux I__1964 (
            .O(N__15904),
            .I(N__15898));
    InMux I__1963 (
            .O(N__15901),
            .I(N__15895));
    InMux I__1962 (
            .O(N__15898),
            .I(N__15892));
    LocalMux I__1961 (
            .O(N__15895),
            .I(N__15887));
    LocalMux I__1960 (
            .O(N__15892),
            .I(N__15887));
    Span4Mux_v I__1959 (
            .O(N__15887),
            .I(N__15884));
    Span4Mux_h I__1958 (
            .O(N__15884),
            .I(N__15881));
    Odrv4 I__1957 (
            .O(N__15881),
            .I(SYNTHESIZED_WIRE_12_9));
    InMux I__1956 (
            .O(N__15878),
            .I(N__15872));
    InMux I__1955 (
            .O(N__15877),
            .I(N__15869));
    InMux I__1954 (
            .O(N__15876),
            .I(N__15866));
    InMux I__1953 (
            .O(N__15875),
            .I(N__15863));
    LocalMux I__1952 (
            .O(N__15872),
            .I(N__15860));
    LocalMux I__1951 (
            .O(N__15869),
            .I(N__15854));
    LocalMux I__1950 (
            .O(N__15866),
            .I(N__15854));
    LocalMux I__1949 (
            .O(N__15863),
            .I(N__15849));
    Span4Mux_v I__1948 (
            .O(N__15860),
            .I(N__15849));
    CascadeMux I__1947 (
            .O(N__15859),
            .I(N__15845));
    Span4Mux_h I__1946 (
            .O(N__15854),
            .I(N__15842));
    Sp12to4 I__1945 (
            .O(N__15849),
            .I(N__15839));
    InMux I__1944 (
            .O(N__15848),
            .I(N__15834));
    InMux I__1943 (
            .O(N__15845),
            .I(N__15834));
    Odrv4 I__1942 (
            .O(N__15842),
            .I(SYNTHESIZED_WIRE_4_6));
    Odrv12 I__1941 (
            .O(N__15839),
            .I(SYNTHESIZED_WIRE_4_6));
    LocalMux I__1940 (
            .O(N__15834),
            .I(SYNTHESIZED_WIRE_4_6));
    InMux I__1939 (
            .O(N__15827),
            .I(N__15821));
    InMux I__1938 (
            .O(N__15826),
            .I(N__15818));
    InMux I__1937 (
            .O(N__15825),
            .I(N__15813));
    InMux I__1936 (
            .O(N__15824),
            .I(N__15813));
    LocalMux I__1935 (
            .O(N__15821),
            .I(N__15808));
    LocalMux I__1934 (
            .O(N__15818),
            .I(N__15808));
    LocalMux I__1933 (
            .O(N__15813),
            .I(N__15802));
    Span4Mux_h I__1932 (
            .O(N__15808),
            .I(N__15802));
    CascadeMux I__1931 (
            .O(N__15807),
            .I(N__15798));
    Span4Mux_h I__1930 (
            .O(N__15802),
            .I(N__15795));
    InMux I__1929 (
            .O(N__15801),
            .I(N__15792));
    InMux I__1928 (
            .O(N__15798),
            .I(N__15789));
    Odrv4 I__1927 (
            .O(N__15795),
            .I(SYNTHESIZED_WIRE_4_5));
    LocalMux I__1926 (
            .O(N__15792),
            .I(SYNTHESIZED_WIRE_4_5));
    LocalMux I__1925 (
            .O(N__15789),
            .I(SYNTHESIZED_WIRE_4_5));
    CascadeMux I__1924 (
            .O(N__15782),
            .I(\b2v_inst.un4_pix_count_intlto6_d_1_0_cascade_ ));
    CascadeMux I__1923 (
            .O(N__15779),
            .I(N__15775));
    CascadeMux I__1922 (
            .O(N__15778),
            .I(N__15770));
    InMux I__1921 (
            .O(N__15775),
            .I(N__15767));
    CascadeMux I__1920 (
            .O(N__15774),
            .I(N__15764));
    InMux I__1919 (
            .O(N__15773),
            .I(N__15761));
    InMux I__1918 (
            .O(N__15770),
            .I(N__15758));
    LocalMux I__1917 (
            .O(N__15767),
            .I(N__15755));
    InMux I__1916 (
            .O(N__15764),
            .I(N__15752));
    LocalMux I__1915 (
            .O(N__15761),
            .I(N__15749));
    LocalMux I__1914 (
            .O(N__15758),
            .I(N__15744));
    Span4Mux_v I__1913 (
            .O(N__15755),
            .I(N__15744));
    LocalMux I__1912 (
            .O(N__15752),
            .I(N__15741));
    Odrv4 I__1911 (
            .O(N__15749),
            .I(SYNTHESIZED_WIRE_4_10_rep1));
    Odrv4 I__1910 (
            .O(N__15744),
            .I(SYNTHESIZED_WIRE_4_10_rep1));
    Odrv4 I__1909 (
            .O(N__15741),
            .I(SYNTHESIZED_WIRE_4_10_rep1));
    CascadeMux I__1908 (
            .O(N__15734),
            .I(N__15731));
    InMux I__1907 (
            .O(N__15731),
            .I(N__15726));
    InMux I__1906 (
            .O(N__15730),
            .I(N__15722));
    InMux I__1905 (
            .O(N__15729),
            .I(N__15719));
    LocalMux I__1904 (
            .O(N__15726),
            .I(N__15716));
    InMux I__1903 (
            .O(N__15725),
            .I(N__15713));
    LocalMux I__1902 (
            .O(N__15722),
            .I(N__15710));
    LocalMux I__1901 (
            .O(N__15719),
            .I(N__15707));
    Span4Mux_h I__1900 (
            .O(N__15716),
            .I(N__15704));
    LocalMux I__1899 (
            .O(N__15713),
            .I(N__15699));
    Span4Mux_h I__1898 (
            .O(N__15710),
            .I(N__15699));
    Span4Mux_h I__1897 (
            .O(N__15707),
            .I(N__15696));
    Span4Mux_h I__1896 (
            .O(N__15704),
            .I(N__15693));
    Span4Mux_h I__1895 (
            .O(N__15699),
            .I(N__15690));
    Odrv4 I__1894 (
            .O(N__15696),
            .I(b2v_inst4_pix_count_int_fast_11));
    Odrv4 I__1893 (
            .O(N__15693),
            .I(b2v_inst4_pix_count_int_fast_11));
    Odrv4 I__1892 (
            .O(N__15690),
            .I(b2v_inst4_pix_count_int_fast_11));
    InMux I__1891 (
            .O(N__15683),
            .I(N__15678));
    CascadeMux I__1890 (
            .O(N__15682),
            .I(N__15675));
    InMux I__1889 (
            .O(N__15681),
            .I(N__15671));
    LocalMux I__1888 (
            .O(N__15678),
            .I(N__15668));
    InMux I__1887 (
            .O(N__15675),
            .I(N__15665));
    InMux I__1886 (
            .O(N__15674),
            .I(N__15662));
    LocalMux I__1885 (
            .O(N__15671),
            .I(N__15659));
    Span4Mux_v I__1884 (
            .O(N__15668),
            .I(N__15654));
    LocalMux I__1883 (
            .O(N__15665),
            .I(N__15654));
    LocalMux I__1882 (
            .O(N__15662),
            .I(N__15649));
    Span4Mux_h I__1881 (
            .O(N__15659),
            .I(N__15649));
    Span4Mux_h I__1880 (
            .O(N__15654),
            .I(N__15646));
    Odrv4 I__1879 (
            .O(N__15649),
            .I(b2v_inst4_pix_count_int_fast_12));
    Odrv4 I__1878 (
            .O(N__15646),
            .I(b2v_inst4_pix_count_int_fast_12));
    InMux I__1877 (
            .O(N__15641),
            .I(N__15638));
    LocalMux I__1876 (
            .O(N__15638),
            .I(N__15635));
    Span4Mux_h I__1875 (
            .O(N__15635),
            .I(N__15631));
    CascadeMux I__1874 (
            .O(N__15634),
            .I(N__15628));
    Span4Mux_h I__1873 (
            .O(N__15631),
            .I(N__15625));
    InMux I__1872 (
            .O(N__15628),
            .I(N__15622));
    Odrv4 I__1871 (
            .O(N__15625),
            .I(b2v_inst_un4_pix_count_intlto12_0));
    LocalMux I__1870 (
            .O(N__15622),
            .I(b2v_inst_un4_pix_count_intlto12_0));
    InMux I__1869 (
            .O(N__15617),
            .I(N__15613));
    InMux I__1868 (
            .O(N__15616),
            .I(N__15610));
    LocalMux I__1867 (
            .O(N__15613),
            .I(N__15606));
    LocalMux I__1866 (
            .O(N__15610),
            .I(N__15603));
    InMux I__1865 (
            .O(N__15609),
            .I(N__15600));
    Span4Mux_v I__1864 (
            .O(N__15606),
            .I(N__15593));
    Span4Mux_h I__1863 (
            .O(N__15603),
            .I(N__15588));
    LocalMux I__1862 (
            .O(N__15600),
            .I(N__15588));
    InMux I__1861 (
            .O(N__15599),
            .I(N__15585));
    InMux I__1860 (
            .O(N__15598),
            .I(N__15582));
    InMux I__1859 (
            .O(N__15597),
            .I(N__15577));
    InMux I__1858 (
            .O(N__15596),
            .I(N__15577));
    Odrv4 I__1857 (
            .O(N__15593),
            .I(SYNTHESIZED_WIRE_4_10));
    Odrv4 I__1856 (
            .O(N__15588),
            .I(SYNTHESIZED_WIRE_4_10));
    LocalMux I__1855 (
            .O(N__15585),
            .I(SYNTHESIZED_WIRE_4_10));
    LocalMux I__1854 (
            .O(N__15582),
            .I(SYNTHESIZED_WIRE_4_10));
    LocalMux I__1853 (
            .O(N__15577),
            .I(SYNTHESIZED_WIRE_4_10));
    InMux I__1852 (
            .O(N__15566),
            .I(N__15561));
    CascadeMux I__1851 (
            .O(N__15565),
            .I(N__15558));
    InMux I__1850 (
            .O(N__15564),
            .I(N__15555));
    LocalMux I__1849 (
            .O(N__15561),
            .I(N__15552));
    InMux I__1848 (
            .O(N__15558),
            .I(N__15549));
    LocalMux I__1847 (
            .O(N__15555),
            .I(N__15543));
    Span4Mux_v I__1846 (
            .O(N__15552),
            .I(N__15538));
    LocalMux I__1845 (
            .O(N__15549),
            .I(N__15538));
    InMux I__1844 (
            .O(N__15548),
            .I(N__15533));
    InMux I__1843 (
            .O(N__15547),
            .I(N__15533));
    CascadeMux I__1842 (
            .O(N__15546),
            .I(N__15530));
    Span4Mux_v I__1841 (
            .O(N__15543),
            .I(N__15526));
    Span4Mux_h I__1840 (
            .O(N__15538),
            .I(N__15521));
    LocalMux I__1839 (
            .O(N__15533),
            .I(N__15521));
    InMux I__1838 (
            .O(N__15530),
            .I(N__15518));
    InMux I__1837 (
            .O(N__15529),
            .I(N__15515));
    Odrv4 I__1836 (
            .O(N__15526),
            .I(SYNTHESIZED_WIRE_4_9));
    Odrv4 I__1835 (
            .O(N__15521),
            .I(SYNTHESIZED_WIRE_4_9));
    LocalMux I__1834 (
            .O(N__15518),
            .I(SYNTHESIZED_WIRE_4_9));
    LocalMux I__1833 (
            .O(N__15515),
            .I(SYNTHESIZED_WIRE_4_9));
    CascadeMux I__1832 (
            .O(N__15506),
            .I(b2v_inst_un4_pix_count_intlto12_0_cascade_));
    InMux I__1831 (
            .O(N__15503),
            .I(N__15496));
    InMux I__1830 (
            .O(N__15502),
            .I(N__15492));
    InMux I__1829 (
            .O(N__15501),
            .I(N__15487));
    InMux I__1828 (
            .O(N__15500),
            .I(N__15487));
    InMux I__1827 (
            .O(N__15499),
            .I(N__15484));
    LocalMux I__1826 (
            .O(N__15496),
            .I(N__15481));
    InMux I__1825 (
            .O(N__15495),
            .I(N__15478));
    LocalMux I__1824 (
            .O(N__15492),
            .I(N__15474));
    LocalMux I__1823 (
            .O(N__15487),
            .I(N__15471));
    LocalMux I__1822 (
            .O(N__15484),
            .I(N__15468));
    Span4Mux_v I__1821 (
            .O(N__15481),
            .I(N__15463));
    LocalMux I__1820 (
            .O(N__15478),
            .I(N__15463));
    InMux I__1819 (
            .O(N__15477),
            .I(N__15460));
    Span4Mux_v I__1818 (
            .O(N__15474),
            .I(N__15455));
    Span4Mux_v I__1817 (
            .O(N__15471),
            .I(N__15455));
    Span4Mux_h I__1816 (
            .O(N__15468),
            .I(N__15450));
    Span4Mux_h I__1815 (
            .O(N__15463),
            .I(N__15450));
    LocalMux I__1814 (
            .O(N__15460),
            .I(SYNTHESIZED_WIRE_4_8));
    Odrv4 I__1813 (
            .O(N__15455),
            .I(SYNTHESIZED_WIRE_4_8));
    Odrv4 I__1812 (
            .O(N__15450),
            .I(SYNTHESIZED_WIRE_4_8));
    InMux I__1811 (
            .O(N__15443),
            .I(N__15440));
    LocalMux I__1810 (
            .O(N__15440),
            .I(N__15437));
    Odrv12 I__1809 (
            .O(N__15437),
            .I(N_457_i));
    InMux I__1808 (
            .O(N__15434),
            .I(N__15431));
    LocalMux I__1807 (
            .O(N__15431),
            .I(\b2v_inst1.N_48 ));
    CascadeMux I__1806 (
            .O(N__15428),
            .I(\b2v_inst1.N_44_cascade_ ));
    InMux I__1805 (
            .O(N__15425),
            .I(N__15422));
    LocalMux I__1804 (
            .O(N__15422),
            .I(\b2v_inst.un4_pix_count_intlto10_1_0Z0Z_0 ));
    CascadeMux I__1803 (
            .O(N__15419),
            .I(\b2v_inst.un4_pix_count_intlt8_cascade_ ));
    InMux I__1802 (
            .O(N__15416),
            .I(N__15413));
    LocalMux I__1801 (
            .O(N__15413),
            .I(\b2v_inst.un4_pix_count_intlto15_1_aZ0Z0 ));
    InMux I__1800 (
            .O(N__15410),
            .I(N__15406));
    InMux I__1799 (
            .O(N__15409),
            .I(N__15403));
    LocalMux I__1798 (
            .O(N__15406),
            .I(\b2v_inst.un4_pix_count_intlt16 ));
    LocalMux I__1797 (
            .O(N__15403),
            .I(\b2v_inst.un4_pix_count_intlt16 ));
    CascadeMux I__1796 (
            .O(N__15398),
            .I(N__15393));
    InMux I__1795 (
            .O(N__15397),
            .I(N__15387));
    InMux I__1794 (
            .O(N__15396),
            .I(N__15387));
    InMux I__1793 (
            .O(N__15393),
            .I(N__15384));
    InMux I__1792 (
            .O(N__15392),
            .I(N__15381));
    LocalMux I__1791 (
            .O(N__15387),
            .I(N__15378));
    LocalMux I__1790 (
            .O(N__15384),
            .I(N__15371));
    LocalMux I__1789 (
            .O(N__15381),
            .I(N__15371));
    Span4Mux_h I__1788 (
            .O(N__15378),
            .I(N__15368));
    InMux I__1787 (
            .O(N__15377),
            .I(N__15363));
    InMux I__1786 (
            .O(N__15376),
            .I(N__15363));
    Odrv4 I__1785 (
            .O(N__15371),
            .I(SYNTHESIZED_WIRE_4_12));
    Odrv4 I__1784 (
            .O(N__15368),
            .I(SYNTHESIZED_WIRE_4_12));
    LocalMux I__1783 (
            .O(N__15363),
            .I(SYNTHESIZED_WIRE_4_12));
    CascadeMux I__1782 (
            .O(N__15356),
            .I(N__15353));
    InMux I__1781 (
            .O(N__15353),
            .I(N__15349));
    InMux I__1780 (
            .O(N__15352),
            .I(N__15346));
    LocalMux I__1779 (
            .O(N__15349),
            .I(N__15337));
    LocalMux I__1778 (
            .O(N__15346),
            .I(N__15337));
    InMux I__1777 (
            .O(N__15345),
            .I(N__15332));
    InMux I__1776 (
            .O(N__15344),
            .I(N__15332));
    InMux I__1775 (
            .O(N__15343),
            .I(N__15327));
    InMux I__1774 (
            .O(N__15342),
            .I(N__15327));
    Odrv4 I__1773 (
            .O(N__15337),
            .I(SYNTHESIZED_WIRE_4_11));
    LocalMux I__1772 (
            .O(N__15332),
            .I(SYNTHESIZED_WIRE_4_11));
    LocalMux I__1771 (
            .O(N__15327),
            .I(SYNTHESIZED_WIRE_4_11));
    InMux I__1770 (
            .O(N__15320),
            .I(N__15316));
    InMux I__1769 (
            .O(N__15319),
            .I(N__15313));
    LocalMux I__1768 (
            .O(N__15316),
            .I(N__15310));
    LocalMux I__1767 (
            .O(N__15313),
            .I(N__15307));
    Span4Mux_h I__1766 (
            .O(N__15310),
            .I(N__15302));
    Span4Mux_v I__1765 (
            .O(N__15307),
            .I(N__15299));
    InMux I__1764 (
            .O(N__15306),
            .I(N__15294));
    InMux I__1763 (
            .O(N__15305),
            .I(N__15294));
    Odrv4 I__1762 (
            .O(N__15302),
            .I(SYNTHESIZED_WIRE_4_9_rep1));
    Odrv4 I__1761 (
            .O(N__15299),
            .I(SYNTHESIZED_WIRE_4_9_rep1));
    LocalMux I__1760 (
            .O(N__15294),
            .I(SYNTHESIZED_WIRE_4_9_rep1));
    CascadeMux I__1759 (
            .O(N__15287),
            .I(\b2v_inst1.r_RX_Bytece_0_4_cascade_ ));
    CascadeMux I__1758 (
            .O(N__15284),
            .I(\b2v_inst.un4_pix_count_intlto10_1_d_0_xZ0Z1_cascade_ ));
    InMux I__1757 (
            .O(N__15281),
            .I(N__15277));
    InMux I__1756 (
            .O(N__15280),
            .I(N__15274));
    LocalMux I__1755 (
            .O(N__15277),
            .I(N__15266));
    LocalMux I__1754 (
            .O(N__15274),
            .I(N__15266));
    InMux I__1753 (
            .O(N__15273),
            .I(N__15263));
    InMux I__1752 (
            .O(N__15272),
            .I(N__15257));
    InMux I__1751 (
            .O(N__15271),
            .I(N__15257));
    Span4Mux_h I__1750 (
            .O(N__15266),
            .I(N__15254));
    LocalMux I__1749 (
            .O(N__15263),
            .I(N__15251));
    InMux I__1748 (
            .O(N__15262),
            .I(N__15248));
    LocalMux I__1747 (
            .O(N__15257),
            .I(SYNTHESIZED_WIRE_4_0));
    Odrv4 I__1746 (
            .O(N__15254),
            .I(SYNTHESIZED_WIRE_4_0));
    Odrv4 I__1745 (
            .O(N__15251),
            .I(SYNTHESIZED_WIRE_4_0));
    LocalMux I__1744 (
            .O(N__15248),
            .I(SYNTHESIZED_WIRE_4_0));
    CascadeMux I__1743 (
            .O(N__15239),
            .I(N__15233));
    InMux I__1742 (
            .O(N__15238),
            .I(N__15230));
    InMux I__1741 (
            .O(N__15237),
            .I(N__15227));
    InMux I__1740 (
            .O(N__15236),
            .I(N__15220));
    InMux I__1739 (
            .O(N__15233),
            .I(N__15220));
    LocalMux I__1738 (
            .O(N__15230),
            .I(N__15215));
    LocalMux I__1737 (
            .O(N__15227),
            .I(N__15215));
    InMux I__1736 (
            .O(N__15226),
            .I(N__15212));
    InMux I__1735 (
            .O(N__15225),
            .I(N__15209));
    LocalMux I__1734 (
            .O(N__15220),
            .I(SYNTHESIZED_WIRE_4_3));
    Odrv12 I__1733 (
            .O(N__15215),
            .I(SYNTHESIZED_WIRE_4_3));
    LocalMux I__1732 (
            .O(N__15212),
            .I(SYNTHESIZED_WIRE_4_3));
    LocalMux I__1731 (
            .O(N__15209),
            .I(SYNTHESIZED_WIRE_4_3));
    CascadeMux I__1730 (
            .O(N__15200),
            .I(N__15194));
    CascadeMux I__1729 (
            .O(N__15199),
            .I(N__15190));
    CascadeMux I__1728 (
            .O(N__15198),
            .I(N__15187));
    InMux I__1727 (
            .O(N__15197),
            .I(N__15184));
    InMux I__1726 (
            .O(N__15194),
            .I(N__15181));
    InMux I__1725 (
            .O(N__15193),
            .I(N__15178));
    InMux I__1724 (
            .O(N__15190),
            .I(N__15175));
    InMux I__1723 (
            .O(N__15187),
            .I(N__15172));
    LocalMux I__1722 (
            .O(N__15184),
            .I(N__15166));
    LocalMux I__1721 (
            .O(N__15181),
            .I(N__15166));
    LocalMux I__1720 (
            .O(N__15178),
            .I(N__15163));
    LocalMux I__1719 (
            .O(N__15175),
            .I(N__15158));
    LocalMux I__1718 (
            .O(N__15172),
            .I(N__15158));
    InMux I__1717 (
            .O(N__15171),
            .I(N__15155));
    Span4Mux_h I__1716 (
            .O(N__15166),
            .I(N__15152));
    Span4Mux_v I__1715 (
            .O(N__15163),
            .I(N__15147));
    Span4Mux_h I__1714 (
            .O(N__15158),
            .I(N__15147));
    LocalMux I__1713 (
            .O(N__15155),
            .I(SYNTHESIZED_WIRE_4_1));
    Odrv4 I__1712 (
            .O(N__15152),
            .I(SYNTHESIZED_WIRE_4_1));
    Odrv4 I__1711 (
            .O(N__15147),
            .I(SYNTHESIZED_WIRE_4_1));
    InMux I__1710 (
            .O(N__15140),
            .I(N__15136));
    InMux I__1709 (
            .O(N__15139),
            .I(N__15133));
    LocalMux I__1708 (
            .O(N__15136),
            .I(N__15127));
    LocalMux I__1707 (
            .O(N__15133),
            .I(N__15127));
    InMux I__1706 (
            .O(N__15132),
            .I(N__15124));
    Span4Mux_h I__1705 (
            .O(N__15127),
            .I(N__15118));
    LocalMux I__1704 (
            .O(N__15124),
            .I(N__15115));
    InMux I__1703 (
            .O(N__15123),
            .I(N__15108));
    InMux I__1702 (
            .O(N__15122),
            .I(N__15108));
    InMux I__1701 (
            .O(N__15121),
            .I(N__15108));
    Odrv4 I__1700 (
            .O(N__15118),
            .I(SYNTHESIZED_WIRE_4_2));
    Odrv4 I__1699 (
            .O(N__15115),
            .I(SYNTHESIZED_WIRE_4_2));
    LocalMux I__1698 (
            .O(N__15108),
            .I(SYNTHESIZED_WIRE_4_2));
    CascadeMux I__1697 (
            .O(N__15101),
            .I(\b2v_inst.dir_mem_316lt6_0_cascade_ ));
    InMux I__1696 (
            .O(N__15098),
            .I(N__15095));
    LocalMux I__1695 (
            .O(N__15095),
            .I(\b2v_inst.dir_mem_316lt7 ));
    InMux I__1694 (
            .O(N__15092),
            .I(N__15089));
    LocalMux I__1693 (
            .O(N__15089),
            .I(N__15084));
    InMux I__1692 (
            .O(N__15088),
            .I(N__15081));
    InMux I__1691 (
            .O(N__15087),
            .I(N__15078));
    Span4Mux_v I__1690 (
            .O(N__15084),
            .I(N__15073));
    LocalMux I__1689 (
            .O(N__15081),
            .I(N__15073));
    LocalMux I__1688 (
            .O(N__15078),
            .I(\b2v_inst.un1_indice_cry_1_c_RNIUSJGZ0 ));
    Odrv4 I__1687 (
            .O(N__15073),
            .I(\b2v_inst.un1_indice_cry_1_c_RNIUSJGZ0 ));
    InMux I__1686 (
            .O(N__15068),
            .I(N__15065));
    LocalMux I__1685 (
            .O(N__15065),
            .I(SYNTHESIZED_WIRE_4_fast_10));
    InMux I__1684 (
            .O(N__15062),
            .I(N__15059));
    LocalMux I__1683 (
            .O(N__15059),
            .I(N__15056));
    Odrv4 I__1682 (
            .O(N__15056),
            .I(SYNTHESIZED_WIRE_4_fast_9));
    CascadeMux I__1681 (
            .O(N__15053),
            .I(\b2v_inst.N_9_cascade_ ));
    InMux I__1680 (
            .O(N__15050),
            .I(N__15047));
    LocalMux I__1679 (
            .O(N__15047),
            .I(N__15044));
    Span4Mux_h I__1678 (
            .O(N__15044),
            .I(N__15038));
    InMux I__1677 (
            .O(N__15043),
            .I(N__15035));
    InMux I__1676 (
            .O(N__15042),
            .I(N__15030));
    InMux I__1675 (
            .O(N__15041),
            .I(N__15030));
    Odrv4 I__1674 (
            .O(N__15038),
            .I(b2v_inst4_pix_count_int_fast_5));
    LocalMux I__1673 (
            .O(N__15035),
            .I(b2v_inst4_pix_count_int_fast_5));
    LocalMux I__1672 (
            .O(N__15030),
            .I(b2v_inst4_pix_count_int_fast_5));
    InMux I__1671 (
            .O(N__15023),
            .I(N__15020));
    LocalMux I__1670 (
            .O(N__15020),
            .I(N__15014));
    InMux I__1669 (
            .O(N__15019),
            .I(N__15007));
    InMux I__1668 (
            .O(N__15018),
            .I(N__15007));
    InMux I__1667 (
            .O(N__15017),
            .I(N__15007));
    Odrv12 I__1666 (
            .O(N__15014),
            .I(b2v_inst4_pix_count_int_fast_6));
    LocalMux I__1665 (
            .O(N__15007),
            .I(b2v_inst4_pix_count_int_fast_6));
    InMux I__1664 (
            .O(N__15002),
            .I(N__14999));
    LocalMux I__1663 (
            .O(N__14999),
            .I(N__14996));
    Odrv12 I__1662 (
            .O(N__14996),
            .I(\b2v_inst.un4_pix_count_intlto6_1_xZ0Z1 ));
    InMux I__1661 (
            .O(N__14993),
            .I(N__14990));
    LocalMux I__1660 (
            .O(N__14990),
            .I(N__14987));
    Span4Mux_h I__1659 (
            .O(N__14987),
            .I(N__14984));
    Odrv4 I__1658 (
            .O(N__14984),
            .I(\b2v_inst.un4_pix_count_intlto6_1_xZ0Z0 ));
    InMux I__1657 (
            .O(N__14981),
            .I(N__14978));
    LocalMux I__1656 (
            .O(N__14978),
            .I(N__14975));
    Span4Mux_h I__1655 (
            .O(N__14975),
            .I(N__14972));
    Span4Mux_h I__1654 (
            .O(N__14972),
            .I(N__14969));
    Odrv4 I__1653 (
            .O(N__14969),
            .I(\b2v_inst.un4_pix_count_intlto6_dZ0Z_1 ));
    InMux I__1652 (
            .O(N__14966),
            .I(\b2v_inst.un8_dir_mem_1_cry_4 ));
    InMux I__1651 (
            .O(N__14963),
            .I(\b2v_inst.un8_dir_mem_1_cry_5 ));
    InMux I__1650 (
            .O(N__14960),
            .I(\b2v_inst.un8_dir_mem_1_cry_6 ));
    InMux I__1649 (
            .O(N__14957),
            .I(bfn_7_7_0_));
    InMux I__1648 (
            .O(N__14954),
            .I(\b2v_inst.un8_dir_mem_1_cry_8 ));
    InMux I__1647 (
            .O(N__14951),
            .I(\b2v_inst.un8_dir_mem_1_cry_9 ));
    InMux I__1646 (
            .O(N__14948),
            .I(\b2v_inst.un8_dir_mem_1_cry_10 ));
    InMux I__1645 (
            .O(N__14945),
            .I(N__14942));
    LocalMux I__1644 (
            .O(N__14942),
            .I(\b2v_inst1.N_40 ));
    InMux I__1643 (
            .O(N__14939),
            .I(\b2v_inst.un8_dir_mem_1_cry_0 ));
    InMux I__1642 (
            .O(N__14936),
            .I(\b2v_inst.un8_dir_mem_1_cry_1 ));
    InMux I__1641 (
            .O(N__14933),
            .I(\b2v_inst.un8_dir_mem_1_cry_2 ));
    InMux I__1640 (
            .O(N__14930),
            .I(\b2v_inst.un8_dir_mem_1_cry_3 ));
    IoInMux I__1639 (
            .O(N__14927),
            .I(N__14924));
    LocalMux I__1638 (
            .O(N__14924),
            .I(N__14921));
    Span4Mux_s1_h I__1637 (
            .O(N__14921),
            .I(N__14918));
    Span4Mux_h I__1636 (
            .O(N__14918),
            .I(N__14915));
    Span4Mux_h I__1635 (
            .O(N__14915),
            .I(N__14912));
    Odrv4 I__1634 (
            .O(N__14912),
            .I(\b2v_inst.N_305_1 ));
    CEMux I__1633 (
            .O(N__14909),
            .I(N__14906));
    LocalMux I__1632 (
            .O(N__14906),
            .I(N__14903));
    Span4Mux_v I__1631 (
            .O(N__14903),
            .I(N__14900));
    Odrv4 I__1630 (
            .O(N__14900),
            .I(\b2v_inst.un1_state_36_0 ));
    InMux I__1629 (
            .O(N__14897),
            .I(N__14892));
    InMux I__1628 (
            .O(N__14896),
            .I(N__14889));
    InMux I__1627 (
            .O(N__14895),
            .I(N__14886));
    LocalMux I__1626 (
            .O(N__14892),
            .I(N__14881));
    LocalMux I__1625 (
            .O(N__14889),
            .I(N__14881));
    LocalMux I__1624 (
            .O(N__14886),
            .I(\b2v_inst4.stateZ0Z_0 ));
    Odrv12 I__1623 (
            .O(N__14881),
            .I(\b2v_inst4.stateZ0Z_0 ));
    InMux I__1622 (
            .O(N__14876),
            .I(N__14872));
    InMux I__1621 (
            .O(N__14875),
            .I(N__14869));
    LocalMux I__1620 (
            .O(N__14872),
            .I(N__14866));
    LocalMux I__1619 (
            .O(N__14869),
            .I(N__14861));
    Span4Mux_h I__1618 (
            .O(N__14866),
            .I(N__14858));
    InMux I__1617 (
            .O(N__14865),
            .I(N__14853));
    InMux I__1616 (
            .O(N__14864),
            .I(N__14853));
    Odrv12 I__1615 (
            .O(N__14861),
            .I(SYNTHESIZED_WIRE_9));
    Odrv4 I__1614 (
            .O(N__14858),
            .I(SYNTHESIZED_WIRE_9));
    LocalMux I__1613 (
            .O(N__14853),
            .I(SYNTHESIZED_WIRE_9));
    CascadeMux I__1612 (
            .O(N__14846),
            .I(N__14843));
    InMux I__1611 (
            .O(N__14843),
            .I(N__14840));
    LocalMux I__1610 (
            .O(N__14840),
            .I(N__14837));
    Odrv4 I__1609 (
            .O(N__14837),
            .I(\b2v_inst.un1_state_36_0_a2_0_1_mbZ0Z_1 ));
    InMux I__1608 (
            .O(N__14834),
            .I(N__14825));
    InMux I__1607 (
            .O(N__14833),
            .I(N__14825));
    InMux I__1606 (
            .O(N__14832),
            .I(N__14825));
    LocalMux I__1605 (
            .O(N__14825),
            .I(N__14822));
    Span4Mux_h I__1604 (
            .O(N__14822),
            .I(N__14819));
    Odrv4 I__1603 (
            .O(N__14819),
            .I(\b2v_inst4.un1_pix_count_int_cry_9_c_RNIB86JZ0 ));
    InMux I__1602 (
            .O(N__14816),
            .I(N__14813));
    LocalMux I__1601 (
            .O(N__14813),
            .I(N__14808));
    InMux I__1600 (
            .O(N__14812),
            .I(N__14803));
    InMux I__1599 (
            .O(N__14811),
            .I(N__14803));
    Span4Mux_h I__1598 (
            .O(N__14808),
            .I(N__14800));
    LocalMux I__1597 (
            .O(N__14803),
            .I(N__14797));
    Odrv4 I__1596 (
            .O(N__14800),
            .I(\b2v_inst4.un1_pix_count_int_cry_8_c_RNI25BIZ0 ));
    Odrv4 I__1595 (
            .O(N__14797),
            .I(\b2v_inst4.un1_pix_count_int_cry_8_c_RNI25BIZ0 ));
    CascadeMux I__1594 (
            .O(N__14792),
            .I(N__14780));
    InMux I__1593 (
            .O(N__14791),
            .I(N__14774));
    InMux I__1592 (
            .O(N__14790),
            .I(N__14771));
    InMux I__1591 (
            .O(N__14789),
            .I(N__14768));
    InMux I__1590 (
            .O(N__14788),
            .I(N__14765));
    InMux I__1589 (
            .O(N__14787),
            .I(N__14762));
    InMux I__1588 (
            .O(N__14786),
            .I(N__14755));
    InMux I__1587 (
            .O(N__14785),
            .I(N__14755));
    InMux I__1586 (
            .O(N__14784),
            .I(N__14755));
    InMux I__1585 (
            .O(N__14783),
            .I(N__14740));
    InMux I__1584 (
            .O(N__14780),
            .I(N__14740));
    InMux I__1583 (
            .O(N__14779),
            .I(N__14740));
    InMux I__1582 (
            .O(N__14778),
            .I(N__14740));
    InMux I__1581 (
            .O(N__14777),
            .I(N__14740));
    LocalMux I__1580 (
            .O(N__14774),
            .I(N__14737));
    LocalMux I__1579 (
            .O(N__14771),
            .I(N__14734));
    LocalMux I__1578 (
            .O(N__14768),
            .I(N__14731));
    LocalMux I__1577 (
            .O(N__14765),
            .I(N__14726));
    LocalMux I__1576 (
            .O(N__14762),
            .I(N__14726));
    LocalMux I__1575 (
            .O(N__14755),
            .I(N__14723));
    InMux I__1574 (
            .O(N__14754),
            .I(N__14714));
    InMux I__1573 (
            .O(N__14753),
            .I(N__14714));
    InMux I__1572 (
            .O(N__14752),
            .I(N__14714));
    InMux I__1571 (
            .O(N__14751),
            .I(N__14714));
    LocalMux I__1570 (
            .O(N__14740),
            .I(N__14711));
    Span4Mux_h I__1569 (
            .O(N__14737),
            .I(N__14708));
    Span4Mux_h I__1568 (
            .O(N__14734),
            .I(N__14705));
    Span4Mux_h I__1567 (
            .O(N__14731),
            .I(N__14698));
    Span4Mux_h I__1566 (
            .O(N__14726),
            .I(N__14698));
    Span4Mux_h I__1565 (
            .O(N__14723),
            .I(N__14698));
    LocalMux I__1564 (
            .O(N__14714),
            .I(\b2v_inst4.un1_pix_count_int_0_sqmuxa_0 ));
    Odrv4 I__1563 (
            .O(N__14711),
            .I(\b2v_inst4.un1_pix_count_int_0_sqmuxa_0 ));
    Odrv4 I__1562 (
            .O(N__14708),
            .I(\b2v_inst4.un1_pix_count_int_0_sqmuxa_0 ));
    Odrv4 I__1561 (
            .O(N__14705),
            .I(\b2v_inst4.un1_pix_count_int_0_sqmuxa_0 ));
    Odrv4 I__1560 (
            .O(N__14698),
            .I(\b2v_inst4.un1_pix_count_int_0_sqmuxa_0 ));
    InMux I__1559 (
            .O(N__14687),
            .I(N__14684));
    LocalMux I__1558 (
            .O(N__14684),
            .I(N__14680));
    InMux I__1557 (
            .O(N__14683),
            .I(N__14677));
    Span4Mux_h I__1556 (
            .O(N__14680),
            .I(N__14674));
    LocalMux I__1555 (
            .O(N__14677),
            .I(N__14671));
    Odrv4 I__1554 (
            .O(N__14674),
            .I(\b2v_inst4.un1_pix_count_int_cry_10_c_RNIKMUJZ0 ));
    Odrv4 I__1553 (
            .O(N__14671),
            .I(\b2v_inst4.un1_pix_count_int_cry_10_c_RNIKMUJZ0 ));
    InMux I__1552 (
            .O(N__14666),
            .I(N__14663));
    LocalMux I__1551 (
            .O(N__14663),
            .I(N__14660));
    Odrv4 I__1550 (
            .O(N__14660),
            .I(\b2v_inst.ignorar_ancho_1_RNOZ0Z_0 ));
    CascadeMux I__1549 (
            .O(N__14657),
            .I(\b2v_inst.N_482_cascade_ ));
    CEMux I__1548 (
            .O(N__14654),
            .I(N__14651));
    LocalMux I__1547 (
            .O(N__14651),
            .I(N__14648));
    Odrv4 I__1546 (
            .O(N__14648),
            .I(\b2v_inst.un1_state_34_0 ));
    InMux I__1545 (
            .O(N__14645),
            .I(N__14642));
    LocalMux I__1544 (
            .O(N__14642),
            .I(N__14637));
    InMux I__1543 (
            .O(N__14641),
            .I(N__14632));
    InMux I__1542 (
            .O(N__14640),
            .I(N__14632));
    Span4Mux_v I__1541 (
            .O(N__14637),
            .I(N__14629));
    LocalMux I__1540 (
            .O(N__14632),
            .I(N__14626));
    Odrv4 I__1539 (
            .O(N__14629),
            .I(\b2v_inst.un1_cuenta_pixel_cry_8_c_RNIMU4IZ0 ));
    Odrv4 I__1538 (
            .O(N__14626),
            .I(\b2v_inst.un1_cuenta_pixel_cry_8_c_RNIMU4IZ0 ));
    InMux I__1537 (
            .O(N__14621),
            .I(N__14618));
    LocalMux I__1536 (
            .O(N__14618),
            .I(N__14613));
    InMux I__1535 (
            .O(N__14617),
            .I(N__14610));
    InMux I__1534 (
            .O(N__14616),
            .I(N__14607));
    Span4Mux_h I__1533 (
            .O(N__14613),
            .I(N__14604));
    LocalMux I__1532 (
            .O(N__14610),
            .I(N__14601));
    LocalMux I__1531 (
            .O(N__14607),
            .I(\b2v_inst.cuenta_pixel_RNIVBL9Z0Z_10 ));
    Odrv4 I__1530 (
            .O(N__14604),
            .I(\b2v_inst.cuenta_pixel_RNIVBL9Z0Z_10 ));
    Odrv4 I__1529 (
            .O(N__14601),
            .I(\b2v_inst.cuenta_pixel_RNIVBL9Z0Z_10 ));
    CascadeMux I__1528 (
            .O(N__14594),
            .I(N__14591));
    InMux I__1527 (
            .O(N__14591),
            .I(N__14587));
    CascadeMux I__1526 (
            .O(N__14590),
            .I(N__14584));
    LocalMux I__1525 (
            .O(N__14587),
            .I(N__14580));
    InMux I__1524 (
            .O(N__14584),
            .I(N__14577));
    InMux I__1523 (
            .O(N__14583),
            .I(N__14574));
    Span4Mux_h I__1522 (
            .O(N__14580),
            .I(N__14571));
    LocalMux I__1521 (
            .O(N__14577),
            .I(N__14568));
    LocalMux I__1520 (
            .O(N__14574),
            .I(\b2v_inst.un1_cuenta_pixel_cry_7_c_RNIKR3IZ0 ));
    Odrv4 I__1519 (
            .O(N__14571),
            .I(\b2v_inst.un1_cuenta_pixel_cry_7_c_RNIKR3IZ0 ));
    Odrv4 I__1518 (
            .O(N__14568),
            .I(\b2v_inst.un1_cuenta_pixel_cry_7_c_RNIKR3IZ0 ));
    InMux I__1517 (
            .O(N__14561),
            .I(N__14558));
    LocalMux I__1516 (
            .O(N__14558),
            .I(N__14554));
    InMux I__1515 (
            .O(N__14557),
            .I(N__14551));
    Span4Mux_h I__1514 (
            .O(N__14554),
            .I(N__14548));
    LocalMux I__1513 (
            .O(N__14551),
            .I(\b2v_inst.cuenta_pixel_5_i_a2_1_1_0_5 ));
    Odrv4 I__1512 (
            .O(N__14548),
            .I(\b2v_inst.cuenta_pixel_5_i_a2_1_1_0_5 ));
    InMux I__1511 (
            .O(N__14543),
            .I(N__14540));
    LocalMux I__1510 (
            .O(N__14540),
            .I(N__14536));
    InMux I__1509 (
            .O(N__14539),
            .I(N__14533));
    Odrv4 I__1508 (
            .O(N__14536),
            .I(\b2v_inst.N_325 ));
    LocalMux I__1507 (
            .O(N__14533),
            .I(\b2v_inst.N_325 ));
    InMux I__1506 (
            .O(N__14528),
            .I(N__14525));
    LocalMux I__1505 (
            .O(N__14525),
            .I(N__14522));
    Odrv4 I__1504 (
            .O(N__14522),
            .I(\b2v_inst.un1_state_36_0_rn_1 ));
    InMux I__1503 (
            .O(N__14519),
            .I(N__14516));
    LocalMux I__1502 (
            .O(N__14516),
            .I(N__14513));
    Odrv4 I__1501 (
            .O(N__14513),
            .I(\b2v_inst.un1_state_36_0_sn ));
    CascadeMux I__1500 (
            .O(N__14510),
            .I(\b2v_inst.N_325_cascade_ ));
    InMux I__1499 (
            .O(N__14507),
            .I(\b2v_inst.un1_indice_cry_6 ));
    InMux I__1498 (
            .O(N__14504),
            .I(\b2v_inst.un1_indice_cry_7 ));
    InMux I__1497 (
            .O(N__14501),
            .I(bfn_6_7_0_));
    InMux I__1496 (
            .O(N__14498),
            .I(\b2v_inst.un1_indice_cry_9 ));
    InMux I__1495 (
            .O(N__14495),
            .I(\b2v_inst.un1_indice_cry_10 ));
    InMux I__1494 (
            .O(N__14492),
            .I(N__14489));
    LocalMux I__1493 (
            .O(N__14489),
            .I(\b2v_inst.ignorar_ancho_1_RNOZ0Z_1 ));
    InMux I__1492 (
            .O(N__14486),
            .I(N__14483));
    LocalMux I__1491 (
            .O(N__14483),
            .I(\b2v_inst.ignorar_ancho_1_RNOZ0Z_2 ));
    InMux I__1490 (
            .O(N__14480),
            .I(\b2v_inst.un2_dir_mem_3_cry_2 ));
    InMux I__1489 (
            .O(N__14477),
            .I(\b2v_inst.un2_dir_mem_3_cry_3 ));
    InMux I__1488 (
            .O(N__14474),
            .I(\b2v_inst.un2_dir_mem_3_cry_4 ));
    InMux I__1487 (
            .O(N__14471),
            .I(\b2v_inst.un1_indice_cry_1 ));
    InMux I__1486 (
            .O(N__14468),
            .I(\b2v_inst.un1_indice_cry_2 ));
    InMux I__1485 (
            .O(N__14465),
            .I(\b2v_inst.un1_indice_cry_3 ));
    InMux I__1484 (
            .O(N__14462),
            .I(\b2v_inst.un1_indice_cry_4 ));
    InMux I__1483 (
            .O(N__14459),
            .I(\b2v_inst.un1_indice_cry_5 ));
    InMux I__1482 (
            .O(N__14456),
            .I(\b2v_inst4.un1_pix_count_int_cry_18 ));
    CascadeMux I__1481 (
            .O(N__14453),
            .I(N__14449));
    CascadeMux I__1480 (
            .O(N__14452),
            .I(N__14446));
    CascadeBuf I__1479 (
            .O(N__14449),
            .I(N__14443));
    CascadeBuf I__1478 (
            .O(N__14446),
            .I(N__14440));
    CascadeMux I__1477 (
            .O(N__14443),
            .I(N__14437));
    CascadeMux I__1476 (
            .O(N__14440),
            .I(N__14434));
    CascadeBuf I__1475 (
            .O(N__14437),
            .I(N__14431));
    CascadeBuf I__1474 (
            .O(N__14434),
            .I(N__14428));
    CascadeMux I__1473 (
            .O(N__14431),
            .I(N__14425));
    CascadeMux I__1472 (
            .O(N__14428),
            .I(N__14422));
    CascadeBuf I__1471 (
            .O(N__14425),
            .I(N__14419));
    CascadeBuf I__1470 (
            .O(N__14422),
            .I(N__14416));
    CascadeMux I__1469 (
            .O(N__14419),
            .I(N__14413));
    CascadeMux I__1468 (
            .O(N__14416),
            .I(N__14410));
    CascadeBuf I__1467 (
            .O(N__14413),
            .I(N__14407));
    CascadeBuf I__1466 (
            .O(N__14410),
            .I(N__14404));
    CascadeMux I__1465 (
            .O(N__14407),
            .I(N__14401));
    CascadeMux I__1464 (
            .O(N__14404),
            .I(N__14398));
    CascadeBuf I__1463 (
            .O(N__14401),
            .I(N__14395));
    CascadeBuf I__1462 (
            .O(N__14398),
            .I(N__14392));
    CascadeMux I__1461 (
            .O(N__14395),
            .I(N__14389));
    CascadeMux I__1460 (
            .O(N__14392),
            .I(N__14386));
    CascadeBuf I__1459 (
            .O(N__14389),
            .I(N__14383));
    CascadeBuf I__1458 (
            .O(N__14386),
            .I(N__14380));
    CascadeMux I__1457 (
            .O(N__14383),
            .I(N__14377));
    CascadeMux I__1456 (
            .O(N__14380),
            .I(N__14374));
    InMux I__1455 (
            .O(N__14377),
            .I(N__14371));
    InMux I__1454 (
            .O(N__14374),
            .I(N__14368));
    LocalMux I__1453 (
            .O(N__14371),
            .I(N__14365));
    LocalMux I__1452 (
            .O(N__14368),
            .I(SYNTHESIZED_WIRE_12_1));
    Odrv4 I__1451 (
            .O(N__14365),
            .I(SYNTHESIZED_WIRE_12_1));
    CascadeMux I__1450 (
            .O(N__14360),
            .I(N__14357));
    CascadeBuf I__1449 (
            .O(N__14357),
            .I(N__14353));
    CascadeMux I__1448 (
            .O(N__14356),
            .I(N__14350));
    CascadeMux I__1447 (
            .O(N__14353),
            .I(N__14347));
    CascadeBuf I__1446 (
            .O(N__14350),
            .I(N__14344));
    CascadeBuf I__1445 (
            .O(N__14347),
            .I(N__14341));
    CascadeMux I__1444 (
            .O(N__14344),
            .I(N__14338));
    CascadeMux I__1443 (
            .O(N__14341),
            .I(N__14335));
    CascadeBuf I__1442 (
            .O(N__14338),
            .I(N__14332));
    CascadeBuf I__1441 (
            .O(N__14335),
            .I(N__14329));
    CascadeMux I__1440 (
            .O(N__14332),
            .I(N__14326));
    CascadeMux I__1439 (
            .O(N__14329),
            .I(N__14323));
    CascadeBuf I__1438 (
            .O(N__14326),
            .I(N__14320));
    CascadeBuf I__1437 (
            .O(N__14323),
            .I(N__14317));
    CascadeMux I__1436 (
            .O(N__14320),
            .I(N__14314));
    CascadeMux I__1435 (
            .O(N__14317),
            .I(N__14311));
    CascadeBuf I__1434 (
            .O(N__14314),
            .I(N__14308));
    CascadeBuf I__1433 (
            .O(N__14311),
            .I(N__14305));
    CascadeMux I__1432 (
            .O(N__14308),
            .I(N__14302));
    CascadeMux I__1431 (
            .O(N__14305),
            .I(N__14299));
    CascadeBuf I__1430 (
            .O(N__14302),
            .I(N__14296));
    CascadeBuf I__1429 (
            .O(N__14299),
            .I(N__14293));
    CascadeMux I__1428 (
            .O(N__14296),
            .I(N__14290));
    CascadeMux I__1427 (
            .O(N__14293),
            .I(N__14287));
    CascadeBuf I__1426 (
            .O(N__14290),
            .I(N__14284));
    InMux I__1425 (
            .O(N__14287),
            .I(N__14281));
    CascadeMux I__1424 (
            .O(N__14284),
            .I(N__14278));
    LocalMux I__1423 (
            .O(N__14281),
            .I(N__14275));
    InMux I__1422 (
            .O(N__14278),
            .I(N__14272));
    Span4Mux_h I__1421 (
            .O(N__14275),
            .I(N__14269));
    LocalMux I__1420 (
            .O(N__14272),
            .I(SYNTHESIZED_WIRE_12_7));
    Odrv4 I__1419 (
            .O(N__14269),
            .I(SYNTHESIZED_WIRE_12_7));
    CascadeMux I__1418 (
            .O(N__14264),
            .I(N__14260));
    CascadeMux I__1417 (
            .O(N__14263),
            .I(N__14257));
    CascadeBuf I__1416 (
            .O(N__14260),
            .I(N__14254));
    CascadeBuf I__1415 (
            .O(N__14257),
            .I(N__14251));
    CascadeMux I__1414 (
            .O(N__14254),
            .I(N__14248));
    CascadeMux I__1413 (
            .O(N__14251),
            .I(N__14245));
    CascadeBuf I__1412 (
            .O(N__14248),
            .I(N__14242));
    CascadeBuf I__1411 (
            .O(N__14245),
            .I(N__14239));
    CascadeMux I__1410 (
            .O(N__14242),
            .I(N__14236));
    CascadeMux I__1409 (
            .O(N__14239),
            .I(N__14233));
    CascadeBuf I__1408 (
            .O(N__14236),
            .I(N__14230));
    CascadeBuf I__1407 (
            .O(N__14233),
            .I(N__14227));
    CascadeMux I__1406 (
            .O(N__14230),
            .I(N__14224));
    CascadeMux I__1405 (
            .O(N__14227),
            .I(N__14221));
    CascadeBuf I__1404 (
            .O(N__14224),
            .I(N__14218));
    CascadeBuf I__1403 (
            .O(N__14221),
            .I(N__14215));
    CascadeMux I__1402 (
            .O(N__14218),
            .I(N__14212));
    CascadeMux I__1401 (
            .O(N__14215),
            .I(N__14209));
    CascadeBuf I__1400 (
            .O(N__14212),
            .I(N__14206));
    CascadeBuf I__1399 (
            .O(N__14209),
            .I(N__14203));
    CascadeMux I__1398 (
            .O(N__14206),
            .I(N__14200));
    CascadeMux I__1397 (
            .O(N__14203),
            .I(N__14197));
    CascadeBuf I__1396 (
            .O(N__14200),
            .I(N__14194));
    CascadeBuf I__1395 (
            .O(N__14197),
            .I(N__14191));
    CascadeMux I__1394 (
            .O(N__14194),
            .I(N__14188));
    CascadeMux I__1393 (
            .O(N__14191),
            .I(N__14185));
    InMux I__1392 (
            .O(N__14188),
            .I(N__14182));
    InMux I__1391 (
            .O(N__14185),
            .I(N__14179));
    LocalMux I__1390 (
            .O(N__14182),
            .I(N__14176));
    LocalMux I__1389 (
            .O(N__14179),
            .I(SYNTHESIZED_WIRE_12_0));
    Odrv4 I__1388 (
            .O(N__14176),
            .I(SYNTHESIZED_WIRE_12_0));
    CascadeMux I__1387 (
            .O(N__14171),
            .I(N__14167));
    CascadeMux I__1386 (
            .O(N__14170),
            .I(N__14164));
    CascadeBuf I__1385 (
            .O(N__14167),
            .I(N__14161));
    CascadeBuf I__1384 (
            .O(N__14164),
            .I(N__14158));
    CascadeMux I__1383 (
            .O(N__14161),
            .I(N__14155));
    CascadeMux I__1382 (
            .O(N__14158),
            .I(N__14152));
    CascadeBuf I__1381 (
            .O(N__14155),
            .I(N__14149));
    CascadeBuf I__1380 (
            .O(N__14152),
            .I(N__14146));
    CascadeMux I__1379 (
            .O(N__14149),
            .I(N__14143));
    CascadeMux I__1378 (
            .O(N__14146),
            .I(N__14140));
    CascadeBuf I__1377 (
            .O(N__14143),
            .I(N__14137));
    CascadeBuf I__1376 (
            .O(N__14140),
            .I(N__14134));
    CascadeMux I__1375 (
            .O(N__14137),
            .I(N__14131));
    CascadeMux I__1374 (
            .O(N__14134),
            .I(N__14128));
    CascadeBuf I__1373 (
            .O(N__14131),
            .I(N__14125));
    CascadeBuf I__1372 (
            .O(N__14128),
            .I(N__14122));
    CascadeMux I__1371 (
            .O(N__14125),
            .I(N__14119));
    CascadeMux I__1370 (
            .O(N__14122),
            .I(N__14116));
    CascadeBuf I__1369 (
            .O(N__14119),
            .I(N__14113));
    CascadeBuf I__1368 (
            .O(N__14116),
            .I(N__14110));
    CascadeMux I__1367 (
            .O(N__14113),
            .I(N__14107));
    CascadeMux I__1366 (
            .O(N__14110),
            .I(N__14104));
    CascadeBuf I__1365 (
            .O(N__14107),
            .I(N__14101));
    CascadeBuf I__1364 (
            .O(N__14104),
            .I(N__14098));
    CascadeMux I__1363 (
            .O(N__14101),
            .I(N__14095));
    CascadeMux I__1362 (
            .O(N__14098),
            .I(N__14092));
    InMux I__1361 (
            .O(N__14095),
            .I(N__14089));
    InMux I__1360 (
            .O(N__14092),
            .I(N__14086));
    LocalMux I__1359 (
            .O(N__14089),
            .I(SYNTHESIZED_WIRE_12_8));
    LocalMux I__1358 (
            .O(N__14086),
            .I(SYNTHESIZED_WIRE_12_8));
    InMux I__1357 (
            .O(N__14081),
            .I(\b2v_inst.un2_dir_mem_3_cry_0 ));
    InMux I__1356 (
            .O(N__14078),
            .I(\b2v_inst.un2_dir_mem_3_cry_1 ));
    InMux I__1355 (
            .O(N__14075),
            .I(\b2v_inst4.un1_pix_count_int_cry_9 ));
    InMux I__1354 (
            .O(N__14072),
            .I(\b2v_inst4.un1_pix_count_int_cry_10 ));
    InMux I__1353 (
            .O(N__14069),
            .I(N__14063));
    InMux I__1352 (
            .O(N__14068),
            .I(N__14063));
    LocalMux I__1351 (
            .O(N__14063),
            .I(N__14060));
    Odrv4 I__1350 (
            .O(N__14060),
            .I(\b2v_inst4.un1_pix_count_int_cry_11_c_RNIMPVJZ0 ));
    InMux I__1349 (
            .O(N__14057),
            .I(\b2v_inst4.un1_pix_count_int_cry_11 ));
    InMux I__1348 (
            .O(N__14054),
            .I(\b2v_inst4.un1_pix_count_int_cry_12 ));
    InMux I__1347 (
            .O(N__14051),
            .I(\b2v_inst4.un1_pix_count_int_cry_13 ));
    InMux I__1346 (
            .O(N__14048),
            .I(\b2v_inst4.un1_pix_count_int_cry_14 ));
    InMux I__1345 (
            .O(N__14045),
            .I(bfn_5_15_0_));
    InMux I__1344 (
            .O(N__14042),
            .I(\b2v_inst4.un1_pix_count_int_cry_16 ));
    InMux I__1343 (
            .O(N__14039),
            .I(\b2v_inst4.un1_pix_count_int_cry_17 ));
    InMux I__1342 (
            .O(N__14036),
            .I(N__14033));
    LocalMux I__1341 (
            .O(N__14033),
            .I(N__14029));
    InMux I__1340 (
            .O(N__14032),
            .I(N__14026));
    Span4Mux_v I__1339 (
            .O(N__14029),
            .I(N__14021));
    LocalMux I__1338 (
            .O(N__14026),
            .I(N__14021));
    Span4Mux_h I__1337 (
            .O(N__14021),
            .I(N__14018));
    Odrv4 I__1336 (
            .O(N__14018),
            .I(\b2v_inst4.un1_pix_count_int_cry_0_c_RNIIC2IZ0 ));
    InMux I__1335 (
            .O(N__14015),
            .I(\b2v_inst4.un1_pix_count_int_cry_0 ));
    InMux I__1334 (
            .O(N__14012),
            .I(N__14009));
    LocalMux I__1333 (
            .O(N__14009),
            .I(N__14005));
    InMux I__1332 (
            .O(N__14008),
            .I(N__14002));
    Span4Mux_v I__1331 (
            .O(N__14005),
            .I(N__13997));
    LocalMux I__1330 (
            .O(N__14002),
            .I(N__13997));
    Span4Mux_h I__1329 (
            .O(N__13997),
            .I(N__13994));
    Odrv4 I__1328 (
            .O(N__13994),
            .I(\b2v_inst4.un1_pix_count_int_cry_1_c_RNIKF3IZ0 ));
    InMux I__1327 (
            .O(N__13991),
            .I(\b2v_inst4.un1_pix_count_int_cry_1 ));
    InMux I__1326 (
            .O(N__13988),
            .I(N__13982));
    InMux I__1325 (
            .O(N__13987),
            .I(N__13982));
    LocalMux I__1324 (
            .O(N__13982),
            .I(N__13979));
    Odrv12 I__1323 (
            .O(N__13979),
            .I(\b2v_inst4.un1_pix_count_int_cry_2_c_RNIMI4IZ0 ));
    InMux I__1322 (
            .O(N__13976),
            .I(\b2v_inst4.un1_pix_count_int_cry_2 ));
    InMux I__1321 (
            .O(N__13973),
            .I(\b2v_inst4.un1_pix_count_int_cry_3 ));
    InMux I__1320 (
            .O(N__13970),
            .I(N__13964));
    InMux I__1319 (
            .O(N__13969),
            .I(N__13964));
    LocalMux I__1318 (
            .O(N__13964),
            .I(N__13961));
    Span4Mux_h I__1317 (
            .O(N__13961),
            .I(N__13958));
    Odrv4 I__1316 (
            .O(N__13958),
            .I(\b2v_inst4.un1_pix_count_int_cry_4_c_RNIQO6IZ0 ));
    InMux I__1315 (
            .O(N__13955),
            .I(\b2v_inst4.un1_pix_count_int_cry_4 ));
    InMux I__1314 (
            .O(N__13952),
            .I(N__13949));
    LocalMux I__1313 (
            .O(N__13949),
            .I(N__13945));
    InMux I__1312 (
            .O(N__13948),
            .I(N__13942));
    Span4Mux_v I__1311 (
            .O(N__13945),
            .I(N__13937));
    LocalMux I__1310 (
            .O(N__13942),
            .I(N__13937));
    Span4Mux_h I__1309 (
            .O(N__13937),
            .I(N__13934));
    Odrv4 I__1308 (
            .O(N__13934),
            .I(\b2v_inst4.un1_pix_count_int_cry_5_c_RNISR7IZ0 ));
    InMux I__1307 (
            .O(N__13931),
            .I(\b2v_inst4.un1_pix_count_int_cry_5 ));
    InMux I__1306 (
            .O(N__13928),
            .I(\b2v_inst4.un1_pix_count_int_cry_6 ));
    InMux I__1305 (
            .O(N__13925),
            .I(bfn_5_14_0_));
    InMux I__1304 (
            .O(N__13922),
            .I(\b2v_inst4.un1_pix_count_int_cry_8 ));
    CascadeMux I__1303 (
            .O(N__13919),
            .I(N__13915));
    InMux I__1302 (
            .O(N__13918),
            .I(N__13907));
    InMux I__1301 (
            .O(N__13915),
            .I(N__13907));
    InMux I__1300 (
            .O(N__13914),
            .I(N__13907));
    LocalMux I__1299 (
            .O(N__13907),
            .I(N__13904));
    Odrv12 I__1298 (
            .O(N__13904),
            .I(\b2v_inst.un1_cuenta_pixel_cry_3_c_RNICFVHZ0 ));
    CascadeMux I__1297 (
            .O(N__13901),
            .I(N__13898));
    InMux I__1296 (
            .O(N__13898),
            .I(N__13895));
    LocalMux I__1295 (
            .O(N__13895),
            .I(N__13892));
    Odrv4 I__1294 (
            .O(N__13892),
            .I(\b2v_inst.cuenta_pixelZ0Z_4 ));
    CascadeMux I__1293 (
            .O(N__13889),
            .I(N__13886));
    InMux I__1292 (
            .O(N__13886),
            .I(N__13883));
    LocalMux I__1291 (
            .O(N__13883),
            .I(N__13880));
    Odrv12 I__1290 (
            .O(N__13880),
            .I(\b2v_inst.un7_pix_count_int_0_I_9_c_RNOZ0 ));
    InMux I__1289 (
            .O(N__13877),
            .I(N__13874));
    LocalMux I__1288 (
            .O(N__13874),
            .I(\b2v_inst.pix_count_anteriorZ0Z_10 ));
    CascadeMux I__1287 (
            .O(N__13871),
            .I(N__13868));
    InMux I__1286 (
            .O(N__13868),
            .I(N__13865));
    LocalMux I__1285 (
            .O(N__13865),
            .I(\b2v_inst.pix_count_anteriorZ0Z_11 ));
    InMux I__1284 (
            .O(N__13862),
            .I(N__13859));
    LocalMux I__1283 (
            .O(N__13859),
            .I(N__13856));
    Odrv4 I__1282 (
            .O(N__13856),
            .I(\b2v_inst.pix_count_anteriorZ0Z_17 ));
    CEMux I__1281 (
            .O(N__13853),
            .I(N__13823));
    CEMux I__1280 (
            .O(N__13852),
            .I(N__13823));
    CEMux I__1279 (
            .O(N__13851),
            .I(N__13823));
    CEMux I__1278 (
            .O(N__13850),
            .I(N__13823));
    CEMux I__1277 (
            .O(N__13849),
            .I(N__13823));
    CEMux I__1276 (
            .O(N__13848),
            .I(N__13823));
    CEMux I__1275 (
            .O(N__13847),
            .I(N__13823));
    CEMux I__1274 (
            .O(N__13846),
            .I(N__13823));
    CEMux I__1273 (
            .O(N__13845),
            .I(N__13823));
    CEMux I__1272 (
            .O(N__13844),
            .I(N__13823));
    GlobalMux I__1271 (
            .O(N__13823),
            .I(N__13820));
    gio2CtrlBuf I__1270 (
            .O(N__13820),
            .I(\b2v_inst.N_305_1_g ));
    InMux I__1269 (
            .O(N__13817),
            .I(N__13814));
    LocalMux I__1268 (
            .O(N__13814),
            .I(N__13811));
    Odrv4 I__1267 (
            .O(N__13811),
            .I(\b2v_inst.N_4_i_i_a6_1 ));
    InMux I__1266 (
            .O(N__13808),
            .I(N__13805));
    LocalMux I__1265 (
            .O(N__13805),
            .I(N__13802));
    Span4Mux_v I__1264 (
            .O(N__13802),
            .I(N__13798));
    InMux I__1263 (
            .O(N__13801),
            .I(N__13795));
    Sp12to4 I__1262 (
            .O(N__13798),
            .I(N__13790));
    LocalMux I__1261 (
            .O(N__13795),
            .I(N__13790));
    Odrv12 I__1260 (
            .O(N__13790),
            .I(\b2v_inst4.pix_count_int_RNI0EPTZ0Z_0 ));
    InMux I__1259 (
            .O(N__13787),
            .I(N__13784));
    LocalMux I__1258 (
            .O(N__13784),
            .I(\b2v_inst4.un1_pix_count_int_0_sqmuxa_10 ));
    InMux I__1257 (
            .O(N__13781),
            .I(N__13778));
    LocalMux I__1256 (
            .O(N__13778),
            .I(N__13775));
    Span4Mux_v I__1255 (
            .O(N__13775),
            .I(N__13771));
    InMux I__1254 (
            .O(N__13774),
            .I(N__13768));
    Span4Mux_h I__1253 (
            .O(N__13771),
            .I(N__13763));
    LocalMux I__1252 (
            .O(N__13768),
            .I(N__13763));
    Odrv4 I__1251 (
            .O(N__13763),
            .I(\b2v_inst.cuenta_pixel_RNIT0FMZ0Z_1 ));
    InMux I__1250 (
            .O(N__13760),
            .I(N__13755));
    InMux I__1249 (
            .O(N__13759),
            .I(N__13752));
    CascadeMux I__1248 (
            .O(N__13758),
            .I(N__13749));
    LocalMux I__1247 (
            .O(N__13755),
            .I(N__13744));
    LocalMux I__1246 (
            .O(N__13752),
            .I(N__13740));
    InMux I__1245 (
            .O(N__13749),
            .I(N__13737));
    InMux I__1244 (
            .O(N__13748),
            .I(N__13732));
    InMux I__1243 (
            .O(N__13747),
            .I(N__13732));
    Span4Mux_h I__1242 (
            .O(N__13744),
            .I(N__13729));
    InMux I__1241 (
            .O(N__13743),
            .I(N__13726));
    Span4Mux_h I__1240 (
            .O(N__13740),
            .I(N__13721));
    LocalMux I__1239 (
            .O(N__13737),
            .I(N__13721));
    LocalMux I__1238 (
            .O(N__13732),
            .I(\b2v_inst.cuenta_pixelZ0Z_0 ));
    Odrv4 I__1237 (
            .O(N__13729),
            .I(\b2v_inst.cuenta_pixelZ0Z_0 ));
    LocalMux I__1236 (
            .O(N__13726),
            .I(\b2v_inst.cuenta_pixelZ0Z_0 ));
    Odrv4 I__1235 (
            .O(N__13721),
            .I(\b2v_inst.cuenta_pixelZ0Z_0 ));
    CascadeMux I__1234 (
            .O(N__13712),
            .I(\b2v_inst.cuenta_pixel_5_i_a2_0_2_5_cascade_ ));
    InMux I__1233 (
            .O(N__13709),
            .I(N__13706));
    LocalMux I__1232 (
            .O(N__13706),
            .I(N__13703));
    Odrv4 I__1231 (
            .O(N__13703),
            .I(\b2v_inst.cuenta_pixelZ0Z_2 ));
    InMux I__1230 (
            .O(N__13700),
            .I(N__13697));
    LocalMux I__1229 (
            .O(N__13697),
            .I(N__13694));
    Odrv4 I__1228 (
            .O(N__13694),
            .I(\b2v_inst.cuenta_pixelZ0Z_3 ));
    InMux I__1227 (
            .O(N__13691),
            .I(N__13682));
    InMux I__1226 (
            .O(N__13690),
            .I(N__13682));
    InMux I__1225 (
            .O(N__13689),
            .I(N__13682));
    LocalMux I__1224 (
            .O(N__13682),
            .I(N__13679));
    Odrv4 I__1223 (
            .O(N__13679),
            .I(\b2v_inst.un1_cuenta_pixel_cry_1_c_RNI89THZ0 ));
    CascadeMux I__1222 (
            .O(N__13676),
            .I(N__13672));
    InMux I__1221 (
            .O(N__13675),
            .I(N__13664));
    InMux I__1220 (
            .O(N__13672),
            .I(N__13664));
    InMux I__1219 (
            .O(N__13671),
            .I(N__13664));
    LocalMux I__1218 (
            .O(N__13664),
            .I(N__13661));
    Odrv12 I__1217 (
            .O(N__13661),
            .I(\b2v_inst.un1_cuenta_pixel_cry_2_c_RNIACUHZ0 ));
    InMux I__1216 (
            .O(N__13658),
            .I(N__13652));
    InMux I__1215 (
            .O(N__13657),
            .I(N__13645));
    InMux I__1214 (
            .O(N__13656),
            .I(N__13645));
    InMux I__1213 (
            .O(N__13655),
            .I(N__13645));
    LocalMux I__1212 (
            .O(N__13652),
            .I(N__13642));
    LocalMux I__1211 (
            .O(N__13645),
            .I(N__13639));
    Odrv4 I__1210 (
            .O(N__13642),
            .I(\b2v_inst.un1_cuenta_pixel_cry_4_c_RNIEI0IZ0 ));
    Odrv4 I__1209 (
            .O(N__13639),
            .I(\b2v_inst.un1_cuenta_pixel_cry_4_c_RNIEI0IZ0 ));
    InMux I__1208 (
            .O(N__13634),
            .I(N__13631));
    LocalMux I__1207 (
            .O(N__13631),
            .I(N__13627));
    InMux I__1206 (
            .O(N__13630),
            .I(N__13624));
    Span4Mux_h I__1205 (
            .O(N__13627),
            .I(N__13621));
    LocalMux I__1204 (
            .O(N__13624),
            .I(\b2v_inst.cuenta_pixel_5_i_a2_0_2_5 ));
    Odrv4 I__1203 (
            .O(N__13621),
            .I(\b2v_inst.cuenta_pixel_5_i_a2_0_2_5 ));
    InMux I__1202 (
            .O(N__13616),
            .I(N__13613));
    LocalMux I__1201 (
            .O(N__13613),
            .I(N__13609));
    CascadeMux I__1200 (
            .O(N__13612),
            .I(N__13606));
    Span4Mux_v I__1199 (
            .O(N__13609),
            .I(N__13602));
    InMux I__1198 (
            .O(N__13606),
            .I(N__13597));
    InMux I__1197 (
            .O(N__13605),
            .I(N__13597));
    Odrv4 I__1196 (
            .O(N__13602),
            .I(\b2v_inst.cuenta_pixel_5_i_a2_0_1_5 ));
    LocalMux I__1195 (
            .O(N__13597),
            .I(\b2v_inst.cuenta_pixel_5_i_a2_0_1_5 ));
    CascadeMux I__1194 (
            .O(N__13592),
            .I(N__13589));
    InMux I__1193 (
            .O(N__13589),
            .I(N__13586));
    LocalMux I__1192 (
            .O(N__13586),
            .I(N__13583));
    Odrv4 I__1191 (
            .O(N__13583),
            .I(\b2v_inst.cuenta_pixelZ0Z_5 ));
    InMux I__1190 (
            .O(N__13580),
            .I(N__13577));
    LocalMux I__1189 (
            .O(N__13577),
            .I(N__13574));
    Odrv4 I__1188 (
            .O(N__13574),
            .I(\b2v_inst4.un1_pix_count_int_0_sqmuxa_7 ));
    InMux I__1187 (
            .O(N__13571),
            .I(N__13568));
    LocalMux I__1186 (
            .O(N__13568),
            .I(\b2v_inst4.un1_pix_count_int_0_sqmuxa_13 ));
    CascadeMux I__1185 (
            .O(N__13565),
            .I(\b2v_inst4.un1_pix_count_int_0_sqmuxa_8_cascade_ ));
    InMux I__1184 (
            .O(N__13562),
            .I(N__13559));
    LocalMux I__1183 (
            .O(N__13559),
            .I(\b2v_inst4.un1_pix_count_int_0_sqmuxa_14 ));
    InMux I__1182 (
            .O(N__13556),
            .I(N__13553));
    LocalMux I__1181 (
            .O(N__13553),
            .I(N__13550));
    Span4Mux_v I__1180 (
            .O(N__13550),
            .I(N__13547));
    Odrv4 I__1179 (
            .O(N__13547),
            .I(\b2v_inst.pix_count_anteriorZ0Z_9 ));
    CascadeMux I__1178 (
            .O(N__13544),
            .I(N__13541));
    InMux I__1177 (
            .O(N__13541),
            .I(N__13538));
    LocalMux I__1176 (
            .O(N__13538),
            .I(\b2v_inst.un7_pix_count_int_0_I_51_c_RNOZ0 ));
    CascadeMux I__1175 (
            .O(N__13535),
            .I(\b2v_inst.N_1_0_0_cascade_ ));
    CascadeMux I__1174 (
            .O(N__13532),
            .I(\b2v_inst.N_4_i_i_o6_2_cascade_ ));
    InMux I__1173 (
            .O(N__13529),
            .I(N__13526));
    LocalMux I__1172 (
            .O(N__13526),
            .I(N__13523));
    Span4Mux_h I__1171 (
            .O(N__13523),
            .I(N__13520));
    Odrv4 I__1170 (
            .O(N__13520),
            .I(\b2v_inst.N_7 ));
    CascadeMux I__1169 (
            .O(N__13517),
            .I(N__13514));
    InMux I__1168 (
            .O(N__13514),
            .I(N__13511));
    LocalMux I__1167 (
            .O(N__13511),
            .I(N__13508));
    Odrv4 I__1166 (
            .O(N__13508),
            .I(\b2v_inst.un7_pix_count_int_0_I_21_c_RNOZ0 ));
    InMux I__1165 (
            .O(N__13505),
            .I(N__13502));
    LocalMux I__1164 (
            .O(N__13502),
            .I(\b2v_inst.pix_count_anteriorZ0Z_6 ));
    InMux I__1163 (
            .O(N__13499),
            .I(N__13496));
    LocalMux I__1162 (
            .O(N__13496),
            .I(\b2v_inst.pix_count_anteriorZ0Z_7 ));
    CascadeMux I__1161 (
            .O(N__13493),
            .I(N__13490));
    InMux I__1160 (
            .O(N__13490),
            .I(N__13487));
    LocalMux I__1159 (
            .O(N__13487),
            .I(\b2v_inst.pix_count_anteriorZ0Z_8 ));
    InMux I__1158 (
            .O(N__13484),
            .I(\b2v_inst.un1_cuenta_pixel_cry_3 ));
    InMux I__1157 (
            .O(N__13481),
            .I(\b2v_inst.un1_cuenta_pixel_cry_4 ));
    InMux I__1156 (
            .O(N__13478),
            .I(N__13475));
    LocalMux I__1155 (
            .O(N__13475),
            .I(N__13472));
    Odrv4 I__1154 (
            .O(N__13472),
            .I(\b2v_inst.cuenta_pixelZ0Z_6 ));
    InMux I__1153 (
            .O(N__13469),
            .I(N__13466));
    LocalMux I__1152 (
            .O(N__13466),
            .I(N__13462));
    InMux I__1151 (
            .O(N__13465),
            .I(N__13459));
    Odrv4 I__1150 (
            .O(N__13462),
            .I(\b2v_inst.un1_cuenta_pixel_cry_5_c_RNIGL1IZ0 ));
    LocalMux I__1149 (
            .O(N__13459),
            .I(\b2v_inst.un1_cuenta_pixel_cry_5_c_RNIGL1IZ0 ));
    InMux I__1148 (
            .O(N__13454),
            .I(\b2v_inst.un1_cuenta_pixel_cry_5 ));
    InMux I__1147 (
            .O(N__13451),
            .I(N__13448));
    LocalMux I__1146 (
            .O(N__13448),
            .I(\b2v_inst.cuenta_pixelZ0Z_7 ));
    InMux I__1145 (
            .O(N__13445),
            .I(N__13441));
    InMux I__1144 (
            .O(N__13444),
            .I(N__13438));
    LocalMux I__1143 (
            .O(N__13441),
            .I(\b2v_inst.un1_cuenta_pixel_cry_6_c_RNIIO2IZ0 ));
    LocalMux I__1142 (
            .O(N__13438),
            .I(\b2v_inst.un1_cuenta_pixel_cry_6_c_RNIIO2IZ0 ));
    InMux I__1141 (
            .O(N__13433),
            .I(\b2v_inst.un1_cuenta_pixel_cry_6 ));
    InMux I__1140 (
            .O(N__13430),
            .I(N__13427));
    LocalMux I__1139 (
            .O(N__13427),
            .I(\b2v_inst.cuenta_pixelZ0Z_8 ));
    InMux I__1138 (
            .O(N__13424),
            .I(\b2v_inst.un1_cuenta_pixel_cry_7 ));
    InMux I__1137 (
            .O(N__13421),
            .I(N__13418));
    LocalMux I__1136 (
            .O(N__13418),
            .I(N__13415));
    Odrv12 I__1135 (
            .O(N__13415),
            .I(\b2v_inst.cuenta_pixelZ0Z_9 ));
    InMux I__1134 (
            .O(N__13412),
            .I(bfn_3_11_0_));
    InMux I__1133 (
            .O(N__13409),
            .I(\b2v_inst.un1_cuenta_pixel_cry_9 ));
    InMux I__1132 (
            .O(N__13406),
            .I(N__13403));
    LocalMux I__1131 (
            .O(N__13403),
            .I(\b2v_inst.cuenta_pixelZ0Z_10 ));
    CascadeMux I__1130 (
            .O(N__13400),
            .I(\b2v_inst.un1_state_36_0_a2_0_2_1_cascade_ ));
    InMux I__1129 (
            .O(N__13397),
            .I(N__13394));
    LocalMux I__1128 (
            .O(N__13394),
            .I(N__13389));
    InMux I__1127 (
            .O(N__13393),
            .I(N__13384));
    InMux I__1126 (
            .O(N__13392),
            .I(N__13384));
    Odrv4 I__1125 (
            .O(N__13389),
            .I(\b2v_inst.N_305_2 ));
    LocalMux I__1124 (
            .O(N__13384),
            .I(\b2v_inst.N_305_2 ));
    CascadeMux I__1123 (
            .O(N__13379),
            .I(\b2v_inst.N_305_2_cascade_ ));
    InMux I__1122 (
            .O(N__13376),
            .I(N__13371));
    InMux I__1121 (
            .O(N__13375),
            .I(N__13368));
    InMux I__1120 (
            .O(N__13374),
            .I(N__13365));
    LocalMux I__1119 (
            .O(N__13371),
            .I(N__13362));
    LocalMux I__1118 (
            .O(N__13368),
            .I(\b2v_inst.cuenta_pixelZ0Z_1 ));
    LocalMux I__1117 (
            .O(N__13365),
            .I(\b2v_inst.cuenta_pixelZ0Z_1 ));
    Odrv4 I__1116 (
            .O(N__13362),
            .I(\b2v_inst.cuenta_pixelZ0Z_1 ));
    InMux I__1115 (
            .O(N__13355),
            .I(\b2v_inst.un1_cuenta_pixel_cry_1 ));
    InMux I__1114 (
            .O(N__13352),
            .I(\b2v_inst.un1_cuenta_pixel_cry_2 ));
    InMux I__1113 (
            .O(N__13349),
            .I(N__13346));
    LocalMux I__1112 (
            .O(N__13346),
            .I(\b2v_inst.pix_count_anteriorZ0Z_13 ));
    CascadeMux I__1111 (
            .O(N__13343),
            .I(N__13340));
    InMux I__1110 (
            .O(N__13340),
            .I(N__13337));
    LocalMux I__1109 (
            .O(N__13337),
            .I(N__13334));
    Odrv4 I__1108 (
            .O(N__13334),
            .I(\b2v_inst.un7_pix_count_int_0_I_45_c_RNOZ0 ));
    CascadeMux I__1107 (
            .O(N__13331),
            .I(N__13328));
    InMux I__1106 (
            .O(N__13328),
            .I(N__13325));
    LocalMux I__1105 (
            .O(N__13325),
            .I(\b2v_inst.pix_count_anteriorZ0Z_14 ));
    CascadeMux I__1104 (
            .O(N__13322),
            .I(\b2v_inst4.un1_pix_count_int_0_sqmuxa_5_cascade_ ));
    InMux I__1103 (
            .O(N__13319),
            .I(N__13316));
    LocalMux I__1102 (
            .O(N__13316),
            .I(\b2v_inst.pix_count_anteriorZ0Z_15 ));
    CascadeMux I__1101 (
            .O(N__13313),
            .I(N__13310));
    InMux I__1100 (
            .O(N__13310),
            .I(N__13307));
    LocalMux I__1099 (
            .O(N__13307),
            .I(N__13304));
    Odrv4 I__1098 (
            .O(N__13304),
            .I(\b2v_inst.pix_count_anteriorZ0Z_19 ));
    CascadeMux I__1097 (
            .O(N__13301),
            .I(N__13298));
    InMux I__1096 (
            .O(N__13298),
            .I(N__13295));
    LocalMux I__1095 (
            .O(N__13295),
            .I(N__13292));
    Span4Mux_h I__1094 (
            .O(N__13292),
            .I(N__13289));
    Odrv4 I__1093 (
            .O(N__13289),
            .I(\b2v_inst.pix_count_anteriorZ0Z_16 ));
    InMux I__1092 (
            .O(N__13286),
            .I(N__13283));
    LocalMux I__1091 (
            .O(N__13283),
            .I(\b2v_inst.pix_count_anteriorZ0Z_2 ));
    CascadeMux I__1090 (
            .O(N__13280),
            .I(N__13277));
    InMux I__1089 (
            .O(N__13277),
            .I(N__13274));
    LocalMux I__1088 (
            .O(N__13274),
            .I(\b2v_inst.pix_count_anteriorZ0Z_3 ));
    InMux I__1087 (
            .O(N__13271),
            .I(N__13268));
    LocalMux I__1086 (
            .O(N__13268),
            .I(\b2v_inst.pix_count_anteriorZ0Z_0 ));
    InMux I__1085 (
            .O(N__13265),
            .I(N__13262));
    LocalMux I__1084 (
            .O(N__13262),
            .I(N__13259));
    Odrv4 I__1083 (
            .O(N__13259),
            .I(\b2v_inst.pix_count_anteriorZ0Z_5 ));
    CascadeMux I__1082 (
            .O(N__13256),
            .I(N__13253));
    InMux I__1081 (
            .O(N__13253),
            .I(N__13250));
    LocalMux I__1080 (
            .O(N__13250),
            .I(\b2v_inst.un7_pix_count_int_0_I_33_c_RNOZ0 ));
    InMux I__1079 (
            .O(N__13247),
            .I(N__13244));
    LocalMux I__1078 (
            .O(N__13244),
            .I(\b2v_inst.pix_count_anteriorZ0Z_18 ));
    CascadeMux I__1077 (
            .O(N__13241),
            .I(N__13238));
    InMux I__1076 (
            .O(N__13238),
            .I(N__13235));
    LocalMux I__1075 (
            .O(N__13235),
            .I(N__13232));
    Odrv4 I__1074 (
            .O(N__13232),
            .I(\b2v_inst.un7_pix_count_int_0_I_39_c_RNOZ0 ));
    CascadeMux I__1073 (
            .O(N__13229),
            .I(N__13226));
    InMux I__1072 (
            .O(N__13226),
            .I(N__13223));
    LocalMux I__1071 (
            .O(N__13223),
            .I(\b2v_inst.pix_count_anteriorZ0Z_12 ));
    InMux I__1070 (
            .O(N__13220),
            .I(\b2v_inst.un7_pix_count_int_0_N_2 ));
    CascadeMux I__1069 (
            .O(N__13217),
            .I(N__13214));
    InMux I__1068 (
            .O(N__13214),
            .I(N__13211));
    LocalMux I__1067 (
            .O(N__13211),
            .I(\b2v_inst.un7_pix_count_int_0_I_57_c_RNOZ0 ));
    InMux I__1066 (
            .O(N__13208),
            .I(N__13205));
    LocalMux I__1065 (
            .O(N__13205),
            .I(N__13202));
    Span4Mux_h I__1064 (
            .O(N__13202),
            .I(N__13199));
    Odrv4 I__1063 (
            .O(N__13199),
            .I(\b2v_inst4.un1_pix_count_int_0_sqmuxa_6 ));
    CascadeMux I__1062 (
            .O(N__13196),
            .I(N__13193));
    InMux I__1061 (
            .O(N__13193),
            .I(N__13190));
    LocalMux I__1060 (
            .O(N__13190),
            .I(N__13187));
    Odrv4 I__1059 (
            .O(N__13187),
            .I(\b2v_inst.un7_pix_count_int_0_I_27_c_RNOZ0 ));
    InMux I__1058 (
            .O(N__13184),
            .I(N__13181));
    LocalMux I__1057 (
            .O(N__13181),
            .I(\b2v_inst.pix_count_anteriorZ0Z_4 ));
    InMux I__1056 (
            .O(N__13178),
            .I(N__13175));
    LocalMux I__1055 (
            .O(N__13175),
            .I(\b2v_inst.un7_pix_count_int_0_I_1_c_RNOZ0 ));
    CascadeMux I__1054 (
            .O(N__13172),
            .I(N__13169));
    InMux I__1053 (
            .O(N__13169),
            .I(N__13166));
    LocalMux I__1052 (
            .O(N__13166),
            .I(\b2v_inst.un7_pix_count_int_0_I_15_c_RNOZ0 ));
    InMux I__1051 (
            .O(N__13163),
            .I(N__13156));
    InMux I__1050 (
            .O(N__13162),
            .I(N__13156));
    InMux I__1049 (
            .O(N__13161),
            .I(N__13153));
    LocalMux I__1048 (
            .O(N__13156),
            .I(b2v_inst4_pix_count_int_fast_0));
    LocalMux I__1047 (
            .O(N__13153),
            .I(b2v_inst4_pix_count_int_fast_0));
    InMux I__1046 (
            .O(N__13148),
            .I(N__13145));
    LocalMux I__1045 (
            .O(N__13145),
            .I(\b2v_inst.N_13 ));
    InMux I__1044 (
            .O(N__13142),
            .I(N__13133));
    InMux I__1043 (
            .O(N__13141),
            .I(N__13133));
    InMux I__1042 (
            .O(N__13140),
            .I(N__13133));
    LocalMux I__1041 (
            .O(N__13133),
            .I(b2v_inst4_pix_count_int_fast_2));
    CascadeMux I__1040 (
            .O(N__13130),
            .I(N__13126));
    CascadeMux I__1039 (
            .O(N__13129),
            .I(N__13122));
    InMux I__1038 (
            .O(N__13126),
            .I(N__13115));
    InMux I__1037 (
            .O(N__13125),
            .I(N__13115));
    InMux I__1036 (
            .O(N__13122),
            .I(N__13115));
    LocalMux I__1035 (
            .O(N__13115),
            .I(b2v_inst4_pix_count_int_fast_3));
    CascadeMux I__1034 (
            .O(N__13112),
            .I(N__13109));
    InMux I__1033 (
            .O(N__13109),
            .I(N__13106));
    LocalMux I__1032 (
            .O(N__13106),
            .I(N__13103));
    Odrv4 I__1031 (
            .O(N__13103),
            .I(\b2v_inst.pix_count_anteriorZ0Z_1 ));
    CascadeMux I__1030 (
            .O(N__13100),
            .I(\b2v_inst.un4_pix_count_intlto6_d_1_1_cascade_ ));
    InMux I__1029 (
            .O(N__13097),
            .I(N__13088));
    InMux I__1028 (
            .O(N__13096),
            .I(N__13088));
    InMux I__1027 (
            .O(N__13095),
            .I(N__13088));
    LocalMux I__1026 (
            .O(N__13088),
            .I(b2v_inst4_pix_count_int_fast_1));
    CascadeMux I__1025 (
            .O(N__13085),
            .I(\b2v_inst.N_4_i_i_a3_0_0_cascade_ ));
    defparam IN_MUX_bfv_17_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_13_0_));
    defparam IN_MUX_bfv_9_5_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_5_0_));
    defparam IN_MUX_bfv_9_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_6_0_ (
            .carryinitin(\b2v_inst.un8_dir_mem_2_cry_8 ),
            .carryinitout(bfn_9_6_0_));
    defparam IN_MUX_bfv_7_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_6_0_));
    defparam IN_MUX_bfv_7_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_7_0_ (
            .carryinitin(\b2v_inst.un8_dir_mem_1_cry_7 ),
            .carryinitout(bfn_7_7_0_));
    defparam IN_MUX_bfv_2_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_11_0_));
    defparam IN_MUX_bfv_2_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_12_0_ (
            .carryinitin(\b2v_inst.un7_pix_count_int_0_data_tmp_7 ),
            .carryinitout(bfn_2_12_0_));
    defparam IN_MUX_bfv_13_12_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_12_0_));
    defparam IN_MUX_bfv_13_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_13_0_ (
            .carryinitin(\b2v_inst.un4_cuenta_cry_8 ),
            .carryinitout(bfn_13_13_0_));
    defparam IN_MUX_bfv_8_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_9_0_));
    defparam IN_MUX_bfv_8_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_10_0_ (
            .carryinitin(\b2v_inst.un3_dir_mem_cry_7 ),
            .carryinitout(bfn_8_10_0_));
    defparam IN_MUX_bfv_6_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_5_0_));
    defparam IN_MUX_bfv_6_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_6_0_));
    defparam IN_MUX_bfv_6_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_7_0_ (
            .carryinitin(\b2v_inst.un1_indice_cry_8 ),
            .carryinitout(bfn_6_7_0_));
    defparam IN_MUX_bfv_3_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_10_0_));
    defparam IN_MUX_bfv_3_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_11_0_ (
            .carryinitin(\b2v_inst.un1_cuenta_pixel_cry_8 ),
            .carryinitout(bfn_3_11_0_));
    defparam IN_MUX_bfv_19_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_19_14_0_));
    defparam IN_MUX_bfv_17_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_8_0_));
    defparam IN_MUX_bfv_17_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_9_0_ (
            .carryinitin(\b2v_inst.valor_max_final4_3_cry_7 ),
            .carryinitout(bfn_17_9_0_));
    defparam IN_MUX_bfv_17_5_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_5_0_));
    defparam IN_MUX_bfv_17_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_6_0_ (
            .carryinitin(\b2v_inst.valor_max_final4_2_cry_7 ),
            .carryinitout(bfn_17_6_0_));
    defparam IN_MUX_bfv_18_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_6_0_));
    defparam IN_MUX_bfv_18_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_7_0_ (
            .carryinitin(\b2v_inst.un2_valor_max2_cry_7 ),
            .carryinitout(bfn_18_7_0_));
    defparam IN_MUX_bfv_13_16_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_16_0_));
    defparam IN_MUX_bfv_13_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_17_0_ (
            .carryinitin(\b2v_inst.dir_energia_cry_7 ),
            .carryinitout(bfn_13_17_0_));
    defparam IN_MUX_bfv_15_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_8_0_));
    defparam IN_MUX_bfv_15_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_9_0_ (
            .carryinitin(\b2v_inst.data_a_escribir11_7 ),
            .carryinitout(bfn_15_9_0_));
    defparam IN_MUX_bfv_17_16_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_16_0_));
    defparam IN_MUX_bfv_5_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_13_0_));
    defparam IN_MUX_bfv_5_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_14_0_ (
            .carryinitin(\b2v_inst4.un1_pix_count_int_cry_7 ),
            .carryinitout(bfn_5_14_0_));
    defparam IN_MUX_bfv_5_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_15_0_ (
            .carryinitin(\b2v_inst4.un1_pix_count_int_cry_15 ),
            .carryinitout(bfn_5_15_0_));
    defparam IN_MUX_bfv_14_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_14_0_));
    defparam IN_MUX_bfv_14_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_15_0_ (
            .carryinitin(\b2v_inst.un14_data_ram_energia_o_cry_7 ),
            .carryinitout(bfn_14_15_0_));
    defparam IN_MUX_bfv_13_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_6_0_));
    defparam IN_MUX_bfv_13_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_7_0_ (
            .carryinitin(\b2v_inst.un2_dir_mem_2_cry_7 ),
            .carryinitout(bfn_13_7_0_));
    defparam IN_MUX_bfv_8_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_5_0_));
    defparam IN_MUX_bfv_8_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_6_0_ (
            .carryinitin(\b2v_inst.un2_dir_mem_1_cry_7 ),
            .carryinitout(bfn_8_6_0_));
    defparam IN_MUX_bfv_15_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_10_0_));
    defparam IN_MUX_bfv_15_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_11_0_ (
            .carryinitin(\b2v_inst.eventos_cry_7 ),
            .carryinitout(bfn_15_11_0_));
    defparam IN_MUX_bfv_17_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_10_0_));
    defparam IN_MUX_bfv_17_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_11_0_ (
            .carryinitin(\b2v_inst.valor_max_final4_1_cry_7 ),
            .carryinitout(bfn_17_11_0_));
    defparam IN_MUX_bfv_18_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_8_0_));
    defparam IN_MUX_bfv_18_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_9_0_ (
            .carryinitin(\b2v_inst.valor_max_final4_0_cry_7 ),
            .carryinitout(bfn_18_9_0_));
    defparam IN_MUX_bfv_16_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_6_0_));
    defparam IN_MUX_bfv_16_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_7_0_ (
            .carryinitin(\b2v_inst.un2_valor_max1_cry_7 ),
            .carryinitout(bfn_16_7_0_));
    ICE_GB \b2v_inst.state_RNI9A7V8_0_29  (
            .USERSIGNALTOGLOBALBUFFER(N__14927),
            .GLOBALBUFFEROUTPUT(\b2v_inst.N_305_1_g ));
    ICE_GB reset_ibuf_RNI8255_0 (
            .USERSIGNALTOGLOBALBUFFER(N__24088),
            .GLOBALBUFFEROUTPUT(reset_c_i_g));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam reset_ibuf_RNI8255_LC_1_6_7.C_ON=1'b0;
    defparam reset_ibuf_RNI8255_LC_1_6_7.SEQ_MODE=4'b0000;
    defparam reset_ibuf_RNI8255_LC_1_6_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 reset_ibuf_RNI8255_LC_1_6_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27787),
            .lcout(reset_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un4_pix_count_intlto6_1_x1_LC_1_11_0 .C_ON=1'b0;
    defparam \b2v_inst.un4_pix_count_intlto6_1_x1_LC_1_11_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un4_pix_count_intlto6_1_x1_LC_1_11_0 .LUT_INIT=16'b0000011100001111;
    LogicCell40 \b2v_inst.un4_pix_count_intlto6_1_x1_LC_1_11_0  (
            .in0(N__16747),
            .in1(N__15018),
            .in2(N__16852),
            .in3(N__15043),
            .lcout(\b2v_inst.un4_pix_count_intlto6_1_xZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNO_27_29_LC_1_11_1 .C_ON=1'b0;
    defparam \b2v_inst.state_RNO_27_29_LC_1_11_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNO_27_29_LC_1_11_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \b2v_inst.state_RNO_27_29_LC_1_11_1  (
            .in0(N__15019),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15042),
            .lcout(),
            .ltout(\b2v_inst.N_4_i_i_a3_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNO_19_29_LC_1_11_2 .C_ON=1'b0;
    defparam \b2v_inst.state_RNO_19_29_LC_1_11_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNO_19_29_LC_1_11_2 .LUT_INIT=16'b1111110011101100;
    LogicCell40 \b2v_inst.state_RNO_19_29_LC_1_11_2  (
            .in0(N__16748),
            .in1(N__16847),
            .in2(N__13085),
            .in3(N__13148),
            .lcout(\b2v_inst.N_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un4_pix_count_intlto6_1_x0_LC_1_11_3 .C_ON=1'b0;
    defparam \b2v_inst.un4_pix_count_intlto6_1_x0_LC_1_11_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un4_pix_count_intlto6_1_x0_LC_1_11_3 .LUT_INIT=16'b0000000001110111;
    LogicCell40 \b2v_inst.un4_pix_count_intlto6_1_x0_LC_1_11_3  (
            .in0(N__15017),
            .in1(N__15041),
            .in2(_gnd_net_),
            .in3(N__16843),
            .lcout(\b2v_inst.un4_pix_count_intlto6_1_xZ0Z0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst4.pix_count_int_fast_5_LC_1_11_4 .C_ON=1'b0;
    defparam \b2v_inst4.pix_count_int_fast_5_LC_1_11_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst4.pix_count_int_fast_5_LC_1_11_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \b2v_inst4.pix_count_int_fast_5_LC_1_11_4  (
            .in0(N__14786),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13970),
            .lcout(b2v_inst4_pix_count_int_fast_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34509),
            .ce(),
            .sr(N__38041));
    defparam \b2v_inst4.pix_count_int_fast_6_LC_1_11_5 .C_ON=1'b0;
    defparam \b2v_inst4.pix_count_int_fast_6_LC_1_11_5 .SEQ_MODE=4'b1010;
    defparam \b2v_inst4.pix_count_int_fast_6_LC_1_11_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \b2v_inst4.pix_count_int_fast_6_LC_1_11_5  (
            .in0(_gnd_net_),
            .in1(N__14784),
            .in2(_gnd_net_),
            .in3(N__13952),
            .lcout(b2v_inst4_pix_count_int_fast_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34509),
            .ce(),
            .sr(N__38041));
    defparam \b2v_inst4.pix_count_int_5_LC_1_11_6 .C_ON=1'b0;
    defparam \b2v_inst4.pix_count_int_5_LC_1_11_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst4.pix_count_int_5_LC_1_11_6 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \b2v_inst4.pix_count_int_5_LC_1_11_6  (
            .in0(N__14785),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13969),
            .lcout(SYNTHESIZED_WIRE_4_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34509),
            .ce(),
            .sr(N__38041));
    defparam \b2v_inst.un7_pix_count_int_0_I_15_c_RNO_LC_1_11_7 .C_ON=1'b0;
    defparam \b2v_inst.un7_pix_count_int_0_I_15_c_RNO_LC_1_11_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un7_pix_count_int_0_I_15_c_RNO_LC_1_11_7 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \b2v_inst.un7_pix_count_int_0_I_15_c_RNO_LC_1_11_7  (
            .in0(N__13265),
            .in1(N__16746),
            .in2(N__15807),
            .in3(N__13184),
            .lcout(\b2v_inst.un7_pix_count_int_0_I_15_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.g0_3_LC_1_12_0 .C_ON=1'b0;
    defparam \b2v_inst.g0_3_LC_1_12_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.g0_3_LC_1_12_0 .LUT_INIT=16'b0101111101111111;
    LogicCell40 \b2v_inst.g0_3_LC_1_12_0  (
            .in0(N__13142),
            .in1(N__13097),
            .in2(N__13130),
            .in3(N__13163),
            .lcout(),
            .ltout(\b2v_inst.un4_pix_count_intlto6_d_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.g2_1_LC_1_12_1 .C_ON=1'b0;
    defparam \b2v_inst.g2_1_LC_1_12_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.g2_1_LC_1_12_1 .LUT_INIT=16'b0111011111110111;
    LogicCell40 \b2v_inst.g2_1_LC_1_12_1  (
            .in0(N__15878),
            .in1(N__15801),
            .in2(N__13100),
            .in3(N__16756),
            .lcout(\b2v_inst.g2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un4_pix_count_intlto6_d_1_LC_1_12_2 .C_ON=1'b0;
    defparam \b2v_inst.un4_pix_count_intlto6_d_1_LC_1_12_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un4_pix_count_intlto6_d_1_LC_1_12_2 .LUT_INIT=16'b0101111101111111;
    LogicCell40 \b2v_inst.un4_pix_count_intlto6_d_1_LC_1_12_2  (
            .in0(N__13140),
            .in1(N__13096),
            .in2(N__13129),
            .in3(N__13162),
            .lcout(\b2v_inst.un4_pix_count_intlto6_dZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst4.pix_count_int_fast_1_LC_1_12_3 .C_ON=1'b0;
    defparam \b2v_inst4.pix_count_int_fast_1_LC_1_12_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst4.pix_count_int_fast_1_LC_1_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst4.pix_count_int_fast_1_LC_1_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14036),
            .lcout(b2v_inst4_pix_count_int_fast_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34514),
            .ce(),
            .sr(N__38042));
    defparam \b2v_inst.un7_pix_count_int_0_I_1_c_RNO_LC_1_12_4 .C_ON=1'b0;
    defparam \b2v_inst.un7_pix_count_int_0_I_1_c_RNO_LC_1_12_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un7_pix_count_int_0_I_1_c_RNO_LC_1_12_4 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \b2v_inst.un7_pix_count_int_0_I_1_c_RNO_LC_1_12_4  (
            .in0(N__13161),
            .in1(N__13095),
            .in2(N__13112),
            .in3(N__13271),
            .lcout(\b2v_inst.un7_pix_count_int_0_I_1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst4.pix_count_int_fast_0_LC_1_12_5 .C_ON=1'b0;
    defparam \b2v_inst4.pix_count_int_fast_0_LC_1_12_5 .SEQ_MODE=4'b1010;
    defparam \b2v_inst4.pix_count_int_fast_0_LC_1_12_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \b2v_inst4.pix_count_int_fast_0_LC_1_12_5  (
            .in0(_gnd_net_),
            .in1(N__13808),
            .in2(_gnd_net_),
            .in3(N__14791),
            .lcout(b2v_inst4_pix_count_int_fast_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34514),
            .ce(),
            .sr(N__38042));
    defparam \b2v_inst.state_RNO_28_29_LC_1_12_7 .C_ON=1'b0;
    defparam \b2v_inst.state_RNO_28_29_LC_1_12_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNO_28_29_LC_1_12_7 .LUT_INIT=16'b1100100000000000;
    LogicCell40 \b2v_inst.state_RNO_28_29_LC_1_12_7  (
            .in0(N__15273),
            .in1(N__13141),
            .in2(N__15199),
            .in3(N__13125),
            .lcout(\b2v_inst.N_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst4.pix_count_int_fast_2_LC_1_13_0 .C_ON=1'b0;
    defparam \b2v_inst4.pix_count_int_fast_2_LC_1_13_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst4.pix_count_int_fast_2_LC_1_13_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \b2v_inst4.pix_count_int_fast_2_LC_1_13_0  (
            .in0(N__14778),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14012),
            .lcout(b2v_inst4_pix_count_int_fast_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34523),
            .ce(),
            .sr(N__38043));
    defparam \b2v_inst4.pix_count_int_0_LC_1_13_3 .C_ON=1'b0;
    defparam \b2v_inst4.pix_count_int_0_LC_1_13_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst4.pix_count_int_0_LC_1_13_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \b2v_inst4.pix_count_int_0_LC_1_13_3  (
            .in0(_gnd_net_),
            .in1(N__13801),
            .in2(_gnd_net_),
            .in3(N__14783),
            .lcout(SYNTHESIZED_WIRE_4_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34523),
            .ce(),
            .sr(N__38043));
    defparam \b2v_inst4.pix_count_int_fast_3_LC_1_13_4 .C_ON=1'b0;
    defparam \b2v_inst4.pix_count_int_fast_3_LC_1_13_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst4.pix_count_int_fast_3_LC_1_13_4 .LUT_INIT=16'b0000101000001010;
    LogicCell40 \b2v_inst4.pix_count_int_fast_3_LC_1_13_4  (
            .in0(N__13988),
            .in1(_gnd_net_),
            .in2(N__14792),
            .in3(_gnd_net_),
            .lcout(b2v_inst4_pix_count_int_fast_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34523),
            .ce(),
            .sr(N__38043));
    defparam \b2v_inst4.pix_count_int_3_LC_1_13_5 .C_ON=1'b0;
    defparam \b2v_inst4.pix_count_int_3_LC_1_13_5 .SEQ_MODE=4'b1010;
    defparam \b2v_inst4.pix_count_int_3_LC_1_13_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \b2v_inst4.pix_count_int_3_LC_1_13_5  (
            .in0(_gnd_net_),
            .in1(N__14779),
            .in2(_gnd_net_),
            .in3(N__13987),
            .lcout(SYNTHESIZED_WIRE_4_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34523),
            .ce(),
            .sr(N__38043));
    defparam \b2v_inst4.pix_count_int_fast_11_LC_1_13_6 .C_ON=1'b0;
    defparam \b2v_inst4.pix_count_int_fast_11_LC_1_13_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst4.pix_count_int_fast_11_LC_1_13_6 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \b2v_inst4.pix_count_int_fast_11_LC_1_13_6  (
            .in0(N__14777),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14687),
            .lcout(b2v_inst4_pix_count_int_fast_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34523),
            .ce(),
            .sr(N__38043));
    defparam \b2v_inst4.state_RNI8N511_0_LC_1_14_1 .C_ON=1'b0;
    defparam \b2v_inst4.state_RNI8N511_0_LC_1_14_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst4.state_RNI8N511_0_LC_1_14_1 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \b2v_inst4.state_RNI8N511_0_LC_1_14_1  (
            .in0(N__14897),
            .in1(N__15503),
            .in2(_gnd_net_),
            .in3(N__15875),
            .lcout(\b2v_inst4.un1_pix_count_int_0_sqmuxa_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.pix_count_anterior_1_LC_2_10_0 .C_ON=1'b0;
    defparam \b2v_inst.pix_count_anterior_1_LC_2_10_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.pix_count_anterior_1_LC_2_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.pix_count_anterior_1_LC_2_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15193),
            .lcout(\b2v_inst.pix_count_anteriorZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34511),
            .ce(N__13845),
            .sr(N__38040));
    defparam \b2v_inst.pix_count_anterior_4_LC_2_10_1 .C_ON=1'b0;
    defparam \b2v_inst.pix_count_anterior_4_LC_2_10_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.pix_count_anterior_4_LC_2_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.pix_count_anterior_4_LC_2_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16757),
            .lcout(\b2v_inst.pix_count_anteriorZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34511),
            .ce(N__13845),
            .sr(N__38040));
    defparam \b2v_inst.pix_count_anterior_9_LC_2_10_2 .C_ON=1'b0;
    defparam \b2v_inst.pix_count_anterior_9_LC_2_10_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.pix_count_anterior_9_LC_2_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.pix_count_anterior_9_LC_2_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15566),
            .lcout(\b2v_inst.pix_count_anteriorZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34511),
            .ce(N__13845),
            .sr(N__38040));
    defparam \b2v_inst.cuenta_pixel_7_LC_2_10_3 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_pixel_7_LC_2_10_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.cuenta_pixel_7_LC_2_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.cuenta_pixel_7_LC_2_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13445),
            .lcout(\b2v_inst.cuenta_pixelZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34511),
            .ce(N__13845),
            .sr(N__38040));
    defparam \b2v_inst.cuenta_pixel_8_LC_2_10_5 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_pixel_8_LC_2_10_5 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.cuenta_pixel_8_LC_2_10_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \b2v_inst.cuenta_pixel_8_LC_2_10_5  (
            .in0(N__13397),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14583),
            .lcout(\b2v_inst.cuenta_pixelZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34511),
            .ce(N__13845),
            .sr(N__38040));
    defparam \b2v_inst.un7_pix_count_int_0_I_1_c_LC_2_11_0 .C_ON=1'b1;
    defparam \b2v_inst.un7_pix_count_int_0_I_1_c_LC_2_11_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un7_pix_count_int_0_I_1_c_LC_2_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.un7_pix_count_int_0_I_1_c_LC_2_11_0  (
            .in0(_gnd_net_),
            .in1(N__13178),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_11_0_),
            .carryout(\b2v_inst.un7_pix_count_int_0_data_tmp_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un7_pix_count_int_0_I_27_c_LC_2_11_1 .C_ON=1'b1;
    defparam \b2v_inst.un7_pix_count_int_0_I_27_c_LC_2_11_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un7_pix_count_int_0_I_27_c_LC_2_11_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.un7_pix_count_int_0_I_27_c_LC_2_11_1  (
            .in0(_gnd_net_),
            .in1(N__37300),
            .in2(N__13196),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.un7_pix_count_int_0_data_tmp_0 ),
            .carryout(\b2v_inst.un7_pix_count_int_0_data_tmp_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un7_pix_count_int_0_I_15_c_LC_2_11_2 .C_ON=1'b1;
    defparam \b2v_inst.un7_pix_count_int_0_I_15_c_LC_2_11_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un7_pix_count_int_0_I_15_c_LC_2_11_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.un7_pix_count_int_0_I_15_c_LC_2_11_2  (
            .in0(_gnd_net_),
            .in1(N__37296),
            .in2(N__13172),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.un7_pix_count_int_0_data_tmp_1 ),
            .carryout(\b2v_inst.un7_pix_count_int_0_data_tmp_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un7_pix_count_int_0_I_21_c_LC_2_11_3 .C_ON=1'b1;
    defparam \b2v_inst.un7_pix_count_int_0_I_21_c_LC_2_11_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un7_pix_count_int_0_I_21_c_LC_2_11_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.un7_pix_count_int_0_I_21_c_LC_2_11_3  (
            .in0(_gnd_net_),
            .in1(N__37299),
            .in2(N__13517),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.un7_pix_count_int_0_data_tmp_2 ),
            .carryout(\b2v_inst.un7_pix_count_int_0_data_tmp_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un7_pix_count_int_0_I_51_c_LC_2_11_4 .C_ON=1'b1;
    defparam \b2v_inst.un7_pix_count_int_0_I_51_c_LC_2_11_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un7_pix_count_int_0_I_51_c_LC_2_11_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.un7_pix_count_int_0_I_51_c_LC_2_11_4  (
            .in0(_gnd_net_),
            .in1(N__37298),
            .in2(N__13544),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.un7_pix_count_int_0_data_tmp_3 ),
            .carryout(\b2v_inst.un7_pix_count_int_0_data_tmp_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un7_pix_count_int_0_I_9_c_LC_2_11_5 .C_ON=1'b1;
    defparam \b2v_inst.un7_pix_count_int_0_I_9_c_LC_2_11_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un7_pix_count_int_0_I_9_c_LC_2_11_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.un7_pix_count_int_0_I_9_c_LC_2_11_5  (
            .in0(_gnd_net_),
            .in1(N__37302),
            .in2(N__13889),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.un7_pix_count_int_0_data_tmp_4 ),
            .carryout(\b2v_inst.un7_pix_count_int_0_data_tmp_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un7_pix_count_int_0_I_39_c_LC_2_11_6 .C_ON=1'b1;
    defparam \b2v_inst.un7_pix_count_int_0_I_39_c_LC_2_11_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un7_pix_count_int_0_I_39_c_LC_2_11_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.un7_pix_count_int_0_I_39_c_LC_2_11_6  (
            .in0(_gnd_net_),
            .in1(N__37297),
            .in2(N__13241),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.un7_pix_count_int_0_data_tmp_5 ),
            .carryout(\b2v_inst.un7_pix_count_int_0_data_tmp_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un7_pix_count_int_0_I_45_c_LC_2_11_7 .C_ON=1'b1;
    defparam \b2v_inst.un7_pix_count_int_0_I_45_c_LC_2_11_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un7_pix_count_int_0_I_45_c_LC_2_11_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.un7_pix_count_int_0_I_45_c_LC_2_11_7  (
            .in0(_gnd_net_),
            .in1(N__37301),
            .in2(N__13343),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.un7_pix_count_int_0_data_tmp_6 ),
            .carryout(\b2v_inst.un7_pix_count_int_0_data_tmp_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un7_pix_count_int_0_I_57_c_LC_2_12_0 .C_ON=1'b1;
    defparam \b2v_inst.un7_pix_count_int_0_I_57_c_LC_2_12_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un7_pix_count_int_0_I_57_c_LC_2_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.un7_pix_count_int_0_I_57_c_LC_2_12_0  (
            .in0(_gnd_net_),
            .in1(N__37265),
            .in2(N__13217),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_12_0_),
            .carryout(\b2v_inst.un7_pix_count_int_0_data_tmp_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un7_pix_count_int_0_I_33_c_LC_2_12_1 .C_ON=1'b1;
    defparam \b2v_inst.un7_pix_count_int_0_I_33_c_LC_2_12_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un7_pix_count_int_0_I_33_c_LC_2_12_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.un7_pix_count_int_0_I_33_c_LC_2_12_1  (
            .in0(_gnd_net_),
            .in1(N__37264),
            .in2(N__13256),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.un7_pix_count_int_0_data_tmp_8 ),
            .carryout(\b2v_inst.un7_pix_count_int_0_N_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un7_pix_count_int_0_N_2_THRU_LUT4_0_LC_2_12_2 .C_ON=1'b0;
    defparam \b2v_inst.un7_pix_count_int_0_N_2_THRU_LUT4_0_LC_2_12_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un7_pix_count_int_0_N_2_THRU_LUT4_0_LC_2_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.un7_pix_count_int_0_N_2_THRU_LUT4_0_LC_2_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13220),
            .lcout(\b2v_inst.un7_pix_count_int_0_N_2_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un7_pix_count_int_0_I_57_c_RNO_LC_2_12_3 .C_ON=1'b0;
    defparam \b2v_inst.un7_pix_count_int_0_I_57_c_RNO_LC_2_12_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un7_pix_count_int_0_I_57_c_RNO_LC_2_12_3 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \b2v_inst.un7_pix_count_int_0_I_57_c_RNO_LC_2_12_3  (
            .in0(N__17610),
            .in1(N__17445),
            .in2(N__13301),
            .in3(N__13862),
            .lcout(\b2v_inst.un7_pix_count_int_0_I_57_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.g0_5_LC_2_12_5 .C_ON=1'b0;
    defparam \b2v_inst.g0_5_LC_2_12_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.g0_5_LC_2_12_5 .LUT_INIT=16'b0011011111111111;
    LogicCell40 \b2v_inst.g0_5_LC_2_12_5  (
            .in0(N__15262),
            .in1(N__15226),
            .in2(N__15198),
            .in3(N__15132),
            .lcout(\b2v_inst.un4_pix_count_intlto6_d_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst4.state_RNI9BF02_0_LC_2_12_7 .C_ON=1'b0;
    defparam \b2v_inst4.state_RNI9BF02_0_LC_2_12_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst4.state_RNI9BF02_0_LC_2_12_7 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \b2v_inst4.state_RNI9BF02_0_LC_2_12_7  (
            .in0(N__13208),
            .in1(N__14876),
            .in2(_gnd_net_),
            .in3(N__15641),
            .lcout(\b2v_inst4.un1_pix_count_int_0_sqmuxa_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un7_pix_count_int_0_I_27_c_RNO_LC_2_13_0 .C_ON=1'b0;
    defparam \b2v_inst.un7_pix_count_int_0_I_27_c_RNO_LC_2_13_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un7_pix_count_int_0_I_27_c_RNO_LC_2_13_0 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \b2v_inst.un7_pix_count_int_0_I_27_c_RNO_LC_2_13_0  (
            .in0(N__15225),
            .in1(N__13286),
            .in2(N__13280),
            .in3(N__15121),
            .lcout(\b2v_inst.un7_pix_count_int_0_I_27_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.pix_count_anterior_2_LC_2_13_1 .C_ON=1'b0;
    defparam \b2v_inst.pix_count_anterior_2_LC_2_13_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.pix_count_anterior_2_LC_2_13_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst.pix_count_anterior_2_LC_2_13_1  (
            .in0(N__15123),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst.pix_count_anteriorZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34515),
            .ce(N__13846),
            .sr(N__38046));
    defparam \b2v_inst.pix_count_anterior_3_LC_2_13_2 .C_ON=1'b0;
    defparam \b2v_inst.pix_count_anterior_3_LC_2_13_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.pix_count_anterior_3_LC_2_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.pix_count_anterior_3_LC_2_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15236),
            .lcout(\b2v_inst.pix_count_anteriorZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34515),
            .ce(N__13846),
            .sr(N__38046));
    defparam \b2v_inst4.pix_count_int_RNIQK3K1_0_LC_2_13_3 .C_ON=1'b0;
    defparam \b2v_inst4.pix_count_int_RNIQK3K1_0_LC_2_13_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst4.pix_count_int_RNIQK3K1_0_LC_2_13_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst4.pix_count_int_RNIQK3K1_0_LC_2_13_3  (
            .in0(N__15122),
            .in1(N__15271),
            .in2(N__15239),
            .in3(N__15824),
            .lcout(\b2v_inst4.un1_pix_count_int_0_sqmuxa_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.pix_count_anterior_0_LC_2_13_4 .C_ON=1'b0;
    defparam \b2v_inst.pix_count_anterior_0_LC_2_13_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.pix_count_anterior_0_LC_2_13_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst.pix_count_anterior_0_LC_2_13_4  (
            .in0(N__15272),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst.pix_count_anteriorZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34515),
            .ce(N__13846),
            .sr(N__38046));
    defparam \b2v_inst.pix_count_anterior_5_LC_2_13_5 .C_ON=1'b0;
    defparam \b2v_inst.pix_count_anterior_5_LC_2_13_5 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.pix_count_anterior_5_LC_2_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.pix_count_anterior_5_LC_2_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15825),
            .lcout(\b2v_inst.pix_count_anteriorZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34515),
            .ce(N__13846),
            .sr(N__38046));
    defparam \b2v_inst.un7_pix_count_int_0_I_33_c_RNO_LC_2_13_6 .C_ON=1'b0;
    defparam \b2v_inst.un7_pix_count_int_0_I_33_c_RNO_LC_2_13_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un7_pix_count_int_0_I_33_c_RNO_LC_2_13_6 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \b2v_inst.un7_pix_count_int_0_I_33_c_RNO_LC_2_13_6  (
            .in0(N__17500),
            .in1(N__17722),
            .in2(N__13313),
            .in3(N__13247),
            .lcout(\b2v_inst.un7_pix_count_int_0_I_33_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.pix_count_anterior_18_LC_2_13_7 .C_ON=1'b0;
    defparam \b2v_inst.pix_count_anterior_18_LC_2_13_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.pix_count_anterior_18_LC_2_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.pix_count_anterior_18_LC_2_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17501),
            .lcout(\b2v_inst.pix_count_anteriorZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34515),
            .ce(N__13846),
            .sr(N__38046));
    defparam \b2v_inst.un7_pix_count_int_0_I_39_c_RNO_LC_2_14_0 .C_ON=1'b0;
    defparam \b2v_inst.un7_pix_count_int_0_I_39_c_RNO_LC_2_14_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un7_pix_count_int_0_I_39_c_RNO_LC_2_14_0 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \b2v_inst.un7_pix_count_int_0_I_39_c_RNO_LC_2_14_0  (
            .in0(N__15376),
            .in1(N__16474),
            .in2(N__13229),
            .in3(N__13349),
            .lcout(\b2v_inst.un7_pix_count_int_0_I_39_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.pix_count_anterior_12_LC_2_14_1 .C_ON=1'b0;
    defparam \b2v_inst.pix_count_anterior_12_LC_2_14_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.pix_count_anterior_12_LC_2_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.pix_count_anterior_12_LC_2_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15377),
            .lcout(\b2v_inst.pix_count_anteriorZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34524),
            .ce(N__13848),
            .sr(N__38049));
    defparam \b2v_inst.pix_count_anterior_13_LC_2_14_2 .C_ON=1'b0;
    defparam \b2v_inst.pix_count_anterior_13_LC_2_14_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.pix_count_anterior_13_LC_2_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.pix_count_anterior_13_LC_2_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16475),
            .lcout(\b2v_inst.pix_count_anteriorZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34524),
            .ce(N__13848),
            .sr(N__38049));
    defparam \b2v_inst.un7_pix_count_int_0_I_45_c_RNO_LC_2_14_3 .C_ON=1'b0;
    defparam \b2v_inst.un7_pix_count_int_0_I_45_c_RNO_LC_2_14_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un7_pix_count_int_0_I_45_c_RNO_LC_2_14_3 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \b2v_inst.un7_pix_count_int_0_I_45_c_RNO_LC_2_14_3  (
            .in0(N__16408),
            .in1(N__16338),
            .in2(N__13331),
            .in3(N__13319),
            .lcout(\b2v_inst.un7_pix_count_int_0_I_45_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.pix_count_anterior_14_LC_2_14_4 .C_ON=1'b0;
    defparam \b2v_inst.pix_count_anterior_14_LC_2_14_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.pix_count_anterior_14_LC_2_14_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst.pix_count_anterior_14_LC_2_14_4  (
            .in0(N__16340),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst.pix_count_anteriorZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34524),
            .ce(N__13848),
            .sr(N__38049));
    defparam \b2v_inst4.pix_count_int_RNIDQ1Q_1_LC_2_14_5 .C_ON=1'b0;
    defparam \b2v_inst4.pix_count_int_RNIDQ1Q_1_LC_2_14_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst4.pix_count_int_RNIDQ1Q_1_LC_2_14_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \b2v_inst4.pix_count_int_RNIDQ1Q_1_LC_2_14_5  (
            .in0(_gnd_net_),
            .in1(N__15171),
            .in2(_gnd_net_),
            .in3(N__16752),
            .lcout(),
            .ltout(\b2v_inst4.un1_pix_count_int_0_sqmuxa_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst4.pix_count_int_RNII16D3_14_LC_2_14_6 .C_ON=1'b0;
    defparam \b2v_inst4.pix_count_int_RNII16D3_14_LC_2_14_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst4.pix_count_int_RNII16D3_14_LC_2_14_6 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \b2v_inst4.pix_count_int_RNII16D3_14_LC_2_14_6  (
            .in0(N__16339),
            .in1(N__16409),
            .in2(N__13322),
            .in3(N__13787),
            .lcout(\b2v_inst4.un1_pix_count_int_0_sqmuxa_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.pix_count_anterior_15_LC_2_14_7 .C_ON=1'b0;
    defparam \b2v_inst.pix_count_anterior_15_LC_2_14_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.pix_count_anterior_15_LC_2_14_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst.pix_count_anterior_15_LC_2_14_7  (
            .in0(N__16410),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst.pix_count_anteriorZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34524),
            .ce(N__13848),
            .sr(N__38049));
    defparam \b2v_inst.pix_count_anterior_19_LC_2_15_3 .C_ON=1'b0;
    defparam \b2v_inst.pix_count_anterior_19_LC_2_15_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.pix_count_anterior_19_LC_2_15_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.pix_count_anterior_19_LC_2_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17705),
            .lcout(\b2v_inst.pix_count_anteriorZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34525),
            .ce(N__13850),
            .sr(N__38053));
    defparam \b2v_inst.pix_count_anterior_16_LC_2_15_7 .C_ON=1'b0;
    defparam \b2v_inst.pix_count_anterior_16_LC_2_15_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.pix_count_anterior_16_LC_2_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.pix_count_anterior_16_LC_2_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17612),
            .lcout(\b2v_inst.pix_count_anteriorZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34525),
            .ce(N__13850),
            .sr(N__38053));
    defparam \b2v_inst.cuenta_pixel_9_LC_3_8_0 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_pixel_9_LC_3_8_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.cuenta_pixel_9_LC_3_8_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \b2v_inst.cuenta_pixel_9_LC_3_8_0  (
            .in0(N__13393),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14641),
            .lcout(\b2v_inst.cuenta_pixelZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34516),
            .ce(N__13851),
            .sr(N__38047));
    defparam \b2v_inst.cuenta_pixel_0_LC_3_8_1 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_pixel_0_LC_3_8_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.cuenta_pixel_0_LC_3_8_1 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \b2v_inst.cuenta_pixel_0_LC_3_8_1  (
            .in0(_gnd_net_),
            .in1(N__13392),
            .in2(_gnd_net_),
            .in3(N__13747),
            .lcout(\b2v_inst.cuenta_pixelZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34516),
            .ce(N__13851),
            .sr(N__38047));
    defparam \b2v_inst.cuenta_pixel_RNINOUV1_10_LC_3_8_3 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_pixel_RNINOUV1_10_LC_3_8_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.cuenta_pixel_RNINOUV1_10_LC_3_8_3 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \b2v_inst.cuenta_pixel_RNINOUV1_10_LC_3_8_3  (
            .in0(N__14640),
            .in1(N__14617),
            .in2(N__14590),
            .in3(N__13658),
            .lcout(),
            .ltout(\b2v_inst.un1_state_36_0_a2_0_2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.cuenta_pixel_RNIISKR5_0_LC_3_8_4 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_pixel_RNIISKR5_0_LC_3_8_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.cuenta_pixel_RNIISKR5_0_LC_3_8_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst.cuenta_pixel_RNIISKR5_0_LC_3_8_4  (
            .in0(N__13634),
            .in1(N__13616),
            .in2(N__13400),
            .in3(N__14557),
            .lcout(\b2v_inst.N_305_2 ),
            .ltout(\b2v_inst.N_305_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.cuenta_pixel_6_LC_3_8_5 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_pixel_6_LC_3_8_5 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.cuenta_pixel_6_LC_3_8_5 .LUT_INIT=16'b0000110000001100;
    LogicCell40 \b2v_inst.cuenta_pixel_6_LC_3_8_5  (
            .in0(_gnd_net_),
            .in1(N__13469),
            .in2(N__13379),
            .in3(_gnd_net_),
            .lcout(\b2v_inst.cuenta_pixelZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34516),
            .ce(N__13851),
            .sr(N__38047));
    defparam \b2v_inst.cuenta_pixel_1_LC_3_8_6 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_pixel_1_LC_3_8_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.cuenta_pixel_1_LC_3_8_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst.cuenta_pixel_1_LC_3_8_6  (
            .in0(N__13748),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13375),
            .lcout(\b2v_inst.cuenta_pixelZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34516),
            .ce(N__13851),
            .sr(N__38047));
    defparam \b2v_inst.cuenta_pixel_RNIT0FM_1_LC_3_9_1 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_pixel_RNIT0FM_1_LC_3_9_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.cuenta_pixel_RNIT0FM_1_LC_3_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst.cuenta_pixel_RNIT0FM_1_LC_3_9_1  (
            .in0(_gnd_net_),
            .in1(N__13743),
            .in2(_gnd_net_),
            .in3(N__13374),
            .lcout(\b2v_inst.cuenta_pixel_RNIT0FMZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un1_cuenta_pixel_cry_5_c_RNI2E441_LC_3_9_5 .C_ON=1'b0;
    defparam \b2v_inst.un1_cuenta_pixel_cry_5_c_RNI2E441_LC_3_9_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un1_cuenta_pixel_cry_5_c_RNI2E441_LC_3_9_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \b2v_inst.un1_cuenta_pixel_cry_5_c_RNI2E441_LC_3_9_5  (
            .in0(N__13444),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13465),
            .lcout(\b2v_inst.cuenta_pixel_5_i_a2_1_1_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un1_cuenta_pixel_cry_1_c_LC_3_10_0 .C_ON=1'b1;
    defparam \b2v_inst.un1_cuenta_pixel_cry_1_c_LC_3_10_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un1_cuenta_pixel_cry_1_c_LC_3_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.un1_cuenta_pixel_cry_1_c_LC_3_10_0  (
            .in0(_gnd_net_),
            .in1(N__13376),
            .in2(N__13758),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_3_10_0_),
            .carryout(\b2v_inst.un1_cuenta_pixel_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un1_cuenta_pixel_cry_1_c_RNI89TH_LC_3_10_1 .C_ON=1'b1;
    defparam \b2v_inst.un1_cuenta_pixel_cry_1_c_RNI89TH_LC_3_10_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un1_cuenta_pixel_cry_1_c_RNI89TH_LC_3_10_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.un1_cuenta_pixel_cry_1_c_RNI89TH_LC_3_10_1  (
            .in0(_gnd_net_),
            .in1(N__13709),
            .in2(_gnd_net_),
            .in3(N__13355),
            .lcout(\b2v_inst.un1_cuenta_pixel_cry_1_c_RNI89THZ0 ),
            .ltout(),
            .carryin(\b2v_inst.un1_cuenta_pixel_cry_1 ),
            .carryout(\b2v_inst.un1_cuenta_pixel_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un1_cuenta_pixel_cry_2_c_RNIACUH_LC_3_10_2 .C_ON=1'b1;
    defparam \b2v_inst.un1_cuenta_pixel_cry_2_c_RNIACUH_LC_3_10_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un1_cuenta_pixel_cry_2_c_RNIACUH_LC_3_10_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.un1_cuenta_pixel_cry_2_c_RNIACUH_LC_3_10_2  (
            .in0(_gnd_net_),
            .in1(N__13700),
            .in2(_gnd_net_),
            .in3(N__13352),
            .lcout(\b2v_inst.un1_cuenta_pixel_cry_2_c_RNIACUHZ0 ),
            .ltout(),
            .carryin(\b2v_inst.un1_cuenta_pixel_cry_2 ),
            .carryout(\b2v_inst.un1_cuenta_pixel_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un1_cuenta_pixel_cry_3_c_RNICFVH_LC_3_10_3 .C_ON=1'b1;
    defparam \b2v_inst.un1_cuenta_pixel_cry_3_c_RNICFVH_LC_3_10_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un1_cuenta_pixel_cry_3_c_RNICFVH_LC_3_10_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst.un1_cuenta_pixel_cry_3_c_RNICFVH_LC_3_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13901),
            .in3(N__13484),
            .lcout(\b2v_inst.un1_cuenta_pixel_cry_3_c_RNICFVHZ0 ),
            .ltout(),
            .carryin(\b2v_inst.un1_cuenta_pixel_cry_3 ),
            .carryout(\b2v_inst.un1_cuenta_pixel_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un1_cuenta_pixel_cry_4_c_RNIEI0I_LC_3_10_4 .C_ON=1'b1;
    defparam \b2v_inst.un1_cuenta_pixel_cry_4_c_RNIEI0I_LC_3_10_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un1_cuenta_pixel_cry_4_c_RNIEI0I_LC_3_10_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst.un1_cuenta_pixel_cry_4_c_RNIEI0I_LC_3_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13592),
            .in3(N__13481),
            .lcout(\b2v_inst.un1_cuenta_pixel_cry_4_c_RNIEI0IZ0 ),
            .ltout(),
            .carryin(\b2v_inst.un1_cuenta_pixel_cry_4 ),
            .carryout(\b2v_inst.un1_cuenta_pixel_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un1_cuenta_pixel_cry_5_c_RNIGL1I_LC_3_10_5 .C_ON=1'b1;
    defparam \b2v_inst.un1_cuenta_pixel_cry_5_c_RNIGL1I_LC_3_10_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un1_cuenta_pixel_cry_5_c_RNIGL1I_LC_3_10_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.un1_cuenta_pixel_cry_5_c_RNIGL1I_LC_3_10_5  (
            .in0(_gnd_net_),
            .in1(N__13478),
            .in2(_gnd_net_),
            .in3(N__13454),
            .lcout(\b2v_inst.un1_cuenta_pixel_cry_5_c_RNIGL1IZ0 ),
            .ltout(),
            .carryin(\b2v_inst.un1_cuenta_pixel_cry_5 ),
            .carryout(\b2v_inst.un1_cuenta_pixel_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un1_cuenta_pixel_cry_6_c_RNIIO2I_LC_3_10_6 .C_ON=1'b1;
    defparam \b2v_inst.un1_cuenta_pixel_cry_6_c_RNIIO2I_LC_3_10_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un1_cuenta_pixel_cry_6_c_RNIIO2I_LC_3_10_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.un1_cuenta_pixel_cry_6_c_RNIIO2I_LC_3_10_6  (
            .in0(_gnd_net_),
            .in1(N__13451),
            .in2(_gnd_net_),
            .in3(N__13433),
            .lcout(\b2v_inst.un1_cuenta_pixel_cry_6_c_RNIIO2IZ0 ),
            .ltout(),
            .carryin(\b2v_inst.un1_cuenta_pixel_cry_6 ),
            .carryout(\b2v_inst.un1_cuenta_pixel_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un1_cuenta_pixel_cry_7_c_RNIKR3I_LC_3_10_7 .C_ON=1'b1;
    defparam \b2v_inst.un1_cuenta_pixel_cry_7_c_RNIKR3I_LC_3_10_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un1_cuenta_pixel_cry_7_c_RNIKR3I_LC_3_10_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.un1_cuenta_pixel_cry_7_c_RNIKR3I_LC_3_10_7  (
            .in0(_gnd_net_),
            .in1(N__13430),
            .in2(_gnd_net_),
            .in3(N__13424),
            .lcout(\b2v_inst.un1_cuenta_pixel_cry_7_c_RNIKR3IZ0 ),
            .ltout(),
            .carryin(\b2v_inst.un1_cuenta_pixel_cry_7 ),
            .carryout(\b2v_inst.un1_cuenta_pixel_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un1_cuenta_pixel_cry_8_c_RNIMU4I_LC_3_11_0 .C_ON=1'b1;
    defparam \b2v_inst.un1_cuenta_pixel_cry_8_c_RNIMU4I_LC_3_11_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un1_cuenta_pixel_cry_8_c_RNIMU4I_LC_3_11_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.un1_cuenta_pixel_cry_8_c_RNIMU4I_LC_3_11_0  (
            .in0(_gnd_net_),
            .in1(N__13421),
            .in2(_gnd_net_),
            .in3(N__13412),
            .lcout(\b2v_inst.un1_cuenta_pixel_cry_8_c_RNIMU4IZ0 ),
            .ltout(),
            .carryin(bfn_3_11_0_),
            .carryout(\b2v_inst.un1_cuenta_pixel_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.cuenta_pixel_RNIVBL9_10_LC_3_11_1 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_pixel_RNIVBL9_10_LC_3_11_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.cuenta_pixel_RNIVBL9_10_LC_3_11_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \b2v_inst.cuenta_pixel_RNIVBL9_10_LC_3_11_1  (
            .in0(_gnd_net_),
            .in1(N__13406),
            .in2(_gnd_net_),
            .in3(N__13409),
            .lcout(\b2v_inst.cuenta_pixel_RNIVBL9Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.cuenta_pixel_10_LC_3_11_2 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_pixel_10_LC_3_11_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.cuenta_pixel_10_LC_3_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.cuenta_pixel_10_LC_3_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14616),
            .lcout(\b2v_inst.cuenta_pixelZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34497),
            .ce(N__13844),
            .sr(N__38044));
    defparam \b2v_inst4.pix_count_int_9_rep1_LC_3_12_3 .C_ON=1'b0;
    defparam \b2v_inst4.pix_count_int_9_rep1_LC_3_12_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst4.pix_count_int_9_rep1_LC_3_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst4.pix_count_int_9_rep1_LC_3_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14816),
            .lcout(SYNTHESIZED_WIRE_4_9_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34503),
            .ce(),
            .sr(N__38048));
    defparam \b2v_inst.un7_pix_count_int_0_I_51_c_RNO_LC_3_12_4 .C_ON=1'b0;
    defparam \b2v_inst.un7_pix_count_int_0_I_51_c_RNO_LC_3_12_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un7_pix_count_int_0_I_51_c_RNO_LC_3_12_4 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \b2v_inst.un7_pix_count_int_0_I_51_c_RNO_LC_3_12_4  (
            .in0(N__13556),
            .in1(N__15495),
            .in2(N__13493),
            .in3(N__15305),
            .lcout(\b2v_inst.un7_pix_count_int_0_I_51_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNO_26_29_LC_3_12_5 .C_ON=1'b0;
    defparam \b2v_inst.state_RNO_26_29_LC_3_12_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNO_26_29_LC_3_12_5 .LUT_INIT=16'b1100100000000000;
    LogicCell40 \b2v_inst.state_RNO_26_29_LC_3_12_5  (
            .in0(N__15306),
            .in1(N__15725),
            .in2(N__15779),
            .in3(N__15674),
            .lcout(),
            .ltout(\b2v_inst.N_1_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNO_18_29_LC_3_12_6 .C_ON=1'b0;
    defparam \b2v_inst.state_RNO_18_29_LC_3_12_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNO_18_29_LC_3_12_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \b2v_inst.state_RNO_18_29_LC_3_12_6  (
            .in0(N__16429),
            .in1(N__16362),
            .in2(N__13535),
            .in3(N__16499),
            .lcout(),
            .ltout(\b2v_inst.N_4_i_i_o6_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNO_7_29_LC_3_12_7 .C_ON=1'b0;
    defparam \b2v_inst.state_RNO_7_29_LC_3_12_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNO_7_29_LC_3_12_7 .LUT_INIT=16'b1010001010100000;
    LogicCell40 \b2v_inst.state_RNO_7_29_LC_3_12_7  (
            .in0(N__13817),
            .in1(N__16271),
            .in2(N__13532),
            .in3(N__13529),
            .lcout(\b2v_inst.N_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un7_pix_count_int_0_I_21_c_RNO_LC_3_13_0 .C_ON=1'b0;
    defparam \b2v_inst.un7_pix_count_int_0_I_21_c_RNO_LC_3_13_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un7_pix_count_int_0_I_21_c_RNO_LC_3_13_0 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \b2v_inst.un7_pix_count_int_0_I_21_c_RNO_LC_3_13_0  (
            .in0(N__13505),
            .in1(N__16822),
            .in2(N__15859),
            .in3(N__13499),
            .lcout(\b2v_inst.un7_pix_count_int_0_I_21_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.pix_count_anterior_6_LC_3_13_1 .C_ON=1'b0;
    defparam \b2v_inst.pix_count_anterior_6_LC_3_13_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.pix_count_anterior_6_LC_3_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.pix_count_anterior_6_LC_3_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15848),
            .lcout(\b2v_inst.pix_count_anteriorZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34512),
            .ce(N__13849),
            .sr(N__38050));
    defparam \b2v_inst.pix_count_anterior_7_LC_3_13_2 .C_ON=1'b0;
    defparam \b2v_inst.pix_count_anterior_7_LC_3_13_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.pix_count_anterior_7_LC_3_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.pix_count_anterior_7_LC_3_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16824),
            .lcout(\b2v_inst.pix_count_anteriorZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34512),
            .ce(N__13849),
            .sr(N__38050));
    defparam \b2v_inst.pix_count_anterior_8_LC_3_13_4 .C_ON=1'b0;
    defparam \b2v_inst.pix_count_anterior_8_LC_3_13_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.pix_count_anterior_8_LC_3_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.pix_count_anterior_8_LC_3_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15502),
            .lcout(\b2v_inst.pix_count_anteriorZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34512),
            .ce(N__13849),
            .sr(N__38050));
    defparam \b2v_inst4.pix_count_int_RNI5JOL1_9_LC_3_13_5 .C_ON=1'b0;
    defparam \b2v_inst4.pix_count_int_RNI5JOL1_9_LC_3_13_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst4.pix_count_int_RNI5JOL1_9_LC_3_13_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst4.pix_count_int_RNI5JOL1_9_LC_3_13_5  (
            .in0(N__16823),
            .in1(N__16500),
            .in2(N__15565),
            .in3(N__15617),
            .lcout(),
            .ltout(\b2v_inst4.un1_pix_count_int_0_sqmuxa_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst4.pix_count_int_RNIQKHN8_0_LC_3_13_6 .C_ON=1'b0;
    defparam \b2v_inst4.pix_count_int_RNIQKHN8_0_LC_3_13_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst4.pix_count_int_RNIQKHN8_0_LC_3_13_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst4.pix_count_int_RNIQKHN8_0_LC_3_13_6  (
            .in0(N__13580),
            .in1(N__13571),
            .in2(N__13565),
            .in3(N__13562),
            .lcout(\b2v_inst4.un1_pix_count_int_0_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst4.pix_count_int_12_LC_3_14_0 .C_ON=1'b0;
    defparam \b2v_inst4.pix_count_int_12_LC_3_14_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst4.pix_count_int_12_LC_3_14_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \b2v_inst4.pix_count_int_12_LC_3_14_0  (
            .in0(N__14752),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14068),
            .lcout(SYNTHESIZED_WIRE_4_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34517),
            .ce(),
            .sr(N__38054));
    defparam \b2v_inst4.pix_count_int_fast_12_LC_3_14_1 .C_ON=1'b0;
    defparam \b2v_inst4.pix_count_int_fast_12_LC_3_14_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst4.pix_count_int_fast_12_LC_3_14_1 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \b2v_inst4.pix_count_int_fast_12_LC_3_14_1  (
            .in0(N__14069),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14753),
            .lcout(b2v_inst4_pix_count_int_fast_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34517),
            .ce(),
            .sr(N__38054));
    defparam \b2v_inst4.pix_count_int_2_LC_3_14_2 .C_ON=1'b0;
    defparam \b2v_inst4.pix_count_int_2_LC_3_14_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst4.pix_count_int_2_LC_3_14_2 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \b2v_inst4.pix_count_int_2_LC_3_14_2  (
            .in0(N__14754),
            .in1(N__14008),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(SYNTHESIZED_WIRE_4_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34517),
            .ce(),
            .sr(N__38054));
    defparam \b2v_inst4.pix_count_int_6_LC_3_14_3 .C_ON=1'b0;
    defparam \b2v_inst4.pix_count_int_6_LC_3_14_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst4.pix_count_int_6_LC_3_14_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \b2v_inst4.pix_count_int_6_LC_3_14_3  (
            .in0(_gnd_net_),
            .in1(N__14751),
            .in2(_gnd_net_),
            .in3(N__13948),
            .lcout(SYNTHESIZED_WIRE_4_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34517),
            .ce(),
            .sr(N__38054));
    defparam \b2v_inst.state_19_LC_3_14_4 .C_ON=1'b0;
    defparam \b2v_inst.state_19_LC_3_14_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.state_19_LC_3_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.state_19_LC_3_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30977),
            .lcout(\b2v_inst.stateZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34517),
            .ce(),
            .sr(N__38054));
    defparam \b2v_inst.state_32_rep1_LC_3_14_5 .C_ON=1'b0;
    defparam \b2v_inst.state_32_rep1_LC_3_14_5 .SEQ_MODE=4'b1011;
    defparam \b2v_inst.state_32_rep1_LC_3_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.state_32_rep1_LC_3_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21269),
            .lcout(\b2v_inst.state_32_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34517),
            .ce(),
            .sr(N__38054));
    defparam \b2v_inst4.state_0_LC_3_14_6 .C_ON=1'b0;
    defparam \b2v_inst4.state_0_LC_3_14_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst4.state_0_LC_3_14_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \b2v_inst4.state_0_LC_3_14_6  (
            .in0(_gnd_net_),
            .in1(N__14895),
            .in2(_gnd_net_),
            .in3(N__14875),
            .lcout(\b2v_inst4.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34517),
            .ce(),
            .sr(N__38054));
    defparam \b2v_inst4.pix_count_int_1_LC_3_14_7 .C_ON=1'b0;
    defparam \b2v_inst4.pix_count_int_1_LC_3_14_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst4.pix_count_int_1_LC_3_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst4.pix_count_int_1_LC_3_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14032),
            .lcout(SYNTHESIZED_WIRE_4_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34517),
            .ce(),
            .sr(N__38054));
    defparam \b2v_inst4.pix_count_int_RNIIJDN1_17_LC_3_15_5 .C_ON=1'b0;
    defparam \b2v_inst4.pix_count_int_RNIIJDN1_17_LC_3_15_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst4.pix_count_int_RNIIJDN1_17_LC_3_15_5 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \b2v_inst4.pix_count_int_RNIIJDN1_17_LC_3_15_5  (
            .in0(N__17490),
            .in1(N__17594),
            .in2(N__17723),
            .in3(N__17444),
            .lcout(\b2v_inst4.un1_pix_count_int_0_sqmuxa_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.ignorar_ancho_1_RNO_1_LC_5_9_6 .C_ON=1'b0;
    defparam \b2v_inst.ignorar_ancho_1_RNO_1_LC_5_9_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.ignorar_ancho_1_RNO_1_LC_5_9_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \b2v_inst.ignorar_ancho_1_RNO_1_LC_5_9_6  (
            .in0(_gnd_net_),
            .in1(N__13774),
            .in2(_gnd_net_),
            .in3(N__13760),
            .lcout(\b2v_inst.ignorar_ancho_1_RNOZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.cuenta_pixel_RNI70MJ1_0_LC_5_10_0 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_pixel_RNI70MJ1_0_LC_5_10_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.cuenta_pixel_RNI70MJ1_0_LC_5_10_0 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \b2v_inst.cuenta_pixel_RNI70MJ1_0_LC_5_10_0  (
            .in0(N__13781),
            .in1(_gnd_net_),
            .in2(N__13919),
            .in3(N__13759),
            .lcout(\b2v_inst.cuenta_pixel_5_i_a2_0_2_5 ),
            .ltout(\b2v_inst.cuenta_pixel_5_i_a2_0_2_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.ignorar_anterior_RNO_1_LC_5_10_1 .C_ON=1'b0;
    defparam \b2v_inst.ignorar_anterior_RNO_1_LC_5_10_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.ignorar_anterior_RNO_1_LC_5_10_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst.ignorar_anterior_RNO_1_LC_5_10_1  (
            .in0(N__28205),
            .in1(N__13605),
            .in2(N__13712),
            .in3(N__13656),
            .lcout(\b2v_inst.un1_state_36_0_sn ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un1_cuenta_pixel_cry_1_c_RNIILR31_LC_5_10_2 .C_ON=1'b0;
    defparam \b2v_inst.un1_cuenta_pixel_cry_1_c_RNIILR31_LC_5_10_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un1_cuenta_pixel_cry_1_c_RNIILR31_LC_5_10_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \b2v_inst.un1_cuenta_pixel_cry_1_c_RNIILR31_LC_5_10_2  (
            .in0(_gnd_net_),
            .in1(N__13689),
            .in2(_gnd_net_),
            .in3(N__13671),
            .lcout(\b2v_inst.cuenta_pixel_5_i_a2_0_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.cuenta_pixel_2_LC_5_10_3 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_pixel_2_LC_5_10_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.cuenta_pixel_2_LC_5_10_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst.cuenta_pixel_2_LC_5_10_3  (
            .in0(N__13691),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst.cuenta_pixelZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34495),
            .ce(N__13852),
            .sr(N__38045));
    defparam \b2v_inst.cuenta_pixel_3_LC_5_10_4 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_pixel_3_LC_5_10_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.cuenta_pixel_3_LC_5_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.cuenta_pixel_3_LC_5_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13675),
            .lcout(\b2v_inst.cuenta_pixelZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34495),
            .ce(N__13852),
            .sr(N__38045));
    defparam \b2v_inst.ignorar_ancho_1_RNO_2_LC_5_10_5 .C_ON=1'b0;
    defparam \b2v_inst.ignorar_ancho_1_RNO_2_LC_5_10_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.ignorar_ancho_1_RNO_2_LC_5_10_5 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \b2v_inst.ignorar_ancho_1_RNO_2_LC_5_10_5  (
            .in0(N__13690),
            .in1(N__13914),
            .in2(N__13676),
            .in3(N__13655),
            .lcout(\b2v_inst.ignorar_ancho_1_RNOZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.cuenta_pixel_5_LC_5_10_6 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_pixel_5_LC_5_10_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.cuenta_pixel_5_LC_5_10_6 .LUT_INIT=16'b0010101010101010;
    LogicCell40 \b2v_inst.cuenta_pixel_5_LC_5_10_6  (
            .in0(N__13657),
            .in1(N__13630),
            .in2(N__13612),
            .in3(N__14543),
            .lcout(\b2v_inst.cuenta_pixelZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34495),
            .ce(N__13852),
            .sr(N__38045));
    defparam \b2v_inst.cuenta_pixel_4_LC_5_10_7 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_pixel_4_LC_5_10_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.cuenta_pixel_4_LC_5_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.cuenta_pixel_4_LC_5_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13918),
            .lcout(\b2v_inst.cuenta_pixelZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34495),
            .ce(N__13852),
            .sr(N__38045));
    defparam \b2v_inst.un7_pix_count_int_0_I_9_c_RNO_LC_5_11_0 .C_ON=1'b0;
    defparam \b2v_inst.un7_pix_count_int_0_I_9_c_RNO_LC_5_11_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un7_pix_count_int_0_I_9_c_RNO_LC_5_11_0 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \b2v_inst.un7_pix_count_int_0_I_9_c_RNO_LC_5_11_0  (
            .in0(N__15596),
            .in1(N__15342),
            .in2(N__13871),
            .in3(N__13877),
            .lcout(\b2v_inst.un7_pix_count_int_0_I_9_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.pix_count_anterior_10_LC_5_11_1 .C_ON=1'b0;
    defparam \b2v_inst.pix_count_anterior_10_LC_5_11_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.pix_count_anterior_10_LC_5_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.pix_count_anterior_10_LC_5_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15597),
            .lcout(\b2v_inst.pix_count_anteriorZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34477),
            .ce(N__13847),
            .sr(N__38051));
    defparam \b2v_inst.pix_count_anterior_11_LC_5_11_2 .C_ON=1'b0;
    defparam \b2v_inst.pix_count_anterior_11_LC_5_11_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.pix_count_anterior_11_LC_5_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.pix_count_anterior_11_LC_5_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15343),
            .lcout(\b2v_inst.pix_count_anteriorZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34477),
            .ce(N__13847),
            .sr(N__38051));
    defparam \b2v_inst1.r_Clk_Count_RNIGMPV1_0_2_LC_5_11_4 .C_ON=1'b0;
    defparam \b2v_inst1.r_Clk_Count_RNIGMPV1_0_2_LC_5_11_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_Clk_Count_RNIGMPV1_0_2_LC_5_11_4 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \b2v_inst1.r_Clk_Count_RNIGMPV1_0_2_LC_5_11_4  (
            .in0(N__22634),
            .in1(N__22893),
            .in2(N__16913),
            .in3(N__16541),
            .lcout(\b2v_inst1.r_RX_Byte_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.pix_count_anterior_17_LC_5_12_2 .C_ON=1'b0;
    defparam \b2v_inst.pix_count_anterior_17_LC_5_12_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.pix_count_anterior_17_LC_5_12_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst.pix_count_anterior_17_LC_5_12_2  (
            .in0(N__17437),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst.pix_count_anteriorZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34496),
            .ce(N__13853),
            .sr(N__38055));
    defparam \b2v_inst.state_RNO_17_29_LC_5_12_5 .C_ON=1'b0;
    defparam \b2v_inst.state_RNO_17_29_LC_5_12_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNO_17_29_LC_5_12_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \b2v_inst.state_RNO_17_29_LC_5_12_5  (
            .in0(N__28202),
            .in1(N__17713),
            .in2(_gnd_net_),
            .in3(N__17592),
            .lcout(\b2v_inst.N_4_i_i_a6_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.ignorar_anterior_RNO_0_LC_5_12_7 .C_ON=1'b0;
    defparam \b2v_inst.ignorar_anterior_RNO_0_LC_5_12_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.ignorar_anterior_RNO_0_LC_5_12_7 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \b2v_inst.ignorar_anterior_RNO_0_LC_5_12_7  (
            .in0(N__28203),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26004),
            .lcout(\b2v_inst.un1_state_36_0_rn_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst4.pix_count_int_RNI0EPT_0_LC_5_13_0 .C_ON=1'b1;
    defparam \b2v_inst4.pix_count_int_RNI0EPT_0_LC_5_13_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst4.pix_count_int_RNI0EPT_0_LC_5_13_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst4.pix_count_int_RNI0EPT_0_LC_5_13_0  (
            .in0(_gnd_net_),
            .in1(N__15281),
            .in2(N__28760),
            .in3(N__28751),
            .lcout(\b2v_inst4.pix_count_int_RNI0EPTZ0Z_0 ),
            .ltout(),
            .carryin(bfn_5_13_0_),
            .carryout(\b2v_inst4.un1_pix_count_int_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst4.un1_pix_count_int_cry_0_c_RNIIC2I_LC_5_13_1 .C_ON=1'b1;
    defparam \b2v_inst4.un1_pix_count_int_cry_0_c_RNIIC2I_LC_5_13_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst4.un1_pix_count_int_cry_0_c_RNIIC2I_LC_5_13_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst4.un1_pix_count_int_cry_0_c_RNIIC2I_LC_5_13_1  (
            .in0(_gnd_net_),
            .in1(N__15197),
            .in2(_gnd_net_),
            .in3(N__14015),
            .lcout(\b2v_inst4.un1_pix_count_int_cry_0_c_RNIIC2IZ0 ),
            .ltout(),
            .carryin(\b2v_inst4.un1_pix_count_int_cry_0 ),
            .carryout(\b2v_inst4.un1_pix_count_int_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst4.un1_pix_count_int_cry_1_c_RNIKF3I_LC_5_13_2 .C_ON=1'b1;
    defparam \b2v_inst4.un1_pix_count_int_cry_1_c_RNIKF3I_LC_5_13_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst4.un1_pix_count_int_cry_1_c_RNIKF3I_LC_5_13_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst4.un1_pix_count_int_cry_1_c_RNIKF3I_LC_5_13_2  (
            .in0(_gnd_net_),
            .in1(N__15140),
            .in2(_gnd_net_),
            .in3(N__13991),
            .lcout(\b2v_inst4.un1_pix_count_int_cry_1_c_RNIKF3IZ0 ),
            .ltout(),
            .carryin(\b2v_inst4.un1_pix_count_int_cry_1 ),
            .carryout(\b2v_inst4.un1_pix_count_int_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst4.un1_pix_count_int_cry_2_c_RNIMI4I_LC_5_13_3 .C_ON=1'b1;
    defparam \b2v_inst4.un1_pix_count_int_cry_2_c_RNIMI4I_LC_5_13_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst4.un1_pix_count_int_cry_2_c_RNIMI4I_LC_5_13_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst4.un1_pix_count_int_cry_2_c_RNIMI4I_LC_5_13_3  (
            .in0(_gnd_net_),
            .in1(N__15238),
            .in2(_gnd_net_),
            .in3(N__13976),
            .lcout(\b2v_inst4.un1_pix_count_int_cry_2_c_RNIMI4IZ0 ),
            .ltout(),
            .carryin(\b2v_inst4.un1_pix_count_int_cry_2 ),
            .carryout(\b2v_inst4.un1_pix_count_int_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst4.pix_count_int_4_LC_5_13_4 .C_ON=1'b1;
    defparam \b2v_inst4.pix_count_int_4_LC_5_13_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst4.pix_count_int_4_LC_5_13_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst4.pix_count_int_4_LC_5_13_4  (
            .in0(_gnd_net_),
            .in1(N__16727),
            .in2(_gnd_net_),
            .in3(N__13973),
            .lcout(SYNTHESIZED_WIRE_4_4),
            .ltout(),
            .carryin(\b2v_inst4.un1_pix_count_int_cry_3 ),
            .carryout(\b2v_inst4.un1_pix_count_int_cry_4 ),
            .clk(N__34502),
            .ce(),
            .sr(N__38059));
    defparam \b2v_inst4.un1_pix_count_int_cry_4_c_RNIQO6I_LC_5_13_5 .C_ON=1'b1;
    defparam \b2v_inst4.un1_pix_count_int_cry_4_c_RNIQO6I_LC_5_13_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst4.un1_pix_count_int_cry_4_c_RNIQO6I_LC_5_13_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst4.un1_pix_count_int_cry_4_c_RNIQO6I_LC_5_13_5  (
            .in0(_gnd_net_),
            .in1(N__15827),
            .in2(_gnd_net_),
            .in3(N__13955),
            .lcout(\b2v_inst4.un1_pix_count_int_cry_4_c_RNIQO6IZ0 ),
            .ltout(),
            .carryin(\b2v_inst4.un1_pix_count_int_cry_4 ),
            .carryout(\b2v_inst4.un1_pix_count_int_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst4.un1_pix_count_int_cry_5_c_RNISR7I_LC_5_13_6 .C_ON=1'b1;
    defparam \b2v_inst4.un1_pix_count_int_cry_5_c_RNISR7I_LC_5_13_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst4.un1_pix_count_int_cry_5_c_RNISR7I_LC_5_13_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst4.un1_pix_count_int_cry_5_c_RNISR7I_LC_5_13_6  (
            .in0(_gnd_net_),
            .in1(N__15877),
            .in2(_gnd_net_),
            .in3(N__13931),
            .lcout(\b2v_inst4.un1_pix_count_int_cry_5_c_RNISR7IZ0 ),
            .ltout(),
            .carryin(\b2v_inst4.un1_pix_count_int_cry_5 ),
            .carryout(\b2v_inst4.un1_pix_count_int_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst4.pix_count_int_7_LC_5_13_7 .C_ON=1'b1;
    defparam \b2v_inst4.pix_count_int_7_LC_5_13_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst4.pix_count_int_7_LC_5_13_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst4.pix_count_int_7_LC_5_13_7  (
            .in0(_gnd_net_),
            .in1(N__16821),
            .in2(_gnd_net_),
            .in3(N__13928),
            .lcout(SYNTHESIZED_WIRE_4_7),
            .ltout(),
            .carryin(\b2v_inst4.un1_pix_count_int_cry_6 ),
            .carryout(\b2v_inst4.un1_pix_count_int_cry_7 ),
            .clk(N__34502),
            .ce(),
            .sr(N__38059));
    defparam \b2v_inst4.pix_count_int_8_LC_5_14_0 .C_ON=1'b1;
    defparam \b2v_inst4.pix_count_int_8_LC_5_14_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst4.pix_count_int_8_LC_5_14_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst4.pix_count_int_8_LC_5_14_0  (
            .in0(N__14790),
            .in1(N__15477),
            .in2(_gnd_net_),
            .in3(N__13925),
            .lcout(SYNTHESIZED_WIRE_4_8),
            .ltout(),
            .carryin(bfn_5_14_0_),
            .carryout(\b2v_inst4.un1_pix_count_int_cry_8 ),
            .clk(N__34508),
            .ce(),
            .sr(N__38062));
    defparam \b2v_inst4.un1_pix_count_int_cry_8_c_RNI25BI_LC_5_14_1 .C_ON=1'b1;
    defparam \b2v_inst4.un1_pix_count_int_cry_8_c_RNI25BI_LC_5_14_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst4.un1_pix_count_int_cry_8_c_RNI25BI_LC_5_14_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst4.un1_pix_count_int_cry_8_c_RNI25BI_LC_5_14_1  (
            .in0(_gnd_net_),
            .in1(N__15564),
            .in2(_gnd_net_),
            .in3(N__13922),
            .lcout(\b2v_inst4.un1_pix_count_int_cry_8_c_RNI25BIZ0 ),
            .ltout(),
            .carryin(\b2v_inst4.un1_pix_count_int_cry_8 ),
            .carryout(\b2v_inst4.un1_pix_count_int_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst4.un1_pix_count_int_cry_9_c_RNIB86J_LC_5_14_2 .C_ON=1'b1;
    defparam \b2v_inst4.un1_pix_count_int_cry_9_c_RNIB86J_LC_5_14_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst4.un1_pix_count_int_cry_9_c_RNIB86J_LC_5_14_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst4.un1_pix_count_int_cry_9_c_RNIB86J_LC_5_14_2  (
            .in0(_gnd_net_),
            .in1(N__15616),
            .in2(_gnd_net_),
            .in3(N__14075),
            .lcout(\b2v_inst4.un1_pix_count_int_cry_9_c_RNIB86JZ0 ),
            .ltout(),
            .carryin(\b2v_inst4.un1_pix_count_int_cry_9 ),
            .carryout(\b2v_inst4.un1_pix_count_int_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst4.un1_pix_count_int_cry_10_c_RNIKMUJ_LC_5_14_3 .C_ON=1'b1;
    defparam \b2v_inst4.un1_pix_count_int_cry_10_c_RNIKMUJ_LC_5_14_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst4.un1_pix_count_int_cry_10_c_RNIKMUJ_LC_5_14_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst4.un1_pix_count_int_cry_10_c_RNIKMUJ_LC_5_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15356),
            .in3(N__14072),
            .lcout(\b2v_inst4.un1_pix_count_int_cry_10_c_RNIKMUJZ0 ),
            .ltout(),
            .carryin(\b2v_inst4.un1_pix_count_int_cry_10 ),
            .carryout(\b2v_inst4.un1_pix_count_int_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst4.un1_pix_count_int_cry_11_c_RNIMPVJ_LC_5_14_4 .C_ON=1'b1;
    defparam \b2v_inst4.un1_pix_count_int_cry_11_c_RNIMPVJ_LC_5_14_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst4.un1_pix_count_int_cry_11_c_RNIMPVJ_LC_5_14_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst4.un1_pix_count_int_cry_11_c_RNIMPVJ_LC_5_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15398),
            .in3(N__14057),
            .lcout(\b2v_inst4.un1_pix_count_int_cry_11_c_RNIMPVJZ0 ),
            .ltout(),
            .carryin(\b2v_inst4.un1_pix_count_int_cry_11 ),
            .carryout(\b2v_inst4.un1_pix_count_int_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst4.pix_count_int_13_LC_5_14_5 .C_ON=1'b1;
    defparam \b2v_inst4.pix_count_int_13_LC_5_14_5 .SEQ_MODE=4'b1010;
    defparam \b2v_inst4.pix_count_int_13_LC_5_14_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst4.pix_count_int_13_LC_5_14_5  (
            .in0(_gnd_net_),
            .in1(N__16473),
            .in2(_gnd_net_),
            .in3(N__14054),
            .lcout(SYNTHESIZED_WIRE_4_13),
            .ltout(),
            .carryin(\b2v_inst4.un1_pix_count_int_cry_12 ),
            .carryout(\b2v_inst4.un1_pix_count_int_cry_13 ),
            .clk(N__34508),
            .ce(),
            .sr(N__38062));
    defparam \b2v_inst4.pix_count_int_14_LC_5_14_6 .C_ON=1'b1;
    defparam \b2v_inst4.pix_count_int_14_LC_5_14_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst4.pix_count_int_14_LC_5_14_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst4.pix_count_int_14_LC_5_14_6  (
            .in0(_gnd_net_),
            .in1(N__16354),
            .in2(_gnd_net_),
            .in3(N__14051),
            .lcout(SYNTHESIZED_WIRE_4_14),
            .ltout(),
            .carryin(\b2v_inst4.un1_pix_count_int_cry_13 ),
            .carryout(\b2v_inst4.un1_pix_count_int_cry_14 ),
            .clk(N__34508),
            .ce(),
            .sr(N__38062));
    defparam \b2v_inst4.pix_count_int_15_LC_5_14_7 .C_ON=1'b1;
    defparam \b2v_inst4.pix_count_int_15_LC_5_14_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst4.pix_count_int_15_LC_5_14_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst4.pix_count_int_15_LC_5_14_7  (
            .in0(_gnd_net_),
            .in1(N__16407),
            .in2(_gnd_net_),
            .in3(N__14048),
            .lcout(SYNTHESIZED_WIRE_4_15),
            .ltout(),
            .carryin(\b2v_inst4.un1_pix_count_int_cry_14 ),
            .carryout(\b2v_inst4.un1_pix_count_int_cry_15 ),
            .clk(N__34508),
            .ce(),
            .sr(N__38062));
    defparam \b2v_inst4.pix_count_int_16_LC_5_15_0 .C_ON=1'b1;
    defparam \b2v_inst4.pix_count_int_16_LC_5_15_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst4.pix_count_int_16_LC_5_15_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst4.pix_count_int_16_LC_5_15_0  (
            .in0(N__14788),
            .in1(N__17598),
            .in2(_gnd_net_),
            .in3(N__14045),
            .lcout(SYNTHESIZED_WIRE_4_16),
            .ltout(),
            .carryin(bfn_5_15_0_),
            .carryout(\b2v_inst4.un1_pix_count_int_cry_16 ),
            .clk(N__34513),
            .ce(),
            .sr(N__38065));
    defparam \b2v_inst4.pix_count_int_17_LC_5_15_1 .C_ON=1'b1;
    defparam \b2v_inst4.pix_count_int_17_LC_5_15_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst4.pix_count_int_17_LC_5_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst4.pix_count_int_17_LC_5_15_1  (
            .in0(_gnd_net_),
            .in1(N__17432),
            .in2(_gnd_net_),
            .in3(N__14042),
            .lcout(SYNTHESIZED_WIRE_4_17),
            .ltout(),
            .carryin(\b2v_inst4.un1_pix_count_int_cry_16 ),
            .carryout(\b2v_inst4.un1_pix_count_int_cry_17 ),
            .clk(N__34513),
            .ce(),
            .sr(N__38065));
    defparam \b2v_inst4.pix_count_int_18_LC_5_15_2 .C_ON=1'b1;
    defparam \b2v_inst4.pix_count_int_18_LC_5_15_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst4.pix_count_int_18_LC_5_15_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst4.pix_count_int_18_LC_5_15_2  (
            .in0(_gnd_net_),
            .in1(N__17484),
            .in2(_gnd_net_),
            .in3(N__14039),
            .lcout(SYNTHESIZED_WIRE_4_18),
            .ltout(),
            .carryin(\b2v_inst4.un1_pix_count_int_cry_17 ),
            .carryout(\b2v_inst4.un1_pix_count_int_cry_18 ),
            .clk(N__34513),
            .ce(),
            .sr(N__38065));
    defparam \b2v_inst4.pix_count_int_19_LC_5_15_3 .C_ON=1'b0;
    defparam \b2v_inst4.pix_count_int_19_LC_5_15_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst4.pix_count_int_19_LC_5_15_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst4.pix_count_int_19_LC_5_15_3  (
            .in0(N__14787),
            .in1(N__17695),
            .in2(_gnd_net_),
            .in3(N__14456),
            .lcout(SYNTHESIZED_WIRE_4_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34513),
            .ce(),
            .sr(N__38065));
    defparam \b2v_inst1.r_RX_Byte_1_LC_5_16_4 .C_ON=1'b0;
    defparam \b2v_inst1.r_RX_Byte_1_LC_5_16_4 .SEQ_MODE=4'b1000;
    defparam \b2v_inst1.r_RX_Byte_1_LC_5_16_4 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \b2v_inst1.r_RX_Byte_1_LC_5_16_4  (
            .in0(N__27018),
            .in1(N__17299),
            .in2(_gnd_net_),
            .in3(N__14945),
            .lcout(SYNTHESIZED_WIRE_10_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34522),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_RNI2OT15_1_LC_5_18_3 .C_ON=1'b0;
    defparam \b2v_inst.indice_RNI2OT15_1_LC_5_18_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_RNI2OT15_1_LC_5_18_3 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \b2v_inst.indice_RNI2OT15_1_LC_5_18_3  (
            .in0(N__21663),
            .in1(N__35217),
            .in2(N__20168),
            .in3(N__38665),
            .lcout(SYNTHESIZED_WIRE_12_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_RNIKAU15_7_LC_5_18_4 .C_ON=1'b0;
    defparam \b2v_inst.indice_RNIKAU15_7_LC_5_18_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_RNIKAU15_7_LC_5_18_4 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \b2v_inst.indice_RNIKAU15_7_LC_5_18_4  (
            .in0(N__35218),
            .in1(N__21664),
            .in2(N__18893),
            .in3(N__38870),
            .lcout(SYNTHESIZED_WIRE_12_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_RNIVKT15_0_LC_5_18_5 .C_ON=1'b0;
    defparam \b2v_inst.indice_RNIVKT15_0_LC_5_18_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_RNIVKT15_0_LC_5_18_5 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \b2v_inst.indice_RNIVKT15_0_LC_5_18_5  (
            .in0(N__21665),
            .in1(N__39317),
            .in2(N__20384),
            .in3(N__35219),
            .lcout(SYNTHESIZED_WIRE_12_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_RNINDU15_8_LC_5_19_2 .C_ON=1'b0;
    defparam \b2v_inst.indice_RNINDU15_8_LC_5_19_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_RNINDU15_8_LC_5_19_2 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \b2v_inst.indice_RNINDU15_8_LC_5_19_2  (
            .in0(N__35237),
            .in1(N__18569),
            .in2(N__39101),
            .in3(N__21662),
            .lcout(SYNTHESIZED_WIRE_12_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un2_dir_mem_3_cry_0_c_LC_6_5_0 .C_ON=1'b1;
    defparam \b2v_inst.un2_dir_mem_3_cry_0_c_LC_6_5_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un2_dir_mem_3_cry_0_c_LC_6_5_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.un2_dir_mem_3_cry_0_c_LC_6_5_0  (
            .in0(_gnd_net_),
            .in1(N__35701),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_5_0_),
            .carryout(\b2v_inst.un2_dir_mem_3_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_3_RNO_0_6_LC_6_5_1 .C_ON=1'b1;
    defparam \b2v_inst.dir_mem_3_RNO_0_6_LC_6_5_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_3_RNO_0_6_LC_6_5_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.dir_mem_3_RNO_0_6_LC_6_5_1  (
            .in0(_gnd_net_),
            .in1(N__38337),
            .in2(_gnd_net_),
            .in3(N__14081),
            .lcout(\b2v_inst.dir_mem_3_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\b2v_inst.un2_dir_mem_3_cry_0 ),
            .carryout(\b2v_inst.un2_dir_mem_3_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_3_RNO_0_7_LC_6_5_2 .C_ON=1'b1;
    defparam \b2v_inst.dir_mem_3_RNO_0_7_LC_6_5_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_3_RNO_0_7_LC_6_5_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst.dir_mem_3_RNO_0_7_LC_6_5_2  (
            .in0(_gnd_net_),
            .in1(N__38836),
            .in2(N__37303),
            .in3(N__14078),
            .lcout(\b2v_inst.dir_mem_3_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(\b2v_inst.un2_dir_mem_3_cry_1 ),
            .carryout(\b2v_inst.un2_dir_mem_3_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_3_RNO_0_8_LC_6_5_3 .C_ON=1'b1;
    defparam \b2v_inst.dir_mem_3_RNO_0_8_LC_6_5_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_3_RNO_0_8_LC_6_5_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.dir_mem_3_RNO_0_8_LC_6_5_3  (
            .in0(_gnd_net_),
            .in1(N__39058),
            .in2(_gnd_net_),
            .in3(N__14480),
            .lcout(\b2v_inst.dir_mem_3_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(\b2v_inst.un2_dir_mem_3_cry_2 ),
            .carryout(\b2v_inst.un2_dir_mem_3_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_3_RNO_0_9_LC_6_5_4 .C_ON=1'b1;
    defparam \b2v_inst.dir_mem_3_RNO_0_9_LC_6_5_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_3_RNO_0_9_LC_6_5_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.dir_mem_3_RNO_0_9_LC_6_5_4  (
            .in0(_gnd_net_),
            .in1(N__35915),
            .in2(_gnd_net_),
            .in3(N__14477),
            .lcout(\b2v_inst.dir_mem_3_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(\b2v_inst.un2_dir_mem_3_cry_3 ),
            .carryout(\b2v_inst.un2_dir_mem_3_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_3_RNO_0_10_LC_6_5_5 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_3_RNO_0_10_LC_6_5_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_3_RNO_0_10_LC_6_5_5 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \b2v_inst.dir_mem_3_RNO_0_10_LC_6_5_5  (
            .in0(N__36747),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14474),
            .lcout(\b2v_inst.dir_mem_3_RNO_0Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un1_indice_cry_1_c_LC_6_6_0 .C_ON=1'b1;
    defparam \b2v_inst.un1_indice_cry_1_c_LC_6_6_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un1_indice_cry_1_c_LC_6_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.un1_indice_cry_1_c_LC_6_6_0  (
            .in0(_gnd_net_),
            .in1(N__39273),
            .in2(N__38603),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_6_0_),
            .carryout(\b2v_inst.un1_indice_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un1_indice_cry_1_c_RNIUSJG_LC_6_6_1 .C_ON=1'b1;
    defparam \b2v_inst.un1_indice_cry_1_c_RNIUSJG_LC_6_6_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un1_indice_cry_1_c_RNIUSJG_LC_6_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.un1_indice_cry_1_c_RNIUSJG_LC_6_6_1  (
            .in0(_gnd_net_),
            .in1(N__36043),
            .in2(_gnd_net_),
            .in3(N__14471),
            .lcout(\b2v_inst.un1_indice_cry_1_c_RNIUSJGZ0 ),
            .ltout(),
            .carryin(\b2v_inst.un1_indice_cry_1 ),
            .carryout(\b2v_inst.un1_indice_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un1_indice_cry_2_c_RNI00LG_LC_6_6_2 .C_ON=1'b1;
    defparam \b2v_inst.un1_indice_cry_2_c_RNI00LG_LC_6_6_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un1_indice_cry_2_c_RNI00LG_LC_6_6_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.un1_indice_cry_2_c_RNI00LG_LC_6_6_2  (
            .in0(_gnd_net_),
            .in1(N__36512),
            .in2(_gnd_net_),
            .in3(N__14468),
            .lcout(\b2v_inst.un1_indice_cry_2_c_RNI00LGZ0 ),
            .ltout(),
            .carryin(\b2v_inst.un1_indice_cry_2 ),
            .carryout(\b2v_inst.un1_indice_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un1_indice_cry_3_c_RNI23MG_LC_6_6_3 .C_ON=1'b1;
    defparam \b2v_inst.un1_indice_cry_3_c_RNI23MG_LC_6_6_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un1_indice_cry_3_c_RNI23MG_LC_6_6_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.un1_indice_cry_3_c_RNI23MG_LC_6_6_3  (
            .in0(_gnd_net_),
            .in1(N__36363),
            .in2(_gnd_net_),
            .in3(N__14465),
            .lcout(\b2v_inst.un1_indice_cry_3_c_RNI23MGZ0 ),
            .ltout(),
            .carryin(\b2v_inst.un1_indice_cry_3 ),
            .carryout(\b2v_inst.un1_indice_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un1_indice_cry_4_c_RNI46NG_LC_6_6_4 .C_ON=1'b1;
    defparam \b2v_inst.un1_indice_cry_4_c_RNI46NG_LC_6_6_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un1_indice_cry_4_c_RNI46NG_LC_6_6_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.un1_indice_cry_4_c_RNI46NG_LC_6_6_4  (
            .in0(_gnd_net_),
            .in1(N__35710),
            .in2(_gnd_net_),
            .in3(N__14462),
            .lcout(\b2v_inst.un1_indice_cry_4_c_RNI46NGZ0 ),
            .ltout(),
            .carryin(\b2v_inst.un1_indice_cry_4 ),
            .carryout(\b2v_inst.un1_indice_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un1_indice_cry_5_c_RNI69OG_LC_6_6_5 .C_ON=1'b1;
    defparam \b2v_inst.un1_indice_cry_5_c_RNI69OG_LC_6_6_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un1_indice_cry_5_c_RNI69OG_LC_6_6_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.un1_indice_cry_5_c_RNI69OG_LC_6_6_5  (
            .in0(_gnd_net_),
            .in1(N__38326),
            .in2(_gnd_net_),
            .in3(N__14459),
            .lcout(\b2v_inst.un1_indice_cry_5_c_RNI69OGZ0 ),
            .ltout(),
            .carryin(\b2v_inst.un1_indice_cry_5 ),
            .carryout(\b2v_inst.un1_indice_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un1_indice_cry_6_c_RNI8CPG_LC_6_6_6 .C_ON=1'b1;
    defparam \b2v_inst.un1_indice_cry_6_c_RNI8CPG_LC_6_6_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un1_indice_cry_6_c_RNI8CPG_LC_6_6_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.un1_indice_cry_6_c_RNI8CPG_LC_6_6_6  (
            .in0(_gnd_net_),
            .in1(N__38861),
            .in2(_gnd_net_),
            .in3(N__14507),
            .lcout(\b2v_inst.dir_mem_316lto7 ),
            .ltout(),
            .carryin(\b2v_inst.un1_indice_cry_6 ),
            .carryout(\b2v_inst.un1_indice_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un1_indice_cry_7_c_RNIAFQG_LC_6_6_7 .C_ON=1'b1;
    defparam \b2v_inst.un1_indice_cry_7_c_RNIAFQG_LC_6_6_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un1_indice_cry_7_c_RNIAFQG_LC_6_6_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.un1_indice_cry_7_c_RNIAFQG_LC_6_6_7  (
            .in0(_gnd_net_),
            .in1(N__39079),
            .in2(_gnd_net_),
            .in3(N__14504),
            .lcout(\b2v_inst.un1_indice_cry_7_c_RNIAFQGZ0 ),
            .ltout(),
            .carryin(\b2v_inst.un1_indice_cry_7 ),
            .carryout(\b2v_inst.un1_indice_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un1_indice_cry_8_c_RNICIRG_LC_6_7_0 .C_ON=1'b1;
    defparam \b2v_inst.un1_indice_cry_8_c_RNICIRG_LC_6_7_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un1_indice_cry_8_c_RNICIRG_LC_6_7_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.un1_indice_cry_8_c_RNICIRG_LC_6_7_0  (
            .in0(_gnd_net_),
            .in1(N__35938),
            .in2(_gnd_net_),
            .in3(N__14501),
            .lcout(\b2v_inst.un1_indice_cry_8_c_RNICIRGZ0 ),
            .ltout(),
            .carryin(bfn_6_7_0_),
            .carryout(\b2v_inst.un1_indice_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un1_indice_cry_9_c_RNILAJP_LC_6_7_1 .C_ON=1'b1;
    defparam \b2v_inst.un1_indice_cry_9_c_RNILAJP_LC_6_7_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un1_indice_cry_9_c_RNILAJP_LC_6_7_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst.un1_indice_cry_9_c_RNILAJP_LC_6_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__36746),
            .in3(N__14498),
            .lcout(\b2v_inst.un1_indice_cry_9_c_RNILAJPZ0 ),
            .ltout(),
            .carryin(\b2v_inst.un1_indice_cry_9 ),
            .carryout(\b2v_inst.un1_indice_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un1_indice_cry_10_THRU_LUT4_0_LC_6_7_2 .C_ON=1'b0;
    defparam \b2v_inst.un1_indice_cry_10_THRU_LUT4_0_LC_6_7_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un1_indice_cry_10_THRU_LUT4_0_LC_6_7_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.un1_indice_cry_10_THRU_LUT4_0_LC_6_7_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14495),
            .lcout(\b2v_inst.un1_indice_cry_10_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.pix_data_reg_4_LC_6_8_4 .C_ON=1'b0;
    defparam \b2v_inst.pix_data_reg_4_LC_6_8_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.pix_data_reg_4_LC_6_8_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.pix_data_reg_4_LC_6_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27086),
            .lcout(\b2v_inst.pix_data_regZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34498),
            .ce(N__30243),
            .sr(N__38057));
    defparam \b2v_inst.ignorar_ancho_1_RNO_0_LC_6_10_4 .C_ON=1'b0;
    defparam \b2v_inst.ignorar_ancho_1_RNO_0_LC_6_10_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.ignorar_ancho_1_RNO_0_LC_6_10_4 .LUT_INIT=16'b0100011111001111;
    LogicCell40 \b2v_inst.ignorar_ancho_1_RNO_0_LC_6_10_4  (
            .in0(N__14492),
            .in1(N__28204),
            .in2(N__26033),
            .in3(N__14486),
            .lcout(\b2v_inst.ignorar_ancho_1_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst4.pix_count_int_9_LC_6_11_0 .C_ON=1'b0;
    defparam \b2v_inst4.pix_count_int_9_LC_6_11_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst4.pix_count_int_9_LC_6_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst4.pix_count_int_9_LC_6_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14811),
            .lcout(SYNTHESIZED_WIRE_4_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34468),
            .ce(),
            .sr(N__38052));
    defparam \b2v_inst4.pix_count_int_fast_10_LC_6_11_1 .C_ON=1'b0;
    defparam \b2v_inst4.pix_count_int_fast_10_LC_6_11_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst4.pix_count_int_fast_10_LC_6_11_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst4.pix_count_int_fast_10_LC_6_11_1  (
            .in0(N__14834),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(SYNTHESIZED_WIRE_4_fast_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34468),
            .ce(),
            .sr(N__38052));
    defparam \b2v_inst4.pix_count_int_10_LC_6_11_2 .C_ON=1'b0;
    defparam \b2v_inst4.pix_count_int_10_LC_6_11_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst4.pix_count_int_10_LC_6_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst4.pix_count_int_10_LC_6_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14832),
            .lcout(SYNTHESIZED_WIRE_4_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34468),
            .ce(),
            .sr(N__38052));
    defparam \b2v_inst4.pix_count_int_10_rep1_LC_6_11_4 .C_ON=1'b0;
    defparam \b2v_inst4.pix_count_int_10_rep1_LC_6_11_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst4.pix_count_int_10_rep1_LC_6_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst4.pix_count_int_10_rep1_LC_6_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14833),
            .lcout(SYNTHESIZED_WIRE_4_10_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34468),
            .ce(),
            .sr(N__38052));
    defparam \b2v_inst4.pix_count_int_fast_9_LC_6_11_6 .C_ON=1'b0;
    defparam \b2v_inst4.pix_count_int_fast_9_LC_6_11_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst4.pix_count_int_fast_9_LC_6_11_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst4.pix_count_int_fast_9_LC_6_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14812),
            .lcout(SYNTHESIZED_WIRE_4_fast_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34468),
            .ce(),
            .sr(N__38052));
    defparam \b2v_inst4.pix_count_int_11_LC_6_11_7 .C_ON=1'b0;
    defparam \b2v_inst4.pix_count_int_11_LC_6_11_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst4.pix_count_int_11_LC_6_11_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \b2v_inst4.pix_count_int_11_LC_6_11_7  (
            .in0(_gnd_net_),
            .in1(N__14789),
            .in2(_gnd_net_),
            .in3(N__14683),
            .lcout(SYNTHESIZED_WIRE_4_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34468),
            .ce(),
            .sr(N__38052));
    defparam \b2v_inst.un7_pix_count_int_0_I_33_c_RNIGJGQ8_LC_6_12_0 .C_ON=1'b0;
    defparam \b2v_inst.un7_pix_count_int_0_I_33_c_RNIGJGQ8_LC_6_12_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un7_pix_count_int_0_I_33_c_RNIGJGQ8_LC_6_12_0 .LUT_INIT=16'b1111001011110000;
    LogicCell40 \b2v_inst.un7_pix_count_int_0_I_33_c_RNIGJGQ8_LC_6_12_0  (
            .in0(N__17709),
            .in1(N__15410),
            .in2(N__17222),
            .in3(N__17593),
            .lcout(\b2v_inst.N_482 ),
            .ltout(\b2v_inst.N_482_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.ignorar_ancho_1_RNO_LC_6_12_1 .C_ON=1'b0;
    defparam \b2v_inst.ignorar_ancho_1_RNO_LC_6_12_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.ignorar_ancho_1_RNO_LC_6_12_1 .LUT_INIT=16'b0001001100010001;
    LogicCell40 \b2v_inst.ignorar_ancho_1_RNO_LC_6_12_1  (
            .in0(N__28184),
            .in1(N__14666),
            .in2(N__14657),
            .in3(N__14539),
            .lcout(\b2v_inst.un1_state_34_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.ignorar_ancho_1_LC_6_12_2 .C_ON=1'b0;
    defparam \b2v_inst.ignorar_ancho_1_LC_6_12_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.ignorar_ancho_1_LC_6_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.ignorar_ancho_1_LC_6_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28185),
            .lcout(\b2v_inst.ignorar_anchoZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34478),
            .ce(N__14654),
            .sr(N__38058));
    defparam \b2v_inst.cuenta_pixel_RNIBK2I2_10_LC_6_12_4 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_pixel_RNIBK2I2_10_LC_6_12_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.cuenta_pixel_RNIBK2I2_10_LC_6_12_4 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \b2v_inst.cuenta_pixel_RNIBK2I2_10_LC_6_12_4  (
            .in0(N__14645),
            .in1(N__14621),
            .in2(N__14594),
            .in3(N__14561),
            .lcout(\b2v_inst.N_325 ),
            .ltout(\b2v_inst.N_325_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.ignorar_anterior_RNO_LC_6_12_5 .C_ON=1'b0;
    defparam \b2v_inst.ignorar_anterior_RNO_LC_6_12_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.ignorar_anterior_RNO_LC_6_12_5 .LUT_INIT=16'b0010001011100010;
    LogicCell40 \b2v_inst.ignorar_anterior_RNO_LC_6_12_5  (
            .in0(N__14528),
            .in1(N__14519),
            .in2(N__14510),
            .in3(N__28514),
            .lcout(\b2v_inst.un1_state_36_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un7_pix_count_int_0_I_33_c_RNIMVIF1_LC_6_12_6 .C_ON=1'b0;
    defparam \b2v_inst.un7_pix_count_int_0_I_33_c_RNIMVIF1_LC_6_12_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un7_pix_count_int_0_I_33_c_RNIMVIF1_LC_6_12_6 .LUT_INIT=16'b1110000011111111;
    LogicCell40 \b2v_inst.un7_pix_count_int_0_I_33_c_RNIMVIF1_LC_6_12_6  (
            .in0(N__17502),
            .in1(N__17436),
            .in2(N__17727),
            .in3(N__17104),
            .lcout(\b2v_inst.un4_pix_count_intlto19_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNI9A7V8_29_LC_6_12_7 .C_ON=1'b0;
    defparam \b2v_inst.state_RNI9A7V8_29_LC_6_12_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNI9A7V8_29_LC_6_12_7 .LUT_INIT=16'b0000000010101000;
    LogicCell40 \b2v_inst.state_RNI9A7V8_29_LC_6_12_7  (
            .in0(N__28183),
            .in1(N__15409),
            .in2(N__14846),
            .in3(N__17217),
            .lcout(\b2v_inst.N_305_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.ignorar_anterior_LC_6_13_0 .C_ON=1'b0;
    defparam \b2v_inst.ignorar_anterior_LC_6_13_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.ignorar_anterior_LC_6_13_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.ignorar_anterior_LC_6_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28174),
            .lcout(\b2v_inst.ignorar_anteriorZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34488),
            .ce(N__14909),
            .sr(N__38060));
    defparam \b2v_inst1.r_RX_Byte_RNO_0_0_LC_6_14_0 .C_ON=1'b0;
    defparam \b2v_inst1.r_RX_Byte_RNO_0_0_LC_6_14_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_RX_Byte_RNO_0_0_LC_6_14_0 .LUT_INIT=16'b0000111100011101;
    LogicCell40 \b2v_inst1.r_RX_Byte_RNO_0_0_LC_6_14_0  (
            .in0(N__22832),
            .in1(N__16638),
            .in2(N__26716),
            .in3(N__15434),
            .lcout(\b2v_inst1.N_42 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.g1_0_a4_0_LC_6_14_1 .C_ON=1'b0;
    defparam \b2v_inst.g1_0_a4_0_LC_6_14_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.g1_0_a4_0_LC_6_14_1 .LUT_INIT=16'b1000100010000000;
    LogicCell40 \b2v_inst.g1_0_a4_0_LC_6_14_1  (
            .in0(N__15392),
            .in1(N__15352),
            .in2(N__15774),
            .in3(N__15319),
            .lcout(\b2v_inst.N_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst4.state_RNICJOG_0_LC_6_14_3 .C_ON=1'b0;
    defparam \b2v_inst4.state_RNICJOG_0_LC_6_14_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst4.state_RNICJOG_0_LC_6_14_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \b2v_inst4.state_RNICJOG_0_LC_6_14_3  (
            .in0(N__14896),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14864),
            .lcout(\b2v_inst4.pix_count_int_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_RX_DV_LC_6_14_4 .C_ON=1'b0;
    defparam \b2v_inst1.r_RX_DV_LC_6_14_4 .SEQ_MODE=4'b1000;
    defparam \b2v_inst1.r_RX_DV_LC_6_14_4 .LUT_INIT=16'b1010101011100000;
    LogicCell40 \b2v_inst1.r_RX_DV_LC_6_14_4  (
            .in0(N__14865),
            .in1(N__22642),
            .in2(N__22925),
            .in3(N__21165),
            .lcout(SYNTHESIZED_WIRE_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34499),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un1_state_36_0_a2_0_1_mb_1_LC_6_15_2 .C_ON=1'b0;
    defparam \b2v_inst.un1_state_36_0_a2_0_1_mb_1_LC_6_15_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un1_state_36_0_a2_0_1_mb_1_LC_6_15_2 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \b2v_inst.un1_state_36_0_a2_0_1_mb_1_LC_6_15_2  (
            .in0(_gnd_net_),
            .in1(N__17685),
            .in2(_gnd_net_),
            .in3(N__17565),
            .lcout(\b2v_inst.un1_state_36_0_a2_0_1_mbZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un4_pix_count_intlto18_0_LC_6_15_5 .C_ON=1'b0;
    defparam \b2v_inst.un4_pix_count_intlto18_0_LC_6_15_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un4_pix_count_intlto18_0_LC_6_15_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \b2v_inst.un4_pix_count_intlto18_0_LC_6_15_5  (
            .in0(_gnd_net_),
            .in1(N__17483),
            .in2(_gnd_net_),
            .in3(N__17431),
            .lcout(\b2v_inst.un4_pix_count_intlto18Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_RX_Byte_RNO_0_1_LC_6_15_7 .C_ON=1'b0;
    defparam \b2v_inst1.r_RX_Byte_RNO_0_1_LC_6_15_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_RX_Byte_RNO_0_1_LC_6_15_7 .LUT_INIT=16'b0000111100011011;
    LogicCell40 \b2v_inst1.r_RX_Byte_RNO_0_1_LC_6_15_7  (
            .in0(N__16628),
            .in1(N__22829),
            .in2(N__27022),
            .in3(N__15983),
            .lcout(\b2v_inst1.N_40 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_1_LC_7_5_0 .C_ON=1'b0;
    defparam \b2v_inst.indice_1_LC_7_5_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.indice_1_LC_7_5_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \b2v_inst.indice_1_LC_7_5_0  (
            .in0(_gnd_net_),
            .in1(N__22106),
            .in2(_gnd_net_),
            .in3(N__16245),
            .lcout(\b2v_inst.indiceZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34510),
            .ce(N__22033),
            .sr(N__38068));
    defparam \b2v_inst.indice_2_LC_7_5_1 .C_ON=1'b0;
    defparam \b2v_inst.indice_2_LC_7_5_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.indice_2_LC_7_5_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \b2v_inst.indice_2_LC_7_5_1  (
            .in0(N__22107),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15087),
            .lcout(\b2v_inst.indiceZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34510),
            .ce(N__22033),
            .sr(N__38068));
    defparam \b2v_inst.indice_6_LC_7_5_4 .C_ON=1'b0;
    defparam \b2v_inst.indice_6_LC_7_5_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.indice_6_LC_7_5_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \b2v_inst.indice_6_LC_7_5_4  (
            .in0(_gnd_net_),
            .in1(N__22109),
            .in2(_gnd_net_),
            .in3(N__16215),
            .lcout(\b2v_inst.indiceZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34510),
            .ce(N__22033),
            .sr(N__38068));
    defparam \b2v_inst.indice_3_LC_7_5_6 .C_ON=1'b0;
    defparam \b2v_inst.indice_3_LC_7_5_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.indice_3_LC_7_5_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \b2v_inst.indice_3_LC_7_5_6  (
            .in0(_gnd_net_),
            .in1(N__22108),
            .in2(_gnd_net_),
            .in3(N__16071),
            .lcout(\b2v_inst.indiceZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34510),
            .ce(N__22033),
            .sr(N__38068));
    defparam \b2v_inst.un8_dir_mem_1_cry_0_c_LC_7_6_0 .C_ON=1'b1;
    defparam \b2v_inst.un8_dir_mem_1_cry_0_c_LC_7_6_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un8_dir_mem_1_cry_0_c_LC_7_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.un8_dir_mem_1_cry_0_c_LC_7_6_0  (
            .in0(_gnd_net_),
            .in1(N__39304),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_6_0_),
            .carryout(\b2v_inst.un8_dir_mem_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un8_dir_mem_1_cry_0_c_RNI4SNC_LC_7_6_1 .C_ON=1'b1;
    defparam \b2v_inst.un8_dir_mem_1_cry_0_c_RNI4SNC_LC_7_6_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un8_dir_mem_1_cry_0_c_RNI4SNC_LC_7_6_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst.un8_dir_mem_1_cry_0_c_RNI4SNC_LC_7_6_1  (
            .in0(_gnd_net_),
            .in1(N__38573),
            .in2(N__37288),
            .in3(N__14939),
            .lcout(\b2v_inst.un8_dir_mem_1_cry_0_c_RNI4SNCZ0 ),
            .ltout(),
            .carryin(\b2v_inst.un8_dir_mem_1_cry_0 ),
            .carryout(\b2v_inst.un8_dir_mem_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un8_dir_mem_1_cry_1_c_RNI6VOC_LC_7_6_2 .C_ON=1'b1;
    defparam \b2v_inst.un8_dir_mem_1_cry_1_c_RNI6VOC_LC_7_6_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un8_dir_mem_1_cry_1_c_RNI6VOC_LC_7_6_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.un8_dir_mem_1_cry_1_c_RNI6VOC_LC_7_6_2  (
            .in0(_gnd_net_),
            .in1(N__36050),
            .in2(_gnd_net_),
            .in3(N__14936),
            .lcout(\b2v_inst.un8_dir_mem_1_cry_1_c_RNI6VOCZ0 ),
            .ltout(),
            .carryin(\b2v_inst.un8_dir_mem_1_cry_1 ),
            .carryout(\b2v_inst.un8_dir_mem_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un8_dir_mem_1_cry_2_c_RNI82QC_LC_7_6_3 .C_ON=1'b1;
    defparam \b2v_inst.un8_dir_mem_1_cry_2_c_RNI82QC_LC_7_6_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un8_dir_mem_1_cry_2_c_RNI82QC_LC_7_6_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.un8_dir_mem_1_cry_2_c_RNI82QC_LC_7_6_3  (
            .in0(_gnd_net_),
            .in1(N__36499),
            .in2(_gnd_net_),
            .in3(N__14933),
            .lcout(\b2v_inst.un8_dir_mem_1_cry_2_c_RNI82QCZ0 ),
            .ltout(),
            .carryin(\b2v_inst.un8_dir_mem_1_cry_2 ),
            .carryout(\b2v_inst.un8_dir_mem_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un8_dir_mem_1_cry_3_c_RNIA5RC_LC_7_6_4 .C_ON=1'b1;
    defparam \b2v_inst.un8_dir_mem_1_cry_3_c_RNIA5RC_LC_7_6_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un8_dir_mem_1_cry_3_c_RNIA5RC_LC_7_6_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.un8_dir_mem_1_cry_3_c_RNIA5RC_LC_7_6_4  (
            .in0(_gnd_net_),
            .in1(N__36357),
            .in2(_gnd_net_),
            .in3(N__14930),
            .lcout(\b2v_inst.un8_dir_mem_1_cry_3_c_RNIA5RCZ0 ),
            .ltout(),
            .carryin(\b2v_inst.un8_dir_mem_1_cry_3 ),
            .carryout(\b2v_inst.un8_dir_mem_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un8_dir_mem_1_cry_4_c_RNIC8SC_LC_7_6_5 .C_ON=1'b1;
    defparam \b2v_inst.un8_dir_mem_1_cry_4_c_RNIC8SC_LC_7_6_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un8_dir_mem_1_cry_4_c_RNIC8SC_LC_7_6_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.un8_dir_mem_1_cry_4_c_RNIC8SC_LC_7_6_5  (
            .in0(_gnd_net_),
            .in1(N__35690),
            .in2(_gnd_net_),
            .in3(N__14966),
            .lcout(\b2v_inst.un8_dir_mem_1_cry_4_c_RNIC8SCZ0 ),
            .ltout(),
            .carryin(\b2v_inst.un8_dir_mem_1_cry_4 ),
            .carryout(\b2v_inst.un8_dir_mem_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un8_dir_mem_1_cry_5_c_RNIEBTC_LC_7_6_6 .C_ON=1'b1;
    defparam \b2v_inst.un8_dir_mem_1_cry_5_c_RNIEBTC_LC_7_6_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un8_dir_mem_1_cry_5_c_RNIEBTC_LC_7_6_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.un8_dir_mem_1_cry_5_c_RNIEBTC_LC_7_6_6  (
            .in0(_gnd_net_),
            .in1(N__38327),
            .in2(_gnd_net_),
            .in3(N__14963),
            .lcout(\b2v_inst.un8_dir_mem_1_cry_5_c_RNIEBTCZ0 ),
            .ltout(),
            .carryin(\b2v_inst.un8_dir_mem_1_cry_5 ),
            .carryout(\b2v_inst.un8_dir_mem_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un8_dir_mem_1_cry_6_c_RNIGEUC_LC_7_6_7 .C_ON=1'b1;
    defparam \b2v_inst.un8_dir_mem_1_cry_6_c_RNIGEUC_LC_7_6_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un8_dir_mem_1_cry_6_c_RNIGEUC_LC_7_6_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst.un8_dir_mem_1_cry_6_c_RNIGEUC_LC_7_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38860),
            .in3(N__14960),
            .lcout(\b2v_inst.dir_mem_115lto7 ),
            .ltout(),
            .carryin(\b2v_inst.un8_dir_mem_1_cry_6 ),
            .carryout(\b2v_inst.un8_dir_mem_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un8_dir_mem_1_cry_7_c_RNIIHVC_LC_7_7_0 .C_ON=1'b1;
    defparam \b2v_inst.un8_dir_mem_1_cry_7_c_RNIIHVC_LC_7_7_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un8_dir_mem_1_cry_7_c_RNIIHVC_LC_7_7_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.un8_dir_mem_1_cry_7_c_RNIIHVC_LC_7_7_0  (
            .in0(_gnd_net_),
            .in1(N__39080),
            .in2(_gnd_net_),
            .in3(N__14957),
            .lcout(\b2v_inst.un8_dir_mem_1_cry_7_c_RNIIHVCZ0 ),
            .ltout(),
            .carryin(bfn_7_7_0_),
            .carryout(\b2v_inst.un8_dir_mem_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un8_dir_mem_1_cry_8_c_RNIKK0D_LC_7_7_1 .C_ON=1'b1;
    defparam \b2v_inst.un8_dir_mem_1_cry_8_c_RNIKK0D_LC_7_7_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un8_dir_mem_1_cry_8_c_RNIKK0D_LC_7_7_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.un8_dir_mem_1_cry_8_c_RNIKK0D_LC_7_7_1  (
            .in0(_gnd_net_),
            .in1(N__35939),
            .in2(_gnd_net_),
            .in3(N__14954),
            .lcout(\b2v_inst.un8_dir_mem_1_cry_8_c_RNIKK0DZ0 ),
            .ltout(),
            .carryin(\b2v_inst.un8_dir_mem_1_cry_8 ),
            .carryout(\b2v_inst.un8_dir_mem_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un8_dir_mem_1_cry_9_c_RNITCOL_LC_7_7_2 .C_ON=1'b1;
    defparam \b2v_inst.un8_dir_mem_1_cry_9_c_RNITCOL_LC_7_7_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un8_dir_mem_1_cry_9_c_RNITCOL_LC_7_7_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.un8_dir_mem_1_cry_9_c_RNITCOL_LC_7_7_2  (
            .in0(_gnd_net_),
            .in1(N__36710),
            .in2(_gnd_net_),
            .in3(N__14951),
            .lcout(\b2v_inst.un8_dir_mem_1_cry_9_c_RNITCOLZ0 ),
            .ltout(),
            .carryin(\b2v_inst.un8_dir_mem_1_cry_9 ),
            .carryout(\b2v_inst.un8_dir_mem_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un8_dir_mem_1_cry_10_THRU_LUT4_0_LC_7_7_3 .C_ON=1'b0;
    defparam \b2v_inst.un8_dir_mem_1_cry_10_THRU_LUT4_0_LC_7_7_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un8_dir_mem_1_cry_10_THRU_LUT4_0_LC_7_7_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.un8_dir_mem_1_cry_10_THRU_LUT4_0_LC_7_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14948),
            .lcout(\b2v_inst.un8_dir_mem_1_cry_10_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un1_indice_cry_6_c_RNIRCFH4_LC_7_8_0 .C_ON=1'b0;
    defparam \b2v_inst.un1_indice_cry_6_c_RNIRCFH4_LC_7_8_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un1_indice_cry_6_c_RNIRCFH4_LC_7_8_0 .LUT_INIT=16'b1000100010000000;
    LogicCell40 \b2v_inst.un1_indice_cry_6_c_RNIRCFH4_LC_7_8_0  (
            .in0(N__20310),
            .in1(N__18796),
            .in2(N__18780),
            .in3(N__15098),
            .lcout(\b2v_inst.dir_mem_316lt11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un1_indice_cry_10_c_RNIO00U_LC_7_8_3 .C_ON=1'b0;
    defparam \b2v_inst.un1_indice_cry_10_c_RNIO00U_LC_7_8_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un1_indice_cry_10_c_RNIO00U_LC_7_8_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \b2v_inst.un1_indice_cry_10_c_RNIO00U_LC_7_8_3  (
            .in0(_gnd_net_),
            .in1(N__16150),
            .in2(_gnd_net_),
            .in3(N__20337),
            .lcout(\b2v_inst.dir_mem_316lto11_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_RNIJFGT1_0_LC_7_8_6 .C_ON=1'b0;
    defparam \b2v_inst.indice_RNIJFGT1_0_LC_7_8_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_RNIJFGT1_0_LC_7_8_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst.indice_RNIJFGT1_0_LC_7_8_6  (
            .in0(N__15088),
            .in1(N__16072),
            .in2(N__16250),
            .in3(N__18351),
            .lcout(),
            .ltout(\b2v_inst.dir_mem_316lt6_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un1_indice_cry_4_c_RNITUVU2_LC_7_8_7 .C_ON=1'b0;
    defparam \b2v_inst.un1_indice_cry_4_c_RNITUVU2_LC_7_8_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un1_indice_cry_4_c_RNITUVU2_LC_7_8_7 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \b2v_inst.un1_indice_cry_4_c_RNITUVU2_LC_7_8_7  (
            .in0(N__16216),
            .in1(_gnd_net_),
            .in2(N__15101),
            .in3(N__18834),
            .lcout(\b2v_inst.dir_mem_316lt7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_3_2_LC_7_9_0 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_3_2_LC_7_9_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.dir_mem_3_2_LC_7_9_0 .LUT_INIT=16'b1110111100100000;
    LogicCell40 \b2v_inst.dir_mem_3_2_LC_7_9_0  (
            .in0(N__15092),
            .in1(N__18262),
            .in2(N__18323),
            .in3(N__36092),
            .lcout(\b2v_inst.dir_mem_3Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34479),
            .ce(N__18208),
            .sr(_gnd_net_));
    defparam \b2v_inst.g0_0_i_a4_0_LC_7_10_3 .C_ON=1'b0;
    defparam \b2v_inst.g0_0_i_a4_0_LC_7_10_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.g0_0_i_a4_0_LC_7_10_3 .LUT_INIT=16'b1110000000000000;
    LogicCell40 \b2v_inst.g0_0_i_a4_0_LC_7_10_3  (
            .in0(N__15068),
            .in1(N__15062),
            .in2(N__15734),
            .in3(N__15681),
            .lcout(),
            .ltout(\b2v_inst.N_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.g0_0_i_2_LC_7_10_4 .C_ON=1'b0;
    defparam \b2v_inst.g0_0_i_2_LC_7_10_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.g0_0_i_2_LC_7_10_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \b2v_inst.g0_0_i_2_LC_7_10_4  (
            .in0(N__16430),
            .in1(N__16363),
            .in2(N__15053),
            .in3(N__16502),
            .lcout(\b2v_inst.g0_0_iZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un4_pix_count_intlto10_1_0_0_LC_7_11_0 .C_ON=1'b0;
    defparam \b2v_inst.un4_pix_count_intlto10_1_0_0_LC_7_11_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un4_pix_count_intlto10_1_0_0_LC_7_11_0 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \b2v_inst.un4_pix_count_intlto10_1_0_0_LC_7_11_0  (
            .in0(N__16424),
            .in1(N__16358),
            .in2(_gnd_net_),
            .in3(N__16494),
            .lcout(\b2v_inst.un4_pix_count_intlto10_1_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.g0_1_1_LC_7_11_1 .C_ON=1'b0;
    defparam \b2v_inst.g0_1_1_LC_7_11_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.g0_1_1_LC_7_11_1 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \b2v_inst.g0_1_1_LC_7_11_1  (
            .in0(N__15050),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15023),
            .lcout(\b2v_inst.g0_1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un4_pix_count_intlto15_1_a0_LC_7_11_3 .C_ON=1'b0;
    defparam \b2v_inst.un4_pix_count_intlto15_1_a0_LC_7_11_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un4_pix_count_intlto15_1_a0_LC_7_11_3 .LUT_INIT=16'b1000100010000000;
    LogicCell40 \b2v_inst.un4_pix_count_intlto15_1_a0_LC_7_11_3  (
            .in0(N__15344),
            .in1(N__15396),
            .in2(N__15546),
            .in3(N__15599),
            .lcout(\b2v_inst.un4_pix_count_intlto15_1_aZ0Z0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un4_pix_count_intlto6_1_ns_LC_7_11_4 .C_ON=1'b0;
    defparam \b2v_inst.un4_pix_count_intlto6_1_ns_LC_7_11_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un4_pix_count_intlto6_1_ns_LC_7_11_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \b2v_inst.un4_pix_count_intlto6_1_ns_LC_7_11_4  (
            .in0(N__15002),
            .in1(N__14993),
            .in2(_gnd_net_),
            .in3(N__14981),
            .lcout(),
            .ltout(\b2v_inst.un4_pix_count_intlt8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un4_pix_count_intlto10_1_0_LC_7_11_5 .C_ON=1'b0;
    defparam \b2v_inst.un4_pix_count_intlto10_1_0_LC_7_11_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un4_pix_count_intlto10_1_0_LC_7_11_5 .LUT_INIT=16'b0000000011001000;
    LogicCell40 \b2v_inst.un4_pix_count_intlto10_1_0_LC_7_11_5  (
            .in0(N__16266),
            .in1(N__15425),
            .in2(N__15419),
            .in3(N__15416),
            .lcout(\b2v_inst.un4_pix_count_intlt16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNO_25_29_LC_7_11_6 .C_ON=1'b0;
    defparam \b2v_inst.state_RNO_25_29_LC_7_11_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNO_25_29_LC_7_11_6 .LUT_INIT=16'b1000100010000000;
    LogicCell40 \b2v_inst.state_RNO_25_29_LC_7_11_6  (
            .in0(N__15397),
            .in1(N__15345),
            .in2(N__15778),
            .in3(N__15320),
            .lcout(\b2v_inst.state_RNO_25Z0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_RX_Byte_RNO_0_4_LC_7_12_0 .C_ON=1'b0;
    defparam \b2v_inst1.r_RX_Byte_RNO_0_4_LC_7_12_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_RX_Byte_RNO_0_4_LC_7_12_0 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \b2v_inst1.r_RX_Byte_RNO_0_4_LC_7_12_0  (
            .in0(N__17011),
            .in1(_gnd_net_),
            .in2(N__17060),
            .in3(N__16640),
            .lcout(),
            .ltout(\b2v_inst1.r_RX_Bytece_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_RX_Byte_4_LC_7_12_1 .C_ON=1'b0;
    defparam \b2v_inst1.r_RX_Byte_4_LC_7_12_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst1.r_RX_Byte_4_LC_7_12_1 .LUT_INIT=16'b1010110011001100;
    LogicCell40 \b2v_inst1.r_RX_Byte_4_LC_7_12_1  (
            .in0(N__22831),
            .in1(N__26773),
            .in2(N__15287),
            .in3(N__17285),
            .lcout(SYNTHESIZED_WIRE_10_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34469),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_SM_Main_RNIHNPV1_2_LC_7_12_2 .C_ON=1'b0;
    defparam \b2v_inst1.r_SM_Main_RNIHNPV1_2_LC_7_12_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_SM_Main_RNIHNPV1_2_LC_7_12_2 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \b2v_inst1.r_SM_Main_RNIHNPV1_2_LC_7_12_2  (
            .in0(N__16904),
            .in1(N__22627),
            .in2(N__22733),
            .in3(N__16536),
            .lcout(\b2v_inst1.N_47 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un4_pix_count_intlto10_1_d_0_x1_LC_7_12_3 .C_ON=1'b0;
    defparam \b2v_inst.un4_pix_count_intlto10_1_d_0_x1_LC_7_12_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un4_pix_count_intlto10_1_d_0_x1_LC_7_12_3 .LUT_INIT=16'b0000111100011111;
    LogicCell40 \b2v_inst.un4_pix_count_intlto10_1_d_0_x1_LC_7_12_3  (
            .in0(N__15529),
            .in1(N__15598),
            .in2(N__15682),
            .in3(N__15499),
            .lcout(),
            .ltout(\b2v_inst.un4_pix_count_intlto10_1_d_0_xZ0Z1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un4_pix_count_intlto10_1_d_0_ns_LC_7_12_4 .C_ON=1'b0;
    defparam \b2v_inst.un4_pix_count_intlto10_1_d_0_ns_LC_7_12_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un4_pix_count_intlto10_1_d_0_ns_LC_7_12_4 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \b2v_inst.un4_pix_count_intlto10_1_d_0_ns_LC_7_12_4  (
            .in0(N__37217),
            .in1(_gnd_net_),
            .in2(N__15284),
            .in3(N__15730),
            .lcout(\b2v_inst.un4_pix_count_intlto10_1_d_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_RX_Byte_RNO_0_6_LC_7_12_7 .C_ON=1'b0;
    defparam \b2v_inst1.r_RX_Byte_RNO_0_6_LC_7_12_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_RX_Byte_RNO_0_6_LC_7_12_7 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \b2v_inst1.r_RX_Byte_RNO_0_6_LC_7_12_7  (
            .in0(N__16639),
            .in1(N__17056),
            .in2(_gnd_net_),
            .in3(N__17010),
            .lcout(\b2v_inst1.r_RX_Bytece_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNO_24_29_LC_7_13_2 .C_ON=1'b0;
    defparam \b2v_inst.state_RNO_24_29_LC_7_13_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNO_24_29_LC_7_13_2 .LUT_INIT=16'b0011011111111111;
    LogicCell40 \b2v_inst.state_RNO_24_29_LC_7_13_2  (
            .in0(N__15280),
            .in1(N__15237),
            .in2(N__15200),
            .in3(N__15139),
            .lcout(),
            .ltout(\b2v_inst.un4_pix_count_intlto6_d_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNO_13_29_LC_7_13_3 .C_ON=1'b0;
    defparam \b2v_inst.state_RNO_13_29_LC_7_13_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNO_13_29_LC_7_13_3 .LUT_INIT=16'b0111011111110111;
    LogicCell40 \b2v_inst.state_RNO_13_29_LC_7_13_3  (
            .in0(N__15876),
            .in1(N__15826),
            .in2(N__15782),
            .in3(N__16744),
            .lcout(\b2v_inst.g2_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.g0_0_i_a4_0_1_LC_7_13_5 .C_ON=1'b0;
    defparam \b2v_inst.g0_0_i_a4_0_1_LC_7_13_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.g0_0_i_a4_0_1_LC_7_13_5 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \b2v_inst.g0_0_i_a4_0_1_LC_7_13_5  (
            .in0(N__15773),
            .in1(N__15547),
            .in2(N__15634),
            .in3(N__15500),
            .lcout(\b2v_inst.g0_0_i_a4Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un4_pix_count_intlto12_0_LC_7_13_6 .C_ON=1'b0;
    defparam \b2v_inst.un4_pix_count_intlto12_0_LC_7_13_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un4_pix_count_intlto12_0_LC_7_13_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \b2v_inst.un4_pix_count_intlto12_0_LC_7_13_6  (
            .in0(N__15729),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15683),
            .lcout(b2v_inst_un4_pix_count_intlto12_0),
            .ltout(b2v_inst_un4_pix_count_intlto12_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.g1_0_a4_0_1_LC_7_13_7 .C_ON=1'b0;
    defparam \b2v_inst.g1_0_a4_0_1_LC_7_13_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.g1_0_a4_0_1_LC_7_13_7 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \b2v_inst.g1_0_a4_0_1_LC_7_13_7  (
            .in0(N__15609),
            .in1(N__15548),
            .in2(N__15506),
            .in3(N__15501),
            .lcout(\b2v_inst.g1_0_a4Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_SM_Main_ns_2_0__m13_i_o2_LC_7_14_0 .C_ON=1'b0;
    defparam \b2v_inst1.r_SM_Main_ns_2_0__m13_i_o2_LC_7_14_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_SM_Main_ns_2_0__m13_i_o2_LC_7_14_0 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \b2v_inst1.r_SM_Main_ns_2_0__m13_i_o2_LC_7_14_0  (
            .in0(N__16632),
            .in1(N__17041),
            .in2(_gnd_net_),
            .in3(N__16995),
            .lcout(\b2v_inst1.N_49 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNIB55E1_6_LC_7_14_1 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNIB55E1_6_LC_7_14_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNIB55E1_6_LC_7_14_1 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \b2v_inst.data_a_escribir_RNIB55E1_6_LC_7_14_1  (
            .in0(N__37789),
            .in1(N__24740),
            .in2(N__35322),
            .in3(N__37496),
            .lcout(N_457_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_RX_Byte_RNO_1_0_LC_7_14_2 .C_ON=1'b0;
    defparam \b2v_inst1.r_RX_Byte_RNO_1_0_LC_7_14_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_RX_Byte_RNO_1_0_LC_7_14_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \b2v_inst1.r_RX_Byte_RNO_1_0_LC_7_14_2  (
            .in0(_gnd_net_),
            .in1(N__17042),
            .in2(_gnd_net_),
            .in3(N__16996),
            .lcout(\b2v_inst1.N_48 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_Bit_Index_RNIBK4I_1_LC_7_14_3 .C_ON=1'b0;
    defparam \b2v_inst1.r_Bit_Index_RNIBK4I_1_LC_7_14_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_Bit_Index_RNIBK4I_1_LC_7_14_3 .LUT_INIT=16'b0101111101011111;
    LogicCell40 \b2v_inst1.r_Bit_Index_RNIBK4I_1_LC_7_14_3  (
            .in0(N__16997),
            .in1(_gnd_net_),
            .in2(N__17055),
            .in3(_gnd_net_),
            .lcout(\b2v_inst1.N_44 ),
            .ltout(\b2v_inst1.N_44_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_Bit_Index_2_LC_7_14_4 .C_ON=1'b0;
    defparam \b2v_inst1.r_Bit_Index_2_LC_7_14_4 .SEQ_MODE=4'b1000;
    defparam \b2v_inst1.r_Bit_Index_2_LC_7_14_4 .LUT_INIT=16'b0000000011001001;
    LogicCell40 \b2v_inst1.r_Bit_Index_2_LC_7_14_4  (
            .in0(N__16003),
            .in1(N__16630),
            .in2(N__15428),
            .in3(N__16019),
            .lcout(\b2v_inst1.r_Bit_IndexZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34489),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.g1_0_0_2_LC_7_14_5 .C_ON=1'b0;
    defparam \b2v_inst.g1_0_0_2_LC_7_14_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.g1_0_0_2_LC_7_14_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \b2v_inst.g1_0_0_2_LC_7_14_5  (
            .in0(N__16423),
            .in1(N__16350),
            .in2(N__16034),
            .in3(N__16498),
            .lcout(\b2v_inst.g1_0_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_RX_Byte_0_LC_7_14_6 .C_ON=1'b0;
    defparam \b2v_inst1.r_RX_Byte_0_LC_7_14_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst1.r_RX_Byte_0_LC_7_14_6 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \b2v_inst1.r_RX_Byte_0_LC_7_14_6  (
            .in0(N__26712),
            .in1(N__17289),
            .in2(_gnd_net_),
            .in3(N__16025),
            .lcout(SYNTHESIZED_WIRE_10_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34489),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_Bit_Index_0_LC_7_14_7 .C_ON=1'b0;
    defparam \b2v_inst1.r_Bit_Index_0_LC_7_14_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst1.r_Bit_Index_0_LC_7_14_7 .LUT_INIT=16'b0010001000010001;
    LogicCell40 \b2v_inst1.r_Bit_Index_0_LC_7_14_7  (
            .in0(N__16998),
            .in1(N__16015),
            .in2(_gnd_net_),
            .in3(N__16002),
            .lcout(\b2v_inst1.r_Bit_IndexZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34489),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNI75II_29_LC_7_15_0 .C_ON=1'b0;
    defparam \b2v_inst.state_RNI75II_29_LC_7_15_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNI75II_29_LC_7_15_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst.state_RNI75II_29_LC_7_15_0  (
            .in0(_gnd_net_),
            .in1(N__28197),
            .in2(_gnd_net_),
            .in3(N__17714),
            .lcout(\b2v_inst.g3_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_SM_Main_RNIC98H_2_LC_7_15_1 .C_ON=1'b0;
    defparam \b2v_inst1.r_SM_Main_RNIC98H_2_LC_7_15_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_SM_Main_RNIC98H_2_LC_7_15_1 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \b2v_inst1.r_SM_Main_RNIC98H_2_LC_7_15_1  (
            .in0(N__22908),
            .in1(N__22720),
            .in2(_gnd_net_),
            .in3(N__22638),
            .lcout(\b2v_inst1.r_SM_Main_d_4 ),
            .ltout(\b2v_inst1.r_SM_Main_d_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_Bit_Index_1_LC_7_15_2 .C_ON=1'b0;
    defparam \b2v_inst1.r_Bit_Index_1_LC_7_15_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst1.r_Bit_Index_1_LC_7_15_2 .LUT_INIT=16'b0000100100001010;
    LogicCell40 \b2v_inst1.r_Bit_Index_1_LC_7_15_2  (
            .in0(N__17048),
            .in1(N__16004),
            .in2(N__15986),
            .in3(N__17012),
            .lcout(\b2v_inst1.r_Bit_IndexZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34500),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_RX_Byte_RNO_1_1_LC_7_15_3 .C_ON=1'b0;
    defparam \b2v_inst1.r_RX_Byte_RNO_1_1_LC_7_15_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_RX_Byte_RNO_1_1_LC_7_15_3 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \b2v_inst1.r_RX_Byte_RNO_1_1_LC_7_15_3  (
            .in0(_gnd_net_),
            .in1(N__17046),
            .in2(_gnd_net_),
            .in3(N__16999),
            .lcout(\b2v_inst1.N_51 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_RNIQGU15_9_LC_7_15_4 .C_ON=1'b0;
    defparam \b2v_inst.indice_RNIQGU15_9_LC_7_15_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_RNIQGU15_9_LC_7_15_4 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \b2v_inst.indice_RNIQGU15_9_LC_7_15_4  (
            .in0(N__16649),
            .in1(N__21654),
            .in2(N__35952),
            .in3(N__35216),
            .lcout(SYNTHESIZED_WIRE_12_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_RX_Byte_RNO_0_5_LC_7_15_7 .C_ON=1'b0;
    defparam \b2v_inst1.r_RX_Byte_RNO_0_5_LC_7_15_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_RX_Byte_RNO_0_5_LC_7_15_7 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \b2v_inst1.r_RX_Byte_RNO_0_5_LC_7_15_7  (
            .in0(N__16627),
            .in1(N__17047),
            .in2(_gnd_net_),
            .in3(N__17000),
            .lcout(\b2v_inst1.r_RX_Bytece_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_RNIJFHB_0_LC_8_5_0 .C_ON=1'b1;
    defparam \b2v_inst.indice_RNIJFHB_0_LC_8_5_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_RNIJFHB_0_LC_8_5_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst.indice_RNIJFHB_0_LC_8_5_0  (
            .in0(_gnd_net_),
            .in1(N__38574),
            .in2(_gnd_net_),
            .in3(N__39303),
            .lcout(\b2v_inst.indice_RNIJFHBZ0Z_0 ),
            .ltout(),
            .carryin(bfn_8_5_0_),
            .carryout(\b2v_inst.un2_dir_mem_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_RNILHHB_2_LC_8_5_1 .C_ON=1'b1;
    defparam \b2v_inst.indice_RNILHHB_2_LC_8_5_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_RNILHHB_2_LC_8_5_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.indice_RNILHHB_2_LC_8_5_1  (
            .in0(N__38575),
            .in1(N__36044),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst.indice_RNILHHBZ0Z_2 ),
            .ltout(),
            .carryin(\b2v_inst.un2_dir_mem_1_cry_0 ),
            .carryout(\b2v_inst.un2_dir_mem_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un2_dir_mem_1_cry_2_c_LC_8_5_2 .C_ON=1'b1;
    defparam \b2v_inst.un2_dir_mem_1_cry_2_c_LC_8_5_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un2_dir_mem_1_cry_2_c_LC_8_5_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.un2_dir_mem_1_cry_2_c_LC_8_5_2  (
            .in0(_gnd_net_),
            .in1(N__36527),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.un2_dir_mem_1_cry_1 ),
            .carryout(\b2v_inst.un2_dir_mem_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un2_dir_mem_1_cry_3_c_LC_8_5_3 .C_ON=1'b1;
    defparam \b2v_inst.un2_dir_mem_1_cry_3_c_LC_8_5_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un2_dir_mem_1_cry_3_c_LC_8_5_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.un2_dir_mem_1_cry_3_c_LC_8_5_3  (
            .in0(_gnd_net_),
            .in1(N__36337),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.un2_dir_mem_1_cry_2 ),
            .carryout(\b2v_inst.un2_dir_mem_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_1_RNO_0_5_LC_8_5_4 .C_ON=1'b1;
    defparam \b2v_inst.dir_mem_1_RNO_0_5_LC_8_5_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_1_RNO_0_5_LC_8_5_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst.dir_mem_1_RNO_0_5_LC_8_5_4  (
            .in0(_gnd_net_),
            .in1(N__35700),
            .in2(N__37158),
            .in3(N__16049),
            .lcout(\b2v_inst.dir_mem_1_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\b2v_inst.un2_dir_mem_1_cry_3 ),
            .carryout(\b2v_inst.un2_dir_mem_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_1_RNO_0_6_LC_8_5_5 .C_ON=1'b1;
    defparam \b2v_inst.dir_mem_1_RNO_0_6_LC_8_5_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_1_RNO_0_6_LC_8_5_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.dir_mem_1_RNO_0_6_LC_8_5_5  (
            .in0(_gnd_net_),
            .in1(N__38338),
            .in2(_gnd_net_),
            .in3(N__16046),
            .lcout(\b2v_inst.dir_mem_1_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\b2v_inst.un2_dir_mem_1_cry_4 ),
            .carryout(\b2v_inst.un2_dir_mem_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_1_RNO_0_7_LC_8_5_6 .C_ON=1'b1;
    defparam \b2v_inst.dir_mem_1_RNO_0_7_LC_8_5_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_1_RNO_0_7_LC_8_5_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst.dir_mem_1_RNO_0_7_LC_8_5_6  (
            .in0(_gnd_net_),
            .in1(N__38829),
            .in2(N__37159),
            .in3(N__16043),
            .lcout(\b2v_inst.dir_mem_1_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(\b2v_inst.un2_dir_mem_1_cry_5 ),
            .carryout(\b2v_inst.un2_dir_mem_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_1_RNO_0_8_LC_8_5_7 .C_ON=1'b1;
    defparam \b2v_inst.dir_mem_1_RNO_0_8_LC_8_5_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_1_RNO_0_8_LC_8_5_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.dir_mem_1_RNO_0_8_LC_8_5_7  (
            .in0(_gnd_net_),
            .in1(N__39068),
            .in2(_gnd_net_),
            .in3(N__16040),
            .lcout(\b2v_inst.dir_mem_1_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(\b2v_inst.un2_dir_mem_1_cry_6 ),
            .carryout(\b2v_inst.un2_dir_mem_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_1_RNO_0_9_LC_8_6_0 .C_ON=1'b1;
    defparam \b2v_inst.dir_mem_1_RNO_0_9_LC_8_6_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_1_RNO_0_9_LC_8_6_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.dir_mem_1_RNO_0_9_LC_8_6_0  (
            .in0(_gnd_net_),
            .in1(N__35920),
            .in2(_gnd_net_),
            .in3(N__16037),
            .lcout(\b2v_inst.dir_mem_1_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(bfn_8_6_0_),
            .carryout(\b2v_inst.un2_dir_mem_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_1_RNO_0_10_LC_8_6_1 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_1_RNO_0_10_LC_8_6_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_1_RNO_0_10_LC_8_6_1 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \b2v_inst.dir_mem_1_RNO_0_10_LC_8_6_1  (
            .in0(N__36728),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16163),
            .lcout(\b2v_inst.dir_mem_1_RNO_0Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un8_dir_mem_1_cry_1_c_RNIS26J1_LC_8_6_3 .C_ON=1'b0;
    defparam \b2v_inst.un8_dir_mem_1_cry_1_c_RNIS26J1_LC_8_6_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un8_dir_mem_1_cry_1_c_RNIS26J1_LC_8_6_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst.un8_dir_mem_1_cry_1_c_RNIS26J1_LC_8_6_3  (
            .in0(N__19123),
            .in1(N__18013),
            .in2(N__19275),
            .in3(N__17998),
            .lcout(\b2v_inst.dir_mem_115lt6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_RNIEPAH_4_LC_8_6_5 .C_ON=1'b0;
    defparam \b2v_inst.indice_RNIEPAH_4_LC_8_6_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_RNIEPAH_4_LC_8_6_5 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \b2v_inst.indice_RNIEPAH_4_LC_8_6_5  (
            .in0(N__35919),
            .in1(N__38313),
            .in2(_gnd_net_),
            .in3(N__36358),
            .lcout(\b2v_inst.indice_4_i_a2_0_7_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNI3UC9_11_LC_8_6_7 .C_ON=1'b0;
    defparam \b2v_inst.state_RNI3UC9_11_LC_8_6_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNI3UC9_11_LC_8_6_7 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \b2v_inst.state_RNI3UC9_11_LC_8_6_7  (
            .in0(N__25952),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26032),
            .lcout(\b2v_inst.N_442_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_3_0_LC_8_7_0 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_3_0_LC_8_7_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.dir_mem_3_0_LC_8_7_0 .LUT_INIT=16'b1111111000000001;
    LogicCell40 \b2v_inst.dir_mem_3_0_LC_8_7_0  (
            .in0(N__18254),
            .in1(N__20349),
            .in2(N__16160),
            .in3(N__39306),
            .lcout(\b2v_inst.dir_mem_3Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34490),
            .ce(N__18209),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_3_10_LC_8_7_1 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_3_10_LC_8_7_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.dir_mem_3_10_LC_8_7_1 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \b2v_inst.dir_mem_3_10_LC_8_7_1  (
            .in0(N__20350),
            .in1(N__16159),
            .in2(N__16139),
            .in3(N__18255),
            .lcout(\b2v_inst.dir_mem_3Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34490),
            .ce(N__18209),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_3_7_LC_8_7_3 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_3_7_LC_8_7_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.dir_mem_3_7_LC_8_7_3 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \b2v_inst.dir_mem_3_7_LC_8_7_3  (
            .in0(N__18784),
            .in1(N__18313),
            .in2(N__16121),
            .in3(N__18253),
            .lcout(\b2v_inst.dir_mem_3Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34490),
            .ce(N__18209),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_3_8_LC_8_7_4 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_3_8_LC_8_7_4 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.dir_mem_3_8_LC_8_7_4 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \b2v_inst.dir_mem_3_8_LC_8_7_4  (
            .in0(N__18258),
            .in1(N__20320),
            .in2(N__16106),
            .in3(N__18318),
            .lcout(\b2v_inst.dir_mem_3Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34490),
            .ce(N__18209),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_3_9_LC_8_7_5 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_3_9_LC_8_7_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.dir_mem_3_9_LC_8_7_5 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \b2v_inst.dir_mem_3_9_LC_8_7_5  (
            .in0(N__18808),
            .in1(N__18314),
            .in2(N__16091),
            .in3(N__18259),
            .lcout(\b2v_inst.dir_mem_3Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34490),
            .ce(N__18209),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_3_3_LC_8_7_6 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_3_3_LC_8_7_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.dir_mem_3_3_LC_8_7_6 .LUT_INIT=16'b1110111101000000;
    LogicCell40 \b2v_inst.dir_mem_3_3_LC_8_7_6  (
            .in0(N__18256),
            .in1(N__16076),
            .in2(N__18324),
            .in3(N__36565),
            .lcout(\b2v_inst.dir_mem_3Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34490),
            .ce(N__18209),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_3_5_LC_8_7_7 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_3_5_LC_8_7_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.dir_mem_3_5_LC_8_7_7 .LUT_INIT=16'b0101010111000101;
    LogicCell40 \b2v_inst.dir_mem_3_5_LC_8_7_7  (
            .in0(N__35705),
            .in1(N__18841),
            .in2(N__18325),
            .in3(N__18257),
            .lcout(\b2v_inst.dir_mem_3Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34490),
            .ce(N__18209),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_3_1_LC_8_8_2 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_3_1_LC_8_8_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.dir_mem_3_1_LC_8_8_2 .LUT_INIT=16'b1110111100100000;
    LogicCell40 \b2v_inst.dir_mem_3_1_LC_8_8_2  (
            .in0(N__16246),
            .in1(N__18260),
            .in2(N__18322),
            .in3(N__38640),
            .lcout(\b2v_inst.dir_mem_3Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34480),
            .ce(N__18204),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_3_6_LC_8_8_4 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_3_6_LC_8_8_4 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.dir_mem_3_6_LC_8_8_4 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \b2v_inst.dir_mem_3_6_LC_8_8_4  (
            .in0(N__18306),
            .in1(N__16220),
            .in2(N__16193),
            .in3(N__18261),
            .lcout(\b2v_inst.dir_mem_3Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34480),
            .ce(N__18204),
            .sr(_gnd_net_));
    defparam \b2v_inst.un3_dir_mem_cry_0_c_LC_8_9_0 .C_ON=1'b1;
    defparam \b2v_inst.un3_dir_mem_cry_0_c_LC_8_9_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un3_dir_mem_cry_0_c_LC_8_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.un3_dir_mem_cry_0_c_LC_8_9_0  (
            .in0(_gnd_net_),
            .in1(N__39305),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_9_0_),
            .carryout(\b2v_inst.un3_dir_mem_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un3_dir_mem_cry_1_c_LC_8_9_1 .C_ON=1'b1;
    defparam \b2v_inst.un3_dir_mem_cry_1_c_LC_8_9_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un3_dir_mem_cry_1_c_LC_8_9_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.un3_dir_mem_cry_1_c_LC_8_9_1  (
            .in0(_gnd_net_),
            .in1(N__38642),
            .in2(N__37157),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.un3_dir_mem_cry_0 ),
            .carryout(\b2v_inst.un3_dir_mem_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_2_LC_8_9_2 .C_ON=1'b1;
    defparam \b2v_inst.dir_mem_2_LC_8_9_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.dir_mem_2_LC_8_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst.dir_mem_2_LC_8_9_2  (
            .in0(_gnd_net_),
            .in1(N__36103),
            .in2(N__37152),
            .in3(N__16175),
            .lcout(\b2v_inst.dir_memZ0Z_2 ),
            .ltout(),
            .carryin(\b2v_inst.un3_dir_mem_cry_1 ),
            .carryout(\b2v_inst.un3_dir_mem_cry_2 ),
            .clk(N__34470),
            .ce(N__22170),
            .sr(N__38061));
    defparam \b2v_inst.dir_mem_3_LC_8_9_3 .C_ON=1'b1;
    defparam \b2v_inst.dir_mem_3_LC_8_9_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.dir_mem_3_LC_8_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst.dir_mem_3_LC_8_9_3  (
            .in0(_gnd_net_),
            .in1(N__36570),
            .in2(N__37155),
            .in3(N__16172),
            .lcout(\b2v_inst.dir_memZ0Z_3 ),
            .ltout(),
            .carryin(\b2v_inst.un3_dir_mem_cry_2 ),
            .carryout(\b2v_inst.un3_dir_mem_cry_3 ),
            .clk(N__34470),
            .ce(N__22170),
            .sr(N__38061));
    defparam \b2v_inst.dir_mem_4_LC_8_9_4 .C_ON=1'b1;
    defparam \b2v_inst.dir_mem_4_LC_8_9_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.dir_mem_4_LC_8_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst.dir_mem_4_LC_8_9_4  (
            .in0(_gnd_net_),
            .in1(N__36359),
            .in2(N__37153),
            .in3(N__16169),
            .lcout(\b2v_inst.dir_memZ0Z_4 ),
            .ltout(),
            .carryin(\b2v_inst.un3_dir_mem_cry_3 ),
            .carryout(\b2v_inst.un3_dir_mem_cry_4 ),
            .clk(N__34470),
            .ce(N__22170),
            .sr(N__38061));
    defparam \b2v_inst.dir_mem_RNO_0_5_LC_8_9_5 .C_ON=1'b1;
    defparam \b2v_inst.dir_mem_RNO_0_5_LC_8_9_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNO_0_5_LC_8_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst.dir_mem_RNO_0_5_LC_8_9_5  (
            .in0(_gnd_net_),
            .in1(N__37063),
            .in2(N__35715),
            .in3(N__16166),
            .lcout(\b2v_inst.dir_mem_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\b2v_inst.un3_dir_mem_cry_4 ),
            .carryout(\b2v_inst.un3_dir_mem_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_RNO_0_6_LC_8_9_6 .C_ON=1'b1;
    defparam \b2v_inst.dir_mem_RNO_0_6_LC_8_9_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNO_0_6_LC_8_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst.dir_mem_RNO_0_6_LC_8_9_6  (
            .in0(_gnd_net_),
            .in1(N__38359),
            .in2(N__37154),
            .in3(N__16517),
            .lcout(\b2v_inst.dir_mem_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\b2v_inst.un3_dir_mem_cry_5 ),
            .carryout(\b2v_inst.un3_dir_mem_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_7_LC_8_9_7 .C_ON=1'b1;
    defparam \b2v_inst.dir_mem_7_LC_8_9_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.dir_mem_7_LC_8_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst.dir_mem_7_LC_8_9_7  (
            .in0(_gnd_net_),
            .in1(N__38847),
            .in2(N__37156),
            .in3(N__16514),
            .lcout(\b2v_inst.dir_memZ0Z_7 ),
            .ltout(),
            .carryin(\b2v_inst.un3_dir_mem_cry_6 ),
            .carryout(\b2v_inst.un3_dir_mem_cry_7 ),
            .clk(N__34470),
            .ce(N__22170),
            .sr(N__38061));
    defparam \b2v_inst.dir_mem_RNO_0_8_LC_8_10_0 .C_ON=1'b1;
    defparam \b2v_inst.dir_mem_RNO_0_8_LC_8_10_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNO_0_8_LC_8_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst.dir_mem_RNO_0_8_LC_8_10_0  (
            .in0(_gnd_net_),
            .in1(N__39069),
            .in2(N__37151),
            .in3(N__16511),
            .lcout(\b2v_inst.dir_mem_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(bfn_8_10_0_),
            .carryout(\b2v_inst.un3_dir_mem_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_RNO_0_9_LC_8_10_1 .C_ON=1'b1;
    defparam \b2v_inst.dir_mem_RNO_0_9_LC_8_10_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNO_0_9_LC_8_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst.dir_mem_RNO_0_9_LC_8_10_1  (
            .in0(_gnd_net_),
            .in1(N__37056),
            .in2(N__35954),
            .in3(N__16508),
            .lcout(\b2v_inst.dir_mem_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(\b2v_inst.un3_dir_mem_cry_8 ),
            .carryout(\b2v_inst.un3_dir_mem_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_10_LC_8_10_2 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_10_LC_8_10_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.dir_mem_10_LC_8_10_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \b2v_inst.dir_mem_10_LC_8_10_2  (
            .in0(_gnd_net_),
            .in1(N__36745),
            .in2(_gnd_net_),
            .in3(N__16505),
            .lcout(\b2v_inst.dir_memZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34458),
            .ce(N__22187),
            .sr(N__38056));
    defparam \b2v_inst.state_RNO_14_29_LC_8_11_0 .C_ON=1'b0;
    defparam \b2v_inst.state_RNO_14_29_LC_8_11_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNO_14_29_LC_8_11_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst.state_RNO_14_29_LC_8_11_0  (
            .in0(N__16501),
            .in1(N__16425),
            .in2(N__16364),
            .in3(N__16289),
            .lcout(),
            .ltout(\b2v_inst.m29_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNO_5_29_LC_8_11_1 .C_ON=1'b0;
    defparam \b2v_inst.state_RNO_5_29_LC_8_11_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNO_5_29_LC_8_11_1 .LUT_INIT=16'b1111000001000000;
    LogicCell40 \b2v_inst.state_RNO_5_29_LC_8_11_1  (
            .in0(N__16853),
            .in1(N__16283),
            .in2(N__16274),
            .in3(N__16267),
            .lcout(\b2v_inst.o2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_Clk_Count_RNI64771_0_LC_8_11_2 .C_ON=1'b0;
    defparam \b2v_inst1.r_Clk_Count_RNI64771_0_LC_8_11_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_Clk_Count_RNI64771_0_LC_8_11_2 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \b2v_inst1.r_Clk_Count_RNI64771_0_LC_8_11_2  (
            .in0(N__16905),
            .in1(N__21077),
            .in2(_gnd_net_),
            .in3(N__21108),
            .lcout(\b2v_inst1.un22_r_clk_count_ac0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNO_20_29_LC_8_11_5 .C_ON=1'b0;
    defparam \b2v_inst.state_RNO_20_29_LC_8_11_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNO_20_29_LC_8_11_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst.state_RNO_20_29_LC_8_11_5  (
            .in0(N__25686),
            .in1(N__26075),
            .in2(N__25742),
            .in3(N__25439),
            .lcout(\b2v_inst.N_618_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_Clk_Count_RNI4O4Q_0_LC_8_11_7 .C_ON=1'b0;
    defparam \b2v_inst1.r_Clk_Count_RNI4O4Q_0_LC_8_11_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_Clk_Count_RNI4O4Q_0_LC_8_11_7 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \b2v_inst1.r_Clk_Count_RNI4O4Q_0_LC_8_11_7  (
            .in0(N__21109),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16906),
            .lcout(\b2v_inst1.N_119 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNO_22_29_LC_8_12_0 .C_ON=1'b0;
    defparam \b2v_inst.state_RNO_22_29_LC_8_12_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNO_22_29_LC_8_12_0 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \b2v_inst.state_RNO_22_29_LC_8_12_0  (
            .in0(N__30875),
            .in1(N__24658),
            .in2(N__28201),
            .in3(N__25827),
            .lcout(\b2v_inst.G_40_i_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_SM_Main_ns_2_0__m13_i_a3_2_LC_8_12_4 .C_ON=1'b0;
    defparam \b2v_inst1.r_SM_Main_ns_2_0__m13_i_a3_2_LC_8_12_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_SM_Main_ns_2_0__m13_i_a3_2_LC_8_12_4 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \b2v_inst1.r_SM_Main_ns_2_0__m13_i_a3_2_LC_8_12_4  (
            .in0(N__22643),
            .in1(N__21181),
            .in2(N__22924),
            .in3(N__21082),
            .lcout(\b2v_inst1.N_96 ),
            .ltout(\b2v_inst1.N_96_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_Clk_Count_0_LC_8_12_5 .C_ON=1'b0;
    defparam \b2v_inst1.r_Clk_Count_0_LC_8_12_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst1.r_Clk_Count_0_LC_8_12_5 .LUT_INIT=16'b0000001000001100;
    LogicCell40 \b2v_inst1.r_Clk_Count_0_LC_8_12_5  (
            .in0(N__22724),
            .in1(N__21150),
            .in2(N__16577),
            .in3(N__21112),
            .lcout(\b2v_inst1.r_Clk_CountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34459),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.g0_0_i_LC_8_12_6 .C_ON=1'b0;
    defparam \b2v_inst.g0_0_i_LC_8_12_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.g0_0_i_LC_8_12_6 .LUT_INIT=16'b1110111011001110;
    LogicCell40 \b2v_inst.g0_0_i_LC_8_12_6  (
            .in0(N__16574),
            .in1(N__16568),
            .in2(N__16559),
            .in3(N__16848),
            .lcout(\b2v_inst.N_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_Clk_Count_RNO_0_2_LC_8_13_0 .C_ON=1'b0;
    defparam \b2v_inst1.r_Clk_Count_RNO_0_2_LC_8_13_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_Clk_Count_RNO_0_2_LC_8_13_0 .LUT_INIT=16'b1001001100110011;
    LogicCell40 \b2v_inst1.r_Clk_Count_RNO_0_2_LC_8_13_0  (
            .in0(N__21111),
            .in1(N__16902),
            .in2(N__21083),
            .in3(N__21145),
            .lcout(),
            .ltout(\b2v_inst1.N_58_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_Clk_Count_2_LC_8_13_1 .C_ON=1'b0;
    defparam \b2v_inst1.r_Clk_Count_2_LC_8_13_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst1.r_Clk_Count_2_LC_8_13_1 .LUT_INIT=16'b0000111100001010;
    LogicCell40 \b2v_inst1.r_Clk_Count_2_LC_8_13_1  (
            .in0(N__21146),
            .in1(_gnd_net_),
            .in2(N__16544),
            .in3(N__22713),
            .lcout(\b2v_inst1.r_Clk_CountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34471),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_SM_Main_2_LC_8_13_2 .C_ON=1'b0;
    defparam \b2v_inst1.r_SM_Main_2_LC_8_13_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst1.r_SM_Main_2_LC_8_13_2 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \b2v_inst1.r_SM_Main_2_LC_8_13_2  (
            .in0(N__22626),
            .in1(N__20902),
            .in2(_gnd_net_),
            .in3(N__22916),
            .lcout(\b2v_inst1.r_SM_MainZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34471),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_Clk_Count_RNIGMPV1_2_LC_8_13_3 .C_ON=1'b0;
    defparam \b2v_inst1.r_Clk_Count_RNIGMPV1_2_LC_8_13_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_Clk_Count_RNIGMPV1_2_LC_8_13_3 .LUT_INIT=16'b1010110011111100;
    LogicCell40 \b2v_inst1.r_Clk_Count_RNIGMPV1_2_LC_8_13_3  (
            .in0(N__16540),
            .in1(N__22624),
            .in2(N__22923),
            .in3(N__16903),
            .lcout(\b2v_inst1.N_43 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_RX_Byte_6_LC_8_13_4 .C_ON=1'b0;
    defparam \b2v_inst1.r_RX_Byte_6_LC_8_13_4 .SEQ_MODE=4'b1000;
    defparam \b2v_inst1.r_RX_Byte_6_LC_8_13_4 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \b2v_inst1.r_RX_Byte_6_LC_8_13_4  (
            .in0(N__16919),
            .in1(N__22830),
            .in2(N__26761),
            .in3(N__17290),
            .lcout(SYNTHESIZED_WIRE_10_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34471),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_SM_Main_ns_2_0__m16_0_o2_LC_8_13_5 .C_ON=1'b0;
    defparam \b2v_inst1.r_SM_Main_ns_2_0__m16_0_o2_LC_8_13_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_SM_Main_ns_2_0__m16_0_o2_LC_8_13_5 .LUT_INIT=16'b0101010101110111;
    LogicCell40 \b2v_inst1.r_SM_Main_ns_2_0__m16_0_o2_LC_8_13_5  (
            .in0(N__16901),
            .in1(N__21078),
            .in2(_gnd_net_),
            .in3(N__21110),
            .lcout(\b2v_inst1.m16_0_o2 ),
            .ltout(\b2v_inst1.m16_0_o2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_SM_Main_ns_2_0__m13_i_2_LC_8_13_6 .C_ON=1'b0;
    defparam \b2v_inst1.r_SM_Main_ns_2_0__m13_i_2_LC_8_13_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_SM_Main_ns_2_0__m13_i_2_LC_8_13_6 .LUT_INIT=16'b0100110001001000;
    LogicCell40 \b2v_inst1.r_SM_Main_ns_2_0__m13_i_2_LC_8_13_6  (
            .in0(N__22625),
            .in1(N__22915),
            .in2(N__16865),
            .in3(N__17314),
            .lcout(\b2v_inst1.m13_i_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.g1_LC_8_13_7 .C_ON=1'b0;
    defparam \b2v_inst.g1_LC_8_13_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.g1_LC_8_13_7 .LUT_INIT=16'b0010001000110010;
    LogicCell40 \b2v_inst.g1_LC_8_13_7  (
            .in0(N__16862),
            .in1(N__16842),
            .in2(N__16775),
            .in3(N__16745),
            .lcout(\b2v_inst.g1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.g0_1_LC_8_14_1 .C_ON=1'b0;
    defparam \b2v_inst.g0_1_LC_8_14_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.g0_1_LC_8_14_1 .LUT_INIT=16'b1101110000000000;
    LogicCell40 \b2v_inst.g0_1_LC_8_14_1  (
            .in0(N__16688),
            .in1(N__16682),
            .in2(N__16676),
            .in3(N__17611),
            .lcout(\b2v_inst.g3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_energia_RNID0NB2_9_LC_8_14_2 .C_ON=1'b0;
    defparam \b2v_inst.dir_energia_RNID0NB2_9_LC_8_14_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_energia_RNID0NB2_9_LC_8_14_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst.dir_energia_RNID0NB2_9_LC_8_14_2  (
            .in0(N__16667),
            .in1(N__21718),
            .in2(_gnd_net_),
            .in3(N__35819),
            .lcout(\b2v_inst.addr_ram_energia_m0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_RX_Byte_RNO_0_2_LC_8_14_4 .C_ON=1'b0;
    defparam \b2v_inst1.r_RX_Byte_RNO_0_2_LC_8_14_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_RX_Byte_RNO_0_2_LC_8_14_4 .LUT_INIT=16'b0000111000011111;
    LogicCell40 \b2v_inst1.r_RX_Byte_RNO_0_2_LC_8_14_4  (
            .in0(N__16964),
            .in1(N__16631),
            .in2(N__26986),
            .in3(N__22826),
            .lcout(),
            .ltout(\b2v_inst1.N_38_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_RX_Byte_2_LC_8_14_5 .C_ON=1'b0;
    defparam \b2v_inst1.r_RX_Byte_2_LC_8_14_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst1.r_RX_Byte_2_LC_8_14_5 .LUT_INIT=16'b0101111100001010;
    LogicCell40 \b2v_inst1.r_RX_Byte_2_LC_8_14_5  (
            .in0(N__17302),
            .in1(_gnd_net_),
            .in2(N__16643),
            .in3(N__26982),
            .lcout(SYNTHESIZED_WIRE_10_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34481),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_RX_Byte_RNO_0_3_LC_8_14_6 .C_ON=1'b0;
    defparam \b2v_inst1.r_RX_Byte_RNO_0_3_LC_8_14_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_RX_Byte_RNO_0_3_LC_8_14_6 .LUT_INIT=16'b0000111100011011;
    LogicCell40 \b2v_inst1.r_RX_Byte_RNO_0_3_LC_8_14_6  (
            .in0(N__16629),
            .in1(N__22827),
            .in2(N__26800),
            .in3(N__16583),
            .lcout(),
            .ltout(\b2v_inst1.N_36_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_RX_Byte_3_LC_8_14_7 .C_ON=1'b0;
    defparam \b2v_inst1.r_RX_Byte_3_LC_8_14_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst1.r_RX_Byte_3_LC_8_14_7 .LUT_INIT=16'b0101111100001010;
    LogicCell40 \b2v_inst1.r_RX_Byte_3_LC_8_14_7  (
            .in0(N__17303),
            .in1(_gnd_net_),
            .in2(N__17063),
            .in3(N__26796),
            .lcout(SYNTHESIZED_WIRE_10_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34481),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_RX_Byte_RNO_1_2_LC_8_15_1 .C_ON=1'b0;
    defparam \b2v_inst1.r_RX_Byte_RNO_1_2_LC_8_15_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_RX_Byte_RNO_1_2_LC_8_15_1 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \b2v_inst1.r_RX_Byte_RNO_1_2_LC_8_15_1  (
            .in0(_gnd_net_),
            .in1(N__17054),
            .in2(_gnd_net_),
            .in3(N__17009),
            .lcout(\b2v_inst1.N_50 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_RX_Byte_5_LC_8_15_5 .C_ON=1'b0;
    defparam \b2v_inst1.r_RX_Byte_5_LC_8_15_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst1.r_RX_Byte_5_LC_8_15_5 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \b2v_inst1.r_RX_Byte_5_LC_8_15_5  (
            .in0(N__17300),
            .in1(N__28813),
            .in2(N__16958),
            .in3(N__22816),
            .lcout(SYNTHESIZED_WIRE_10_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34491),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNIAD041_9_LC_8_15_6 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNIAD041_9_LC_8_15_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNIAD041_9_LC_8_15_6 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \b2v_inst.data_a_escribir_RNIAD041_9_LC_8_15_6  (
            .in0(N__37467),
            .in1(N__37791),
            .in2(N__32872),
            .in3(N__24677),
            .lcout(N_460_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNI79V31_8_LC_8_15_7 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNI79V31_8_LC_8_15_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNI79V31_8_LC_8_15_7 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \b2v_inst.data_a_escribir_RNI79V31_8_LC_8_15_7  (
            .in0(N__37790),
            .in1(N__24692),
            .in2(N__33398),
            .in3(N__37466),
            .lcout(N_459_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un8_dir_mem_2_cry_1_c_LC_9_5_0 .C_ON=1'b1;
    defparam \b2v_inst.un8_dir_mem_2_cry_1_c_LC_9_5_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un8_dir_mem_2_cry_1_c_LC_9_5_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.un8_dir_mem_2_cry_1_c_LC_9_5_0  (
            .in0(_gnd_net_),
            .in1(N__38587),
            .in2(N__36076),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_5_0_),
            .carryout(\b2v_inst.un8_dir_mem_2_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un8_dir_mem_2_cry_1_c_RNI88LL_LC_9_5_1 .C_ON=1'b1;
    defparam \b2v_inst.un8_dir_mem_2_cry_1_c_RNI88LL_LC_9_5_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un8_dir_mem_2_cry_1_c_RNI88LL_LC_9_5_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.un8_dir_mem_2_cry_1_c_RNI88LL_LC_9_5_1  (
            .in0(_gnd_net_),
            .in1(N__36523),
            .in2(_gnd_net_),
            .in3(N__16928),
            .lcout(\b2v_inst.un8_dir_mem_2_cry_1_c_RNI88LLZ0 ),
            .ltout(),
            .carryin(\b2v_inst.un8_dir_mem_2_cry_1 ),
            .carryout(\b2v_inst.un8_dir_mem_2_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un8_dir_mem_2_cry_2_c_RNIABML_LC_9_5_2 .C_ON=1'b1;
    defparam \b2v_inst.un8_dir_mem_2_cry_2_c_RNIABML_LC_9_5_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un8_dir_mem_2_cry_2_c_RNIABML_LC_9_5_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.un8_dir_mem_2_cry_2_c_RNIABML_LC_9_5_2  (
            .in0(_gnd_net_),
            .in1(N__36309),
            .in2(_gnd_net_),
            .in3(N__16925),
            .lcout(\b2v_inst.un8_dir_mem_2_cry_2_c_RNIABMLZ0 ),
            .ltout(),
            .carryin(\b2v_inst.un8_dir_mem_2_cry_2 ),
            .carryout(\b2v_inst.un8_dir_mem_2_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un8_dir_mem_2_cry_3_c_RNICENL_LC_9_5_3 .C_ON=1'b1;
    defparam \b2v_inst.un8_dir_mem_2_cry_3_c_RNICENL_LC_9_5_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un8_dir_mem_2_cry_3_c_RNICENL_LC_9_5_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.un8_dir_mem_2_cry_3_c_RNICENL_LC_9_5_3  (
            .in0(_gnd_net_),
            .in1(N__35669),
            .in2(_gnd_net_),
            .in3(N__16922),
            .lcout(\b2v_inst.un8_dir_mem_2_cry_3_c_RNICENLZ0 ),
            .ltout(),
            .carryin(\b2v_inst.un8_dir_mem_2_cry_3 ),
            .carryout(\b2v_inst.un8_dir_mem_2_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un8_dir_mem_2_cry_4_c_RNIEHOL_LC_9_5_4 .C_ON=1'b1;
    defparam \b2v_inst.un8_dir_mem_2_cry_4_c_RNIEHOL_LC_9_5_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un8_dir_mem_2_cry_4_c_RNIEHOL_LC_9_5_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.un8_dir_mem_2_cry_4_c_RNIEHOL_LC_9_5_4  (
            .in0(_gnd_net_),
            .in1(N__38342),
            .in2(_gnd_net_),
            .in3(N__17087),
            .lcout(\b2v_inst.un8_dir_mem_2_cry_4_c_RNIEHOLZ0 ),
            .ltout(),
            .carryin(\b2v_inst.un8_dir_mem_2_cry_4 ),
            .carryout(\b2v_inst.un8_dir_mem_2_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un8_dir_mem_2_cry_5_c_RNIGKP5_LC_9_5_5 .C_ON=1'b1;
    defparam \b2v_inst.un8_dir_mem_2_cry_5_c_RNIGKP5_LC_9_5_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un8_dir_mem_2_cry_5_c_RNIGKP5_LC_9_5_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.un8_dir_mem_2_cry_5_c_RNIGKP5_LC_9_5_5  (
            .in0(_gnd_net_),
            .in1(N__38828),
            .in2(_gnd_net_),
            .in3(N__17084),
            .lcout(\b2v_inst.dir_mem_215lto7 ),
            .ltout(),
            .carryin(\b2v_inst.un8_dir_mem_2_cry_5 ),
            .carryout(\b2v_inst.un8_dir_mem_2_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un8_dir_mem_2_cry_6_c_RNIINQ5_LC_9_5_6 .C_ON=1'b1;
    defparam \b2v_inst.un8_dir_mem_2_cry_6_c_RNIINQ5_LC_9_5_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un8_dir_mem_2_cry_6_c_RNIINQ5_LC_9_5_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.un8_dir_mem_2_cry_6_c_RNIINQ5_LC_9_5_6  (
            .in0(_gnd_net_),
            .in1(N__39034),
            .in2(_gnd_net_),
            .in3(N__17081),
            .lcout(\b2v_inst.un8_dir_mem_2_cry_6_c_RNIINQZ0Z5 ),
            .ltout(),
            .carryin(\b2v_inst.un8_dir_mem_2_cry_6 ),
            .carryout(\b2v_inst.un8_dir_mem_2_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un8_dir_mem_2_cry_7_c_RNIKQR5_LC_9_5_7 .C_ON=1'b1;
    defparam \b2v_inst.un8_dir_mem_2_cry_7_c_RNIKQR5_LC_9_5_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un8_dir_mem_2_cry_7_c_RNIKQR5_LC_9_5_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.un8_dir_mem_2_cry_7_c_RNIKQR5_LC_9_5_7  (
            .in0(_gnd_net_),
            .in1(N__35911),
            .in2(_gnd_net_),
            .in3(N__17078),
            .lcout(\b2v_inst.un8_dir_mem_2_cry_7_c_RNIKQRZ0Z5 ),
            .ltout(),
            .carryin(\b2v_inst.un8_dir_mem_2_cry_7 ),
            .carryout(\b2v_inst.un8_dir_mem_2_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un8_dir_mem_2_cry_8_c_RNITIJE_LC_9_6_0 .C_ON=1'b1;
    defparam \b2v_inst.un8_dir_mem_2_cry_8_c_RNITIJE_LC_9_6_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un8_dir_mem_2_cry_8_c_RNITIJE_LC_9_6_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.un8_dir_mem_2_cry_8_c_RNITIJE_LC_9_6_0  (
            .in0(_gnd_net_),
            .in1(N__36727),
            .in2(_gnd_net_),
            .in3(N__17075),
            .lcout(\b2v_inst.un8_dir_mem_2_cry_8_c_RNITIJEZ0 ),
            .ltout(),
            .carryin(bfn_9_6_0_),
            .carryout(\b2v_inst.un8_dir_mem_2_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un8_dir_mem_2_cry_9_THRU_LUT4_0_LC_9_6_1 .C_ON=1'b0;
    defparam \b2v_inst.un8_dir_mem_2_cry_9_THRU_LUT4_0_LC_9_6_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un8_dir_mem_2_cry_9_THRU_LUT4_0_LC_9_6_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.un8_dir_mem_2_cry_9_THRU_LUT4_0_LC_9_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17072),
            .lcout(\b2v_inst.un8_dir_mem_2_cry_9_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_RNIHTLS1_1_LC_9_6_2 .C_ON=1'b0;
    defparam \b2v_inst.indice_RNIHTLS1_1_LC_9_6_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_RNIHTLS1_1_LC_9_6_2 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \b2v_inst.indice_RNIHTLS1_1_LC_9_6_2  (
            .in0(N__19059),
            .in1(N__19035),
            .in2(N__19200),
            .in3(N__38625),
            .lcout(\b2v_inst.dir_mem_215lt6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un8_dir_mem_2_cry_9_c_RNI1HOE_LC_9_6_4 .C_ON=1'b0;
    defparam \b2v_inst.un8_dir_mem_2_cry_9_c_RNI1HOE_LC_9_6_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un8_dir_mem_2_cry_9_c_RNI1HOE_LC_9_6_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \b2v_inst.un8_dir_mem_2_cry_9_c_RNI1HOE_LC_9_6_4  (
            .in0(_gnd_net_),
            .in1(N__20260),
            .in2(_gnd_net_),
            .in3(N__20241),
            .lcout(\b2v_inst.dir_mem_215lto11_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_RNIBT583_1_LC_9_6_6 .C_ON=1'b0;
    defparam \b2v_inst.indice_RNIBT583_1_LC_9_6_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_RNIBT583_1_LC_9_6_6 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \b2v_inst.indice_RNIBT583_1_LC_9_6_6  (
            .in0(N__18997),
            .in1(N__18979),
            .in2(_gnd_net_),
            .in3(N__17069),
            .lcout(\b2v_inst.dir_mem_215lt7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.energia_temp_4_LC_9_7_1 .C_ON=1'b0;
    defparam \b2v_inst.energia_temp_4_LC_9_7_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.energia_temp_4_LC_9_7_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.energia_temp_4_LC_9_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17185),
            .lcout(b2v_inst_energia_temp_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34482),
            .ce(N__26144),
            .sr(N__38069));
    defparam \b2v_inst.energia_temp_5_LC_9_7_3 .C_ON=1'b0;
    defparam \b2v_inst.energia_temp_5_LC_9_7_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.energia_temp_5_LC_9_7_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.energia_temp_5_LC_9_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17149),
            .lcout(b2v_inst_energia_temp_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34482),
            .ce(N__26144),
            .sr(N__38069));
    defparam \b2v_inst.data_a_escribir_RNO_2_5_LC_9_7_5 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_2_5_LC_9_7_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_2_5_LC_9_7_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_2_5_LC_9_7_5  (
            .in0(N__27398),
            .in1(N__29560),
            .in2(_gnd_net_),
            .in3(N__32535),
            .lcout(\b2v_inst.N_273 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un8_dir_mem_1_cry_4_c_RNIMMVC2_LC_9_7_6 .C_ON=1'b0;
    defparam \b2v_inst.un8_dir_mem_1_cry_4_c_RNIMMVC2_LC_9_7_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un8_dir_mem_1_cry_4_c_RNIMMVC2_LC_9_7_6 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \b2v_inst.un8_dir_mem_1_cry_4_c_RNIMMVC2_LC_9_7_6  (
            .in0(N__18112),
            .in1(N__17987),
            .in2(_gnd_net_),
            .in3(N__17120),
            .lcout(\b2v_inst.dir_mem_115lt7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNIQHR9_22_LC_9_8_7 .C_ON=1'b0;
    defparam \b2v_inst.state_RNIQHR9_22_LC_9_8_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNIQHR9_22_LC_9_8_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst.state_RNIQHR9_22_LC_9_8_7  (
            .in0(_gnd_net_),
            .in1(N__27837),
            .in2(_gnd_net_),
            .in3(N__20972),
            .lcout(\b2v_inst.N_362_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_27_LC_9_9_1 .C_ON=1'b0;
    defparam \b2v_inst.state_27_LC_9_9_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.state_27_LC_9_9_1 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \b2v_inst.state_27_LC_9_9_1  (
            .in0(N__22150),
            .in1(N__31622),
            .in2(_gnd_net_),
            .in3(N__23016),
            .lcout(\b2v_inst.stateZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34460),
            .ce(),
            .sr(N__38064));
    defparam \b2v_inst.state_28_LC_9_9_5 .C_ON=1'b0;
    defparam \b2v_inst.state_28_LC_9_9_5 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.state_28_LC_9_9_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \b2v_inst.state_28_LC_9_9_5  (
            .in0(_gnd_net_),
            .in1(N__32051),
            .in2(_gnd_net_),
            .in3(N__23017),
            .lcout(\b2v_inst.stateZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34460),
            .ce(),
            .sr(N__38064));
    defparam \b2v_inst.state_RNO_29_29_LC_9_10_3 .C_ON=1'b0;
    defparam \b2v_inst.state_RNO_29_29_LC_9_10_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNO_29_29_LC_9_10_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst.state_RNO_29_29_LC_9_10_3  (
            .in0(N__31613),
            .in1(N__20947),
            .in2(N__22169),
            .in3(N__26449),
            .lcout(\b2v_inst.N_618_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNO_23_29_LC_9_11_1 .C_ON=1'b0;
    defparam \b2v_inst.state_RNO_23_29_LC_9_11_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNO_23_29_LC_9_11_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \b2v_inst.state_RNO_23_29_LC_9_11_1  (
            .in0(_gnd_net_),
            .in1(N__26074),
            .in2(_gnd_net_),
            .in3(N__25438),
            .lcout(),
            .ltout(\b2v_inst.g0_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNO_11_29_LC_9_11_2 .C_ON=1'b0;
    defparam \b2v_inst.state_RNO_11_29_LC_9_11_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNO_11_29_LC_9_11_2 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \b2v_inst.state_RNO_11_29_LC_9_11_2  (
            .in0(N__25738),
            .in1(N__25685),
            .in2(N__17114),
            .in3(N__17111),
            .lcout(),
            .ltout(\b2v_inst.g0_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNO_4_29_LC_9_11_3 .C_ON=1'b0;
    defparam \b2v_inst.state_RNO_4_29_LC_9_11_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNO_4_29_LC_9_11_3 .LUT_INIT=16'b1111111111011111;
    LogicCell40 \b2v_inst.state_RNO_4_29_LC_9_11_3  (
            .in0(N__17333),
            .in1(N__38259),
            .in2(N__17345),
            .in3(N__17738),
            .lcout(),
            .ltout(\b2v_inst.G_40_i_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNO_1_29_LC_9_11_4 .C_ON=1'b0;
    defparam \b2v_inst.state_RNO_1_29_LC_9_11_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNO_1_29_LC_9_11_4 .LUT_INIT=16'b0000110100001111;
    LogicCell40 \b2v_inst.state_RNO_1_29_LC_9_11_4  (
            .in0(N__17620),
            .in1(N__17342),
            .in2(N__17336),
            .in3(N__17728),
            .lcout(\b2v_inst.state_RNO_1Z0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNO_12_29_LC_9_11_5 .C_ON=1'b0;
    defparam \b2v_inst.state_RNO_12_29_LC_9_11_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNO_12_29_LC_9_11_5 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \b2v_inst.state_RNO_12_29_LC_9_11_5  (
            .in0(N__28332),
            .in1(N__21892),
            .in2(N__19692),
            .in3(N__19526),
            .lcout(\b2v_inst.state_ns_i_0_a2_11_a2_0_3_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNO_21_29_LC_9_11_7 .C_ON=1'b0;
    defparam \b2v_inst.state_RNO_21_29_LC_9_11_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNO_21_29_LC_9_11_7 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \b2v_inst.state_RNO_21_29_LC_9_11_7  (
            .in0(N__28333),
            .in1(N__17327),
            .in2(N__19693),
            .in3(N__21893),
            .lcout(\b2v_inst.state_ns_i_0_a2_11_o2_4_0_3_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_RX_Byte_7_LC_9_12_0 .C_ON=1'b0;
    defparam \b2v_inst1.r_RX_Byte_7_LC_9_12_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst1.r_RX_Byte_7_LC_9_12_0 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \b2v_inst1.r_RX_Byte_7_LC_9_12_0  (
            .in0(N__22828),
            .in1(N__17321),
            .in2(N__26737),
            .in3(N__17301),
            .lcout(SYNTHESIZED_WIRE_10_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34452),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNO_0_10_LC_9_12_2 .C_ON=1'b0;
    defparam \b2v_inst.state_RNO_0_10_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNO_0_10_LC_9_12_2 .LUT_INIT=16'b1010100010100000;
    LogicCell40 \b2v_inst.state_RNO_0_10_LC_9_12_2  (
            .in0(N__17731),
            .in1(N__17524),
            .in2(N__17381),
            .in3(N__17621),
            .lcout(\b2v_inst.pix_count_anterior5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNO_9_29_LC_9_12_3 .C_ON=1'b0;
    defparam \b2v_inst.state_RNO_9_29_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNO_9_29_LC_9_12_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \b2v_inst.state_RNO_9_29_LC_9_12_3  (
            .in0(N__19525),
            .in1(N__17234),
            .in2(_gnd_net_),
            .in3(N__17228),
            .lcout(\b2v_inst.state_ns_i_0_a2_11_o2_4_0_5_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNO_8_29_LC_9_12_4 .C_ON=1'b0;
    defparam \b2v_inst.state_RNO_8_29_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNO_8_29_LC_9_12_4 .LUT_INIT=16'b1100111011111111;
    LogicCell40 \b2v_inst.state_RNO_8_29_LC_9_12_4  (
            .in0(N__17730),
            .in1(N__27058),
            .in2(N__17861),
            .in3(N__17221),
            .lcout(\b2v_inst.g3_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNO_10_29_LC_9_12_6 .C_ON=1'b0;
    defparam \b2v_inst.state_RNO_10_29_LC_9_12_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNO_10_29_LC_9_12_6 .LUT_INIT=16'b1111101011111000;
    LogicCell40 \b2v_inst.state_RNO_10_29_LC_9_12_6  (
            .in0(N__17729),
            .in1(N__17510),
            .in2(N__17201),
            .in3(N__17447),
            .lcout(\b2v_inst.G_40_i_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNIBA4S1_29_LC_9_13_0 .C_ON=1'b0;
    defparam \b2v_inst.state_RNIBA4S1_29_LC_9_13_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNIBA4S1_29_LC_9_13_0 .LUT_INIT=16'b0111011101111111;
    LogicCell40 \b2v_inst.state_RNIBA4S1_29_LC_9_13_0  (
            .in0(N__17732),
            .in1(N__28136),
            .in2(N__17380),
            .in3(N__17613),
            .lcout(),
            .ltout(\b2v_inst.N_430_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNIO4NID_10_LC_9_13_1 .C_ON=1'b0;
    defparam \b2v_inst.state_RNIO4NID_10_LC_9_13_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNIO4NID_10_LC_9_13_1 .LUT_INIT=16'b0011111100111011;
    LogicCell40 \b2v_inst.state_RNIO4NID_10_LC_9_13_1  (
            .in0(N__17525),
            .in1(N__17882),
            .in2(N__17513),
            .in3(N__17376),
            .lcout(\b2v_inst.N_430_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.g1_0_LC_9_13_2 .C_ON=1'b0;
    defparam \b2v_inst.g1_0_LC_9_13_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.g1_0_LC_9_13_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \b2v_inst.g1_0_LC_9_13_2  (
            .in0(_gnd_net_),
            .in1(N__17509),
            .in2(_gnd_net_),
            .in3(N__17446),
            .lcout(\b2v_inst.g1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_10_LC_9_13_4 .C_ON=1'b0;
    defparam \b2v_inst.state_10_LC_9_13_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.state_10_LC_9_13_4 .LUT_INIT=16'b1100111010001010;
    LogicCell40 \b2v_inst.state_10_LC_9_13_4  (
            .in0(N__25484),
            .in1(N__28137),
            .in2(N__30434),
            .in3(N__17360),
            .lcout(\b2v_inst.stateZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34461),
            .ce(),
            .sr(N__38070));
    defparam \b2v_inst.state_RNIMBKA_10_LC_9_13_5 .C_ON=1'b0;
    defparam \b2v_inst.state_RNIMBKA_10_LC_9_13_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNIMBKA_10_LC_9_13_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \b2v_inst.state_RNIMBKA_10_LC_9_13_5  (
            .in0(_gnd_net_),
            .in1(N__28233),
            .in2(_gnd_net_),
            .in3(N__34582),
            .lcout(\b2v_inst.N_481 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_9_LC_9_13_6 .C_ON=1'b0;
    defparam \b2v_inst.state_9_LC_9_13_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.state_9_LC_9_13_6 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \b2v_inst.state_9_LC_9_13_6  (
            .in0(N__28234),
            .in1(N__18629),
            .in2(N__21303),
            .in3(N__23018),
            .lcout(\b2v_inst.stateZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34461),
            .ce(),
            .sr(N__38070));
    defparam \b2v_inst.dir_energia_RNICN7Q1_0_0_LC_9_14_1 .C_ON=1'b0;
    defparam \b2v_inst.dir_energia_RNICN7Q1_0_0_LC_9_14_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_energia_RNICN7Q1_0_0_LC_9_14_1 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \b2v_inst.dir_energia_RNICN7Q1_0_0_LC_9_14_1  (
            .in0(N__39349),
            .in1(N__39122),
            .in2(N__35827),
            .in3(N__36448),
            .lcout(\b2v_inst.state_ns_0_i_o2_7_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_energia_RNIBM7Q1_0_1_LC_9_14_2 .C_ON=1'b0;
    defparam \b2v_inst.dir_energia_RNIBM7Q1_0_1_LC_9_14_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_energia_RNIBM7Q1_0_1_LC_9_14_2 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \b2v_inst.dir_energia_RNIBM7Q1_0_1_LC_9_14_2  (
            .in0(N__38407),
            .in1(N__35570),
            .in2(N__38909),
            .in3(N__38692),
            .lcout(),
            .ltout(\b2v_inst.state_ns_0_i_o2_6_23_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_energia_RNIOG7I4_0_LC_9_14_3 .C_ON=1'b0;
    defparam \b2v_inst.dir_energia_RNIOG7I4_0_LC_9_14_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_energia_RNIOG7I4_0_LC_9_14_3 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \b2v_inst.dir_energia_RNIOG7I4_0_LC_9_14_3  (
            .in0(_gnd_net_),
            .in1(N__21931),
            .in2(N__17354),
            .in3(N__17351),
            .lcout(\b2v_inst.N_512 ),
            .ltout(\b2v_inst.N_512_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNI3EH15_10_LC_9_14_4 .C_ON=1'b0;
    defparam \b2v_inst.state_RNI3EH15_10_LC_9_14_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNI3EH15_10_LC_9_14_4 .LUT_INIT=16'b0000000000010101;
    LogicCell40 \b2v_inst.state_RNI3EH15_10_LC_9_14_4  (
            .in0(N__23912),
            .in1(N__28338),
            .in2(N__17885),
            .in3(N__28238),
            .lcout(\b2v_inst.N_430_tz ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_energia_RNO_0_0_LC_9_14_7 .C_ON=1'b0;
    defparam \b2v_inst.dir_energia_RNO_0_0_LC_9_14_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_energia_RNO_0_0_LC_9_14_7 .LUT_INIT=16'b1100111000001010;
    LogicCell40 \b2v_inst.dir_energia_RNO_0_0_LC_9_14_7  (
            .in0(N__28239),
            .in1(N__34973),
            .in2(N__21302),
            .in3(N__23913),
            .lcout(\b2v_inst.dir_energia_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_energia_RNIBM7Q1_1_LC_9_15_0 .C_ON=1'b0;
    defparam \b2v_inst.dir_energia_RNIBM7Q1_1_LC_9_15_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_energia_RNIBM7Q1_1_LC_9_15_0 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \b2v_inst.dir_energia_RNIBM7Q1_1_LC_9_15_0  (
            .in0(N__38408),
            .in1(N__35571),
            .in2(N__38910),
            .in3(N__38693),
            .lcout(),
            .ltout(\b2v_inst.g0_4_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_fast_RNITQVP4_19_LC_9_15_1 .C_ON=1'b0;
    defparam \b2v_inst.state_fast_RNITQVP4_19_LC_9_15_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_fast_RNITQVP4_19_LC_9_15_1 .LUT_INIT=16'b1111111100000001;
    LogicCell40 \b2v_inst.state_fast_RNITQVP4_19_LC_9_15_1  (
            .in0(N__17831),
            .in1(N__21935),
            .in2(N__17873),
            .in3(N__26950),
            .lcout(),
            .ltout(\b2v_inst.g0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNI9QDMD_29_LC_9_15_2 .C_ON=1'b0;
    defparam \b2v_inst.state_RNI9QDMD_29_LC_9_15_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNI9QDMD_29_LC_9_15_2 .LUT_INIT=16'b1111101011110010;
    LogicCell40 \b2v_inst.state_RNI9QDMD_29_LC_9_15_2  (
            .in0(N__17870),
            .in1(N__17857),
            .in2(N__17840),
            .in3(N__17837),
            .lcout(\b2v_inst.N_352_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_energia_RNICN7Q1_0_LC_9_15_3 .C_ON=1'b0;
    defparam \b2v_inst.dir_energia_RNICN7Q1_0_LC_9_15_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_energia_RNICN7Q1_0_LC_9_15_3 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \b2v_inst.dir_energia_RNICN7Q1_0_LC_9_15_3  (
            .in0(N__39123),
            .in1(N__36449),
            .in2(N__35812),
            .in3(N__39350),
            .lcout(\b2v_inst.g0_4_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.energia_temp_10_LC_9_16_5 .C_ON=1'b0;
    defparam \b2v_inst.energia_temp_10_LC_9_16_5 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.energia_temp_10_LC_9_16_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.energia_temp_10_LC_9_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17821),
            .lcout(b2v_inst_energia_temp_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34492),
            .ce(N__26198),
            .sr(N__38081));
    defparam \b2v_inst.energia_temp_11_LC_9_17_0 .C_ON=1'b0;
    defparam \b2v_inst.energia_temp_11_LC_9_17_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.energia_temp_11_LC_9_17_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.energia_temp_11_LC_9_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17782),
            .lcout(b2v_inst_energia_temp_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34501),
            .ce(N__26206),
            .sr(N__38088));
    defparam \b2v_inst.energia_temp_7_LC_9_17_4 .C_ON=1'b0;
    defparam \b2v_inst.energia_temp_7_LC_9_17_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.energia_temp_7_LC_9_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.energia_temp_7_LC_9_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17765),
            .lcout(b2v_inst_energia_temp_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34501),
            .ce(N__26206),
            .sr(N__38088));
    defparam \b2v_inst.indice_4_LC_10_5_5 .C_ON=1'b0;
    defparam \b2v_inst.indice_4_LC_10_5_5 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.indice_4_LC_10_5_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \b2v_inst.indice_4_LC_10_5_5  (
            .in0(_gnd_net_),
            .in1(N__22096),
            .in2(_gnd_net_),
            .in3(N__18361),
            .lcout(\b2v_inst.indiceZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34493),
            .ce(N__22046),
            .sr(N__38082));
    defparam \b2v_inst.dir_mem_1_3_LC_10_6_0 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_1_3_LC_10_6_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.dir_mem_1_3_LC_10_6_0 .LUT_INIT=16'b1010101011001010;
    LogicCell40 \b2v_inst.dir_mem_1_3_LC_10_6_0  (
            .in0(N__19060),
            .in1(N__18017),
            .in2(N__19179),
            .in3(N__19247),
            .lcout(\b2v_inst.dir_mem_1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34483),
            .ce(N__19112),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_1_4_LC_10_6_1 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_1_4_LC_10_6_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.dir_mem_1_4_LC_10_6_1 .LUT_INIT=16'b1101110010001100;
    LogicCell40 \b2v_inst.dir_mem_1_4_LC_10_6_1  (
            .in0(N__19248),
            .in1(N__19036),
            .in2(N__19180),
            .in3(N__18002),
            .lcout(\b2v_inst.dir_mem_1Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34483),
            .ce(N__19112),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_1_6_LC_10_6_2 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_1_6_LC_10_6_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.dir_mem_1_6_LC_10_6_2 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \b2v_inst.dir_mem_1_6_LC_10_6_2  (
            .in0(N__19168),
            .in1(N__17986),
            .in2(N__17966),
            .in3(N__19246),
            .lcout(\b2v_inst.dir_mem_1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34483),
            .ce(N__19112),
            .sr(_gnd_net_));
    defparam \b2v_inst.un8_dir_mem_2_cry_5_c_RNI14MP3_LC_10_6_6 .C_ON=1'b0;
    defparam \b2v_inst.un8_dir_mem_2_cry_5_c_RNI14MP3_LC_10_6_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un8_dir_mem_2_cry_5_c_RNI14MP3_LC_10_6_6 .LUT_INIT=16'b1000100010000000;
    LogicCell40 \b2v_inst.un8_dir_mem_2_cry_5_c_RNI14MP3_LC_10_6_6  (
            .in0(N__20734),
            .in1(N__20701),
            .in2(N__20779),
            .in3(N__17948),
            .lcout(\b2v_inst.dir_mem_215lt11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un8_dir_mem_1_cry_6_c_RNICBUJ3_LC_10_7_0 .C_ON=1'b0;
    defparam \b2v_inst.un8_dir_mem_1_cry_6_c_RNICBUJ3_LC_10_7_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un8_dir_mem_1_cry_6_c_RNICBUJ3_LC_10_7_0 .LUT_INIT=16'b1000100010000000;
    LogicCell40 \b2v_inst.un8_dir_mem_1_cry_6_c_RNICBUJ3_LC_10_7_0  (
            .in0(N__18166),
            .in1(N__18139),
            .in2(N__17921),
            .in3(N__17942),
            .lcout(\b2v_inst.dir_mem_115lt11 ),
            .ltout(\b2v_inst.dir_mem_115lt11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_1_10_LC_10_7_1 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_1_10_LC_10_7_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.dir_mem_1_10_LC_10_7_1 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \b2v_inst.dir_mem_1_10_LC_10_7_1  (
            .in0(N__18968),
            .in1(N__17936),
            .in2(N__17924),
            .in3(N__18949),
            .lcout(\b2v_inst.dir_mem_1Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34472),
            .ce(N__19104),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_1_0_LC_10_7_3 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_1_0_LC_10_7_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.dir_mem_1_0_LC_10_7_3 .LUT_INIT=16'b1111000011100001;
    LogicCell40 \b2v_inst.dir_mem_1_0_LC_10_7_3  (
            .in0(N__18967),
            .in1(N__19245),
            .in2(N__39316),
            .in3(N__18950),
            .lcout(\b2v_inst.dir_mem_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34472),
            .ce(N__19104),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_1_7_LC_10_7_4 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_1_7_LC_10_7_4 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.dir_mem_1_7_LC_10_7_4 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \b2v_inst.dir_mem_1_7_LC_10_7_4  (
            .in0(N__19242),
            .in1(N__17920),
            .in2(N__17900),
            .in3(N__19167),
            .lcout(\b2v_inst.dir_mem_1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34472),
            .ce(N__19104),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_1_8_LC_10_7_5 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_1_8_LC_10_7_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.dir_mem_1_8_LC_10_7_5 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \b2v_inst.dir_mem_1_8_LC_10_7_5  (
            .in0(N__19165),
            .in1(N__18167),
            .in2(N__18155),
            .in3(N__19243),
            .lcout(\b2v_inst.dir_mem_1Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34472),
            .ce(N__19104),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_1_9_LC_10_7_6 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_1_9_LC_10_7_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.dir_mem_1_9_LC_10_7_6 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \b2v_inst.dir_mem_1_9_LC_10_7_6  (
            .in0(N__19244),
            .in1(N__18140),
            .in2(N__18128),
            .in3(N__19166),
            .lcout(\b2v_inst.dir_mem_1Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34472),
            .ce(N__19104),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_1_5_LC_10_7_7 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_1_5_LC_10_7_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.dir_mem_1_5_LC_10_7_7 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \b2v_inst.dir_mem_1_5_LC_10_7_7  (
            .in0(N__19164),
            .in1(N__18113),
            .in2(N__18089),
            .in3(N__19241),
            .lcout(\b2v_inst.dir_mem_1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34472),
            .ce(N__19104),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_1_LC_10_8_0 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_1_LC_10_8_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.dir_mem_1_LC_10_8_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.dir_mem_1_LC_10_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19282),
            .lcout(\b2v_inst.dir_memZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34462),
            .ce(N__22188),
            .sr(N__38071));
    defparam \b2v_inst.dir_mem_1_RNIGHIR_6_LC_10_9_0 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_1_RNIGHIR_6_LC_10_9_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_1_RNIGHIR_6_LC_10_9_0 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \b2v_inst.dir_mem_1_RNIGHIR_6_LC_10_9_0  (
            .in0(N__25248),
            .in1(N__18074),
            .in2(N__18065),
            .in3(N__25340),
            .lcout(\b2v_inst.addr_ram_iv_i_1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNIFAD9_28_LC_10_9_1 .C_ON=1'b0;
    defparam \b2v_inst.state_RNIFAD9_28_LC_10_9_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNIFAD9_28_LC_10_9_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \b2v_inst.state_RNIFAD9_28_LC_10_9_1  (
            .in0(_gnd_net_),
            .in1(N__22149),
            .in2(_gnd_net_),
            .in3(N__31604),
            .lcout(\b2v_inst.N_450_i_1 ),
            .ltout(\b2v_inst.N_450_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_2_RNI91F21_7_LC_10_9_2 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_2_RNI91F21_7_LC_10_9_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_2_RNI91F21_7_LC_10_9_2 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \b2v_inst.dir_mem_2_RNI91F21_7_LC_10_9_2  (
            .in0(N__20756),
            .in1(N__18050),
            .in2(N__18041),
            .in3(N__22431),
            .lcout(\b2v_inst.addr_ram_iv_i_0_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_2_RNIT4KM_10_LC_10_9_3 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_2_RNIT4KM_10_LC_10_9_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_2_RNIT4KM_10_LC_10_9_3 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \b2v_inst.dir_mem_2_RNIT4KM_10_LC_10_9_3  (
            .in0(N__22430),
            .in1(N__18038),
            .in2(N__20228),
            .in3(N__22499),
            .lcout(\b2v_inst.addr_ram_iv_i_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_1_RNIEFIR_5_LC_10_9_5 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_1_RNIEFIR_5_LC_10_9_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_1_RNIEFIR_5_LC_10_9_5 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \b2v_inst.dir_mem_1_RNIEFIR_5_LC_10_9_5  (
            .in0(N__25339),
            .in1(N__18026),
            .in2(N__18527),
            .in3(N__25249),
            .lcout(\b2v_inst.addr_ram_iv_i_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.cantidad_temp_5_LC_10_10_0 .C_ON=1'b0;
    defparam \b2v_inst.cantidad_temp_5_LC_10_10_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.cantidad_temp_5_LC_10_10_0 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \b2v_inst.cantidad_temp_5_LC_10_10_0  (
            .in0(N__32586),
            .in1(N__34761),
            .in2(N__18512),
            .in3(N__34625),
            .lcout(b2v_inst_cantidad_temp_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34447),
            .ce(),
            .sr(N__38063));
    defparam \b2v_inst.state_0_LC_10_10_2 .C_ON=1'b0;
    defparam \b2v_inst.state_0_LC_10_10_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.state_0_LC_10_10_2 .LUT_INIT=16'b1011101110101010;
    LogicCell40 \b2v_inst.state_0_LC_10_10_2  (
            .in0(N__19691),
            .in1(N__21314),
            .in2(_gnd_net_),
            .in3(N__28339),
            .lcout(\b2v_inst.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34447),
            .ce(),
            .sr(N__38063));
    defparam \b2v_inst.state_24_LC_10_10_4 .C_ON=1'b0;
    defparam \b2v_inst.state_24_LC_10_10_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.state_24_LC_10_10_4 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \b2v_inst.state_24_LC_10_10_4  (
            .in0(N__27059),
            .in1(N__28173),
            .in2(_gnd_net_),
            .in3(N__28526),
            .lcout(\b2v_inst.stateZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34447),
            .ce(),
            .sr(N__38063));
    defparam \b2v_inst.dir_mem_2_RNI3RE21_4_LC_10_11_0 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_2_RNI3RE21_4_LC_10_11_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_2_RNI3RE21_4_LC_10_11_0 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \b2v_inst.dir_mem_2_RNI3RE21_4_LC_10_11_0  (
            .in0(N__18488),
            .in1(N__22531),
            .in2(N__19019),
            .in3(N__22443),
            .lcout(),
            .ltout(\b2v_inst.addr_ram_iv_i_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_RNIN3333_4_LC_10_11_1 .C_ON=1'b0;
    defparam \b2v_inst.indice_RNIN3333_4_LC_10_11_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_RNIN3333_4_LC_10_11_1 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \b2v_inst.indice_RNIN3333_4_LC_10_11_1  (
            .in0(N__18368),
            .in1(N__35166),
            .in2(N__18476),
            .in3(N__36367),
            .lcout(indice_RNIN3333_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_1_RNICDIR_4_LC_10_11_2 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_1_RNICDIR_4_LC_10_11_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_1_RNICDIR_4_LC_10_11_2 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \b2v_inst.dir_mem_1_RNICDIR_4_LC_10_11_2  (
            .in0(N__18377),
            .in1(N__25349),
            .in2(N__18218),
            .in3(N__25260),
            .lcout(\b2v_inst.addr_ram_iv_i_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_3_4_LC_10_11_3 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_3_4_LC_10_11_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.dir_mem_3_4_LC_10_11_3 .LUT_INIT=16'b1010101011001010;
    LogicCell40 \b2v_inst.dir_mem_3_4_LC_10_11_3  (
            .in0(N__36368),
            .in1(N__18362),
            .in2(N__18332),
            .in3(N__18269),
            .lcout(\b2v_inst.dir_mem_3Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34437),
            .ce(N__18203),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNO_15_29_LC_10_12_0 .C_ON=1'b0;
    defparam \b2v_inst.state_RNO_15_29_LC_10_12_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNO_15_29_LC_10_12_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst.state_RNO_15_29_LC_10_12_0  (
            .in0(N__24659),
            .in1(N__33167),
            .in2(N__30931),
            .in3(N__25828),
            .lcout(\b2v_inst.state_ns_i_0_a2_11_o2_4_0_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNO_0_9_LC_10_12_2 .C_ON=1'b0;
    defparam \b2v_inst.state_RNO_0_9_LC_10_12_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNO_0_9_LC_10_12_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \b2v_inst.state_RNO_0_9_LC_10_12_2  (
            .in0(_gnd_net_),
            .in1(N__28337),
            .in2(_gnd_net_),
            .in3(N__34588),
            .lcout(\b2v_inst.state_ns_0_i_a2_0_0_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNO_16_29_LC_10_12_5 .C_ON=1'b0;
    defparam \b2v_inst.state_RNO_16_29_LC_10_12_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNO_16_29_LC_10_12_5 .LUT_INIT=16'b0000000000110010;
    LogicCell40 \b2v_inst.state_RNO_16_29_LC_10_12_5  (
            .in0(N__27959),
            .in1(N__22444),
            .in2(N__26021),
            .in3(N__25267),
            .lcout(),
            .ltout(\b2v_inst.state_ns_i_0_a2_11_o2_4_0_6_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNO_6_29_LC_10_12_6 .C_ON=1'b0;
    defparam \b2v_inst.state_RNO_6_29_LC_10_12_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNO_6_29_LC_10_12_6 .LUT_INIT=16'b0001111111111111;
    LogicCell40 \b2v_inst.state_RNO_6_29_LC_10_12_6  (
            .in0(N__26014),
            .in1(N__27993),
            .in2(N__18620),
            .in3(N__18617),
            .lcout(),
            .ltout(\b2v_inst.N_4_i_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNO_2_29_LC_10_12_7 .C_ON=1'b0;
    defparam \b2v_inst.state_RNO_2_29_LC_10_12_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNO_2_29_LC_10_12_7 .LUT_INIT=16'b0000000100000011;
    LogicCell40 \b2v_inst.state_RNO_2_29_LC_10_12_7  (
            .in0(N__28138),
            .in1(N__18611),
            .in2(N__18602),
            .in3(N__18599),
            .lcout(\b2v_inst.state_RNO_2Z0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_energia_RNIBUMB2_8_LC_10_13_1 .C_ON=1'b0;
    defparam \b2v_inst.dir_energia_RNIBUMB2_8_LC_10_13_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_energia_RNIBUMB2_8_LC_10_13_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst.dir_energia_RNIBUMB2_8_LC_10_13_1  (
            .in0(N__18593),
            .in1(N__39138),
            .in2(_gnd_net_),
            .in3(N__21710),
            .lcout(\b2v_inst.addr_ram_energia_m0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_32_rep1_RNIRV8V_LC_10_13_3 .C_ON=1'b0;
    defparam \b2v_inst.state_32_rep1_RNIRV8V_LC_10_13_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_32_rep1_RNIRV8V_LC_10_13_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \b2v_inst.state_32_rep1_RNIRV8V_LC_10_13_3  (
            .in0(N__25537),
            .in1(N__21258),
            .in2(N__27909),
            .in3(N__20210),
            .lcout(\b2v_inst.N_480 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNO_3_29_LC_10_13_4 .C_ON=1'b0;
    defparam \b2v_inst.state_RNO_3_29_LC_10_13_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNO_3_29_LC_10_13_4 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \b2v_inst.state_RNO_3_29_LC_10_13_4  (
            .in0(N__20211),
            .in1(N__25538),
            .in2(N__21265),
            .in3(N__18557),
            .lcout(),
            .ltout(\b2v_inst.state_ns_i_0_a2_11_o2_4_0_7_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_29_LC_10_13_5 .C_ON=1'b0;
    defparam \b2v_inst.state_29_LC_10_13_5 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.state_29_LC_10_13_5 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \b2v_inst.state_29_LC_10_13_5  (
            .in0(N__18551),
            .in1(N__19388),
            .in2(N__18545),
            .in3(N__18542),
            .lcout(\b2v_inst.stateZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34453),
            .ce(),
            .sr(N__38074));
    defparam \b2v_inst.dir_energia_0_LC_10_14_1 .C_ON=1'b0;
    defparam \b2v_inst.dir_energia_0_LC_10_14_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.dir_energia_0_LC_10_14_1 .LUT_INIT=16'b1000110111011000;
    LogicCell40 \b2v_inst.dir_energia_0_LC_10_14_1  (
            .in0(N__23872),
            .in1(N__18533),
            .in2(N__37133),
            .in3(N__39359),
            .lcout(\b2v_inst.dir_energiaZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34463),
            .ce(N__23800),
            .sr(N__38076));
    defparam \b2v_inst.dir_energia_10_LC_10_14_2 .C_ON=1'b0;
    defparam \b2v_inst.dir_energia_10_LC_10_14_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.dir_energia_10_LC_10_14_2 .LUT_INIT=16'b1111001110101010;
    LogicCell40 \b2v_inst.dir_energia_10_LC_10_14_2  (
            .in0(N__23996),
            .in1(N__23914),
            .in2(N__33686),
            .in3(N__23873),
            .lcout(\b2v_inst.dir_energiaZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34463),
            .ce(N__23800),
            .sr(N__38076));
    defparam \b2v_inst.dir_energia_2_LC_10_14_3 .C_ON=1'b0;
    defparam \b2v_inst.dir_energia_2_LC_10_14_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.dir_energia_2_LC_10_14_3 .LUT_INIT=16'b1101100011111010;
    LogicCell40 \b2v_inst.dir_energia_2_LC_10_14_3  (
            .in0(N__23870),
            .in1(N__33139),
            .in2(N__23588),
            .in3(N__23969),
            .lcout(\b2v_inst.dir_energiaZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34463),
            .ce(N__23800),
            .sr(N__38076));
    defparam \b2v_inst.dir_energia_4_LC_10_14_4 .C_ON=1'b0;
    defparam \b2v_inst.dir_energia_4_LC_10_14_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.dir_energia_4_LC_10_14_4 .LUT_INIT=16'b1011101111110000;
    LogicCell40 \b2v_inst.dir_energia_4_LC_10_14_4  (
            .in0(N__33337),
            .in1(N__23915),
            .in2(N__23555),
            .in3(N__23875),
            .lcout(\b2v_inst.dir_energiaZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34463),
            .ce(N__23800),
            .sr(N__38076));
    defparam \b2v_inst.dir_energia_1_LC_10_14_5 .C_ON=1'b0;
    defparam \b2v_inst.dir_energia_1_LC_10_14_5 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.dir_energia_1_LC_10_14_5 .LUT_INIT=16'b1111011110100010;
    LogicCell40 \b2v_inst.dir_energia_1_LC_10_14_5  (
            .in0(N__23869),
            .in1(N__23967),
            .in2(N__34844),
            .in3(N__23603),
            .lcout(\b2v_inst.dir_energiaZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34463),
            .ce(N__23800),
            .sr(N__38076));
    defparam \b2v_inst.dir_energia_3_LC_10_14_6 .C_ON=1'b0;
    defparam \b2v_inst.dir_energia_3_LC_10_14_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.dir_energia_3_LC_10_14_6 .LUT_INIT=16'b1100111110101010;
    LogicCell40 \b2v_inst.dir_energia_3_LC_10_14_6  (
            .in0(N__23570),
            .in1(N__33256),
            .in2(N__23977),
            .in3(N__23874),
            .lcout(\b2v_inst.dir_energiaZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34463),
            .ce(N__23800),
            .sr(N__38076));
    defparam \b2v_inst.dir_energia_5_LC_10_14_7 .C_ON=1'b0;
    defparam \b2v_inst.dir_energia_5_LC_10_14_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.dir_energia_5_LC_10_14_7 .LUT_INIT=16'b1111011110100010;
    LogicCell40 \b2v_inst.dir_energia_5_LC_10_14_7  (
            .in0(N__23871),
            .in1(N__23968),
            .in2(N__37631),
            .in3(N__23534),
            .lcout(\b2v_inst.dir_energiaZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34463),
            .ce(N__23800),
            .sr(N__38076));
    defparam \b2v_inst.dir_energia_6_LC_10_15_0 .C_ON=1'b0;
    defparam \b2v_inst.dir_energia_6_LC_10_15_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.dir_energia_6_LC_10_15_0 .LUT_INIT=16'b1111010111001100;
    LogicCell40 \b2v_inst.dir_energia_6_LC_10_15_0  (
            .in0(N__23948),
            .in1(N__24056),
            .in2(N__35330),
            .in3(N__23867),
            .lcout(\b2v_inst.dir_energiaZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34473),
            .ce(N__23799),
            .sr(N__38083));
    defparam \b2v_inst.dir_energia_RNI7QMB2_6_LC_10_15_1 .C_ON=1'b0;
    defparam \b2v_inst.dir_energia_RNI7QMB2_6_LC_10_15_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_energia_RNI7QMB2_6_LC_10_15_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst.dir_energia_RNI7QMB2_6_LC_10_15_1  (
            .in0(N__21709),
            .in1(N__18749),
            .in2(_gnd_net_),
            .in3(N__38412),
            .lcout(),
            .ltout(\b2v_inst.addr_ram_energia_m0_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_RNIH7U15_6_LC_10_15_2 .C_ON=1'b0;
    defparam \b2v_inst.indice_RNIH7U15_6_LC_10_15_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_RNIH7U15_6_LC_10_15_2 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \b2v_inst.indice_RNIH7U15_6_LC_10_15_2  (
            .in0(N__38369),
            .in1(N__21636),
            .in2(N__18728),
            .in3(N__35185),
            .lcout(SYNTHESIZED_WIRE_12_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_energia_7_LC_10_15_3 .C_ON=1'b0;
    defparam \b2v_inst.dir_energia_7_LC_10_15_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.dir_energia_7_LC_10_15_3 .LUT_INIT=16'b1101111110001010;
    LogicCell40 \b2v_inst.dir_energia_7_LC_10_15_3  (
            .in0(N__23865),
            .in1(N__35504),
            .in2(N__23976),
            .in3(N__24041),
            .lcout(\b2v_inst.dir_energiaZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34473),
            .ce(N__23799),
            .sr(N__38083));
    defparam \b2v_inst.dir_energia_8_LC_10_15_4 .C_ON=1'b0;
    defparam \b2v_inst.dir_energia_8_LC_10_15_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.dir_energia_8_LC_10_15_4 .LUT_INIT=16'b1111010111001100;
    LogicCell40 \b2v_inst.dir_energia_8_LC_10_15_4  (
            .in0(N__23949),
            .in1(N__24026),
            .in2(N__33397),
            .in3(N__23868),
            .lcout(\b2v_inst.dir_energiaZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34473),
            .ce(N__23799),
            .sr(N__38083));
    defparam \b2v_inst.dir_energia_9_LC_10_15_5 .C_ON=1'b0;
    defparam \b2v_inst.dir_energia_9_LC_10_15_5 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.dir_energia_9_LC_10_15_5 .LUT_INIT=16'b1111011110100010;
    LogicCell40 \b2v_inst.dir_energia_9_LC_10_15_5  (
            .in0(N__23866),
            .in1(N__23950),
            .in2(N__32873),
            .in3(N__24011),
            .lcout(\b2v_inst.dir_energiaZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34473),
            .ce(N__23799),
            .sr(N__38083));
    defparam \b2v_inst.dir_energia_RNI9SMB2_7_LC_10_15_6 .C_ON=1'b0;
    defparam \b2v_inst.dir_energia_RNI9SMB2_7_LC_10_15_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_energia_RNI9SMB2_7_LC_10_15_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst.dir_energia_RNI9SMB2_7_LC_10_15_6  (
            .in0(N__18914),
            .in1(N__38905),
            .in2(_gnd_net_),
            .in3(N__21708),
            .lcout(\b2v_inst.addr_ram_energia_m0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_15_LC_10_16_5 .C_ON=1'b0;
    defparam \b2v_inst.state_15_LC_10_16_5 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.state_15_LC_10_16_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.state_15_LC_10_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19733),
            .lcout(b2v_inst_state_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34484),
            .ce(),
            .sr(N__38089));
    defparam \b2v_inst.energia_temp_12_LC_10_17_6 .C_ON=1'b0;
    defparam \b2v_inst.energia_temp_12_LC_10_17_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.energia_temp_12_LC_10_17_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.energia_temp_12_LC_10_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18874),
            .lcout(b2v_inst_energia_temp_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34494),
            .ce(N__26207),
            .sr(N__38094));
    defparam \b2v_inst.indice_5_LC_11_5_1 .C_ON=1'b0;
    defparam \b2v_inst.indice_5_LC_11_5_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.indice_5_LC_11_5_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \b2v_inst.indice_5_LC_11_5_1  (
            .in0(_gnd_net_),
            .in1(N__22086),
            .in2(_gnd_net_),
            .in3(N__18845),
            .lcout(\b2v_inst.indiceZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34485),
            .ce(N__22057),
            .sr(N__38090));
    defparam \b2v_inst.indice_9_LC_11_5_3 .C_ON=1'b0;
    defparam \b2v_inst.indice_9_LC_11_5_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.indice_9_LC_11_5_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \b2v_inst.indice_9_LC_11_5_3  (
            .in0(_gnd_net_),
            .in1(N__18812),
            .in2(_gnd_net_),
            .in3(N__22088),
            .lcout(\b2v_inst.indiceZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34485),
            .ce(N__22057),
            .sr(N__38090));
    defparam \b2v_inst.indice_7_LC_11_5_4 .C_ON=1'b0;
    defparam \b2v_inst.indice_7_LC_11_5_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.indice_7_LC_11_5_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \b2v_inst.indice_7_LC_11_5_4  (
            .in0(N__22087),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18785),
            .lcout(\b2v_inst.indiceZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34485),
            .ce(N__22057),
            .sr(N__38090));
    defparam \b2v_inst.dir_mem_2_2_LC_11_6_1 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_2_2_LC_11_6_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.dir_mem_2_2_LC_11_6_1 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \b2v_inst.dir_mem_2_2_LC_11_6_1  (
            .in0(N__20679),
            .in1(N__19210),
            .in2(N__21983),
            .in3(N__20638),
            .lcout(\b2v_inst.dir_mem_2Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34474),
            .ce(N__20602),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_2_1_LC_11_6_2 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_2_1_LC_11_6_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.dir_mem_2_1_LC_11_6_2 .LUT_INIT=16'b0000101111110100;
    LogicCell40 \b2v_inst.dir_mem_2_1_LC_11_6_2  (
            .in0(N__20643),
            .in1(N__20684),
            .in2(N__22001),
            .in3(N__38656),
            .lcout(\b2v_inst.dir_mem_2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34474),
            .ce(N__20602),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_2_3_LC_11_6_3 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_2_3_LC_11_6_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.dir_mem_2_3_LC_11_6_3 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \b2v_inst.dir_mem_2_3_LC_11_6_3  (
            .in0(N__20680),
            .in1(N__19067),
            .in2(N__21965),
            .in3(N__20639),
            .lcout(\b2v_inst.dir_mem_2Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34474),
            .ce(N__20602),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_2_4_LC_11_6_5 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_2_4_LC_11_6_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.dir_mem_2_4_LC_11_6_5 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \b2v_inst.dir_mem_2_4_LC_11_6_5  (
            .in0(N__20681),
            .in1(N__19043),
            .in2(N__21950),
            .in3(N__20640),
            .lcout(\b2v_inst.dir_mem_2Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34474),
            .ce(N__20602),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_2_5_LC_11_6_6 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_2_5_LC_11_6_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.dir_mem_2_5_LC_11_6_6 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \b2v_inst.dir_mem_2_5_LC_11_6_6  (
            .in0(N__20641),
            .in1(N__20682),
            .in2(N__22358),
            .in3(N__19004),
            .lcout(\b2v_inst.dir_mem_2Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34474),
            .ce(N__20602),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_2_6_LC_11_6_7 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_2_6_LC_11_6_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.dir_mem_2_6_LC_11_6_7 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \b2v_inst.dir_mem_2_6_LC_11_6_7  (
            .in0(N__20683),
            .in1(N__18986),
            .in2(N__22343),
            .in3(N__20642),
            .lcout(\b2v_inst.dir_mem_2Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34474),
            .ce(N__20602),
            .sr(_gnd_net_));
    defparam \b2v_inst.un8_dir_mem_1_cry_10_c_RNI8DCR_LC_11_7_0 .C_ON=1'b0;
    defparam \b2v_inst.un8_dir_mem_1_cry_10_c_RNI8DCR_LC_11_7_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un8_dir_mem_1_cry_10_c_RNI8DCR_LC_11_7_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \b2v_inst.un8_dir_mem_1_cry_10_c_RNI8DCR_LC_11_7_0  (
            .in0(_gnd_net_),
            .in1(N__18966),
            .in2(_gnd_net_),
            .in3(N__18948),
            .lcout(\b2v_inst.dir_mem_115lto11_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNIULR9_26_LC_11_7_1 .C_ON=1'b0;
    defparam \b2v_inst.state_RNIULR9_26_LC_11_7_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNIULR9_26_LC_11_7_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst.state_RNIULR9_26_LC_11_7_1  (
            .in0(_gnd_net_),
            .in1(N__27839),
            .in2(_gnd_net_),
            .in3(N__20948),
            .lcout(\b2v_inst.N_363_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNISJR9_24_LC_11_7_3 .C_ON=1'b0;
    defparam \b2v_inst.state_RNISJR9_24_LC_11_7_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNISJR9_24_LC_11_7_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst.state_RNISJR9_24_LC_11_7_3  (
            .in0(_gnd_net_),
            .in1(N__27838),
            .in2(_gnd_net_),
            .in3(N__30232),
            .lcout(\b2v_inst.N_463_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_1_RNIKLIR_8_LC_11_7_4 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_1_RNIKLIR_8_LC_11_7_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_1_RNIKLIR_8_LC_11_7_4 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \b2v_inst.dir_mem_1_RNIKLIR_8_LC_11_7_4  (
            .in0(N__18932),
            .in1(N__25358),
            .in2(N__18926),
            .in3(N__25256),
            .lcout(\b2v_inst.addr_ram_iv_i_1_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_RNIBMAH_0_3_LC_11_7_5 .C_ON=1'b0;
    defparam \b2v_inst.indice_RNIBMAH_0_3_LC_11_7_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_RNIBMAH_0_3_LC_11_7_5 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \b2v_inst.indice_RNIBMAH_0_3_LC_11_7_5  (
            .in0(N__35910),
            .in1(N__36347),
            .in2(_gnd_net_),
            .in3(N__36572),
            .lcout(\b2v_inst.un9_indice_0_a2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_1_RNI67IR_1_LC_11_8_0 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_1_RNI67IR_1_LC_11_8_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_1_RNI67IR_1_LC_11_8_0 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \b2v_inst.dir_mem_1_RNI67IR_1_LC_11_8_0  (
            .in0(N__25257),
            .in1(N__19322),
            .in2(N__25366),
            .in3(N__19256),
            .lcout(\b2v_inst.addr_ram_iv_i_0_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_2_RNITKE21_1_LC_11_8_2 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_2_RNITKE21_1_LC_11_8_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_2_RNITKE21_1_LC_11_8_2 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \b2v_inst.dir_mem_2_RNITKE21_1_LC_11_8_2  (
            .in0(N__22406),
            .in1(N__19310),
            .in2(N__19301),
            .in3(N__22511),
            .lcout(\b2v_inst.addr_ram_iv_i_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_1_1_LC_11_8_3 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_1_1_LC_11_8_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.dir_mem_1_1_LC_11_8_3 .LUT_INIT=16'b0000111110001011;
    LogicCell40 \b2v_inst.dir_mem_1_1_LC_11_8_3  (
            .in0(N__19286),
            .in1(N__19178),
            .in2(N__38664),
            .in3(N__19249),
            .lcout(\b2v_inst.dir_mem_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34454),
            .ce(N__19111),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_1_2_LC_11_8_4 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_1_2_LC_11_8_4 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.dir_mem_1_2_LC_11_8_4 .LUT_INIT=16'b1101110010001100;
    LogicCell40 \b2v_inst.dir_mem_1_2_LC_11_8_4  (
            .in0(N__19250),
            .in1(N__19211),
            .in2(N__19181),
            .in3(N__19130),
            .lcout(\b2v_inst.dir_mem_1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34454),
            .ce(N__19111),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNI72D9_24_LC_11_9_0 .C_ON=1'b0;
    defparam \b2v_inst.state_RNI72D9_24_LC_11_9_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNI72D9_24_LC_11_9_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \b2v_inst.state_RNI72D9_24_LC_11_9_0  (
            .in0(_gnd_net_),
            .in1(N__30217),
            .in2(_gnd_net_),
            .in3(N__32896),
            .lcout(\b2v_inst.N_489 ),
            .ltout(\b2v_inst.N_489_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_2_RNI7VE21_6_LC_11_9_1 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_2_RNI7VE21_6_LC_11_9_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_2_RNI7VE21_6_LC_11_9_1 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \b2v_inst.dir_mem_2_RNI7VE21_6_LC_11_9_1  (
            .in0(N__19079),
            .in1(N__21809),
            .in2(N__19070),
            .in3(N__22500),
            .lcout(\b2v_inst.addr_ram_iv_i_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_2_RNIB3F21_8_LC_11_9_3 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_2_RNIB3F21_8_LC_11_9_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_2_RNIB3F21_8_LC_11_9_3 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \b2v_inst.dir_mem_2_RNIB3F21_8_LC_11_9_3  (
            .in0(N__21779),
            .in1(N__22501),
            .in2(N__20723),
            .in3(N__22420),
            .lcout(\b2v_inst.addr_ram_iv_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNI3UC9_22_LC_11_9_4 .C_ON=1'b0;
    defparam \b2v_inst.state_RNI3UC9_22_LC_11_9_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNI3UC9_22_LC_11_9_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \b2v_inst.state_RNI3UC9_22_LC_11_9_4  (
            .in0(_gnd_net_),
            .in1(N__20964),
            .in2(_gnd_net_),
            .in3(N__32024),
            .lcout(\b2v_inst.N_488 ),
            .ltout(\b2v_inst.N_488_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_1_RNIIJIR_7_LC_11_9_5 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_1_RNIIJIR_7_LC_11_9_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_1_RNIIJIR_7_LC_11_9_5 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \b2v_inst.dir_mem_1_RNIIJIR_7_LC_11_9_5  (
            .in0(N__19508),
            .in1(N__19499),
            .in2(N__19484),
            .in3(N__25364),
            .lcout(),
            .ltout(\b2v_inst.addr_ram_iv_i_0_1_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_RNI6J333_7_LC_11_9_6 .C_ON=1'b0;
    defparam \b2v_inst.indice_RNI6J333_7_LC_11_9_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_RNI6J333_7_LC_11_9_6 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \b2v_inst.indice_RNI6J333_7_LC_11_9_6  (
            .in0(N__19481),
            .in1(N__35207),
            .in2(N__19475),
            .in3(N__38843),
            .lcout(indice_RNI6J333_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNO_0_29_LC_11_9_7 .C_ON=1'b0;
    defparam \b2v_inst.state_RNO_0_29_LC_11_9_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNO_0_29_LC_11_9_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst.state_RNO_0_29_LC_11_9_7  (
            .in0(N__22525),
            .in1(N__25255),
            .in2(N__22445),
            .in3(N__25365),
            .lcout(\b2v_inst.state_RNO_0Z0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_26_LC_11_10_3 .C_ON=1'b0;
    defparam \b2v_inst.state_26_LC_11_10_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.state_26_LC_11_10_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \b2v_inst.state_26_LC_11_10_3  (
            .in0(_gnd_net_),
            .in1(N__32899),
            .in2(_gnd_net_),
            .in3(N__23005),
            .lcout(\b2v_inst.stateZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34438),
            .ce(),
            .sr(N__38066));
    defparam \b2v_inst.state_RNIB6D9_26_LC_11_10_4 .C_ON=1'b0;
    defparam \b2v_inst.state_RNIB6D9_26_LC_11_10_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNIB6D9_26_LC_11_10_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \b2v_inst.state_RNIB6D9_26_LC_11_10_4  (
            .in0(_gnd_net_),
            .in1(N__20942),
            .in2(_gnd_net_),
            .in3(N__26441),
            .lcout(\b2v_inst.N_490 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_20_LC_11_10_6 .C_ON=1'b0;
    defparam \b2v_inst.state_20_LC_11_10_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.state_20_LC_11_10_6 .LUT_INIT=16'b0000101000001010;
    LogicCell40 \b2v_inst.state_20_LC_11_10_6  (
            .in0(N__31666),
            .in1(_gnd_net_),
            .in2(N__23015),
            .in3(_gnd_net_),
            .lcout(\b2v_inst.stateZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34438),
            .ce(),
            .sr(N__38066));
    defparam \b2v_inst.state_22_LC_11_10_7 .C_ON=1'b0;
    defparam \b2v_inst.state_22_LC_11_10_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.state_22_LC_11_10_7 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \b2v_inst.state_22_LC_11_10_7  (
            .in0(N__26442),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23004),
            .lcout(\b2v_inst.stateZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34438),
            .ce(),
            .sr(N__38066));
    defparam \b2v_inst.dir_mem_1_RNI45IR_0_LC_11_11_0 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_1_RNI45IR_0_LC_11_11_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_1_RNI45IR_0_LC_11_11_0 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \b2v_inst.dir_mem_1_RNI45IR_0_LC_11_11_0  (
            .in0(N__19376),
            .in1(N__25347),
            .in2(N__19364),
            .in3(N__25259),
            .lcout(\b2v_inst.addr_ram_iv_i_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_2_RNIRIE21_0_LC_11_11_2 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_2_RNIRIE21_0_LC_11_11_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_2_RNIRIE21_0_LC_11_11_2 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \b2v_inst.dir_mem_2_RNIRIE21_0_LC_11_11_2  (
            .in0(N__19532),
            .in1(N__22527),
            .in2(N__20288),
            .in3(N__22438),
            .lcout(\b2v_inst.addr_ram_iv_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_2_RNI1PE21_3_LC_11_11_3 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_2_RNI1PE21_3_LC_11_11_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_2_RNI1PE21_3_LC_11_11_3 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \b2v_inst.dir_mem_2_RNI1PE21_3_LC_11_11_3  (
            .in0(N__22439),
            .in1(N__19346),
            .in2(N__22532),
            .in3(N__19334),
            .lcout(),
            .ltout(\b2v_inst.addr_ram_iv_i_0_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_RNIIU233_3_LC_11_11_4 .C_ON=1'b0;
    defparam \b2v_inst.indice_RNIIU233_3_LC_11_11_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_RNIIU233_3_LC_11_11_4 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \b2v_inst.indice_RNIIU233_3_LC_11_11_4  (
            .in0(N__19538),
            .in1(N__35172),
            .in2(N__19661),
            .in3(N__36573),
            .lcout(indice_RNIIU233_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_1_RNIABIR_3_LC_11_11_5 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_1_RNIABIR_3_LC_11_11_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_1_RNIABIR_3_LC_11_11_5 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \b2v_inst.dir_mem_1_RNIABIR_3_LC_11_11_5  (
            .in0(N__25258),
            .in1(N__19565),
            .in2(N__25363),
            .in3(N__19550),
            .lcout(\b2v_inst.addr_ram_iv_i_0_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_0_LC_11_11_7 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_0_LC_11_11_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.dir_mem_0_LC_11_11_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst.dir_mem_0_LC_11_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39322),
            .lcout(\b2v_inst.dir_memZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34428),
            .ce(N__22186),
            .sr(N__38072));
    defparam \b2v_inst.state_RNIEIRN_4_LC_11_12_0 .C_ON=1'b0;
    defparam \b2v_inst.state_RNIEIRN_4_LC_11_12_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNIEIRN_4_LC_11_12_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst.state_RNIEIRN_4_LC_11_12_0  (
            .in0(N__25457),
            .in1(N__23450),
            .in2(N__23430),
            .in3(N__28045),
            .lcout(\b2v_inst.N_618_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_3_LC_11_12_1 .C_ON=1'b0;
    defparam \b2v_inst.state_3_LC_11_12_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.state_3_LC_11_12_1 .LUT_INIT=16'b1111101011110000;
    LogicCell40 \b2v_inst.state_3_LC_11_12_1  (
            .in0(N__28046),
            .in1(_gnd_net_),
            .in2(N__23458),
            .in3(N__30422),
            .lcout(b2v_inst_state_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34439),
            .ce(),
            .sr(N__38075));
    defparam \b2v_inst.state_7_LC_11_12_2 .C_ON=1'b0;
    defparam \b2v_inst.state_7_LC_11_12_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.state_7_LC_11_12_2 .LUT_INIT=16'b1111101011110000;
    LogicCell40 \b2v_inst.state_7_LC_11_12_2  (
            .in0(N__25458),
            .in1(_gnd_net_),
            .in2(N__23431),
            .in3(N__30421),
            .lcout(b2v_inst_state_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34439),
            .ce(),
            .sr(N__38075));
    defparam \b2v_inst.state_4_LC_11_12_3 .C_ON=1'b0;
    defparam \b2v_inst.state_4_LC_11_12_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.state_4_LC_11_12_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \b2v_inst.state_4_LC_11_12_3  (
            .in0(_gnd_net_),
            .in1(N__21878),
            .in2(_gnd_net_),
            .in3(N__22968),
            .lcout(b2v_inst_state_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34439),
            .ce(),
            .sr(N__38075));
    defparam \b2v_inst.state_8_LC_11_12_4 .C_ON=1'b0;
    defparam \b2v_inst.state_8_LC_11_12_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.state_8_LC_11_12_4 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \b2v_inst.state_8_LC_11_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22995),
            .in3(N__34626),
            .lcout(b2v_inst_state_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34439),
            .ce(),
            .sr(N__38075));
    defparam \b2v_inst9.fsm_state_ns_i_i_0_a2_2_2_0_LC_11_12_5 .C_ON=1'b0;
    defparam \b2v_inst9.fsm_state_ns_i_i_0_a2_2_2_0_LC_11_12_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst9.fsm_state_ns_i_i_0_a2_2_2_0_LC_11_12_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst9.fsm_state_ns_i_i_0_a2_2_2_0_LC_11_12_5  (
            .in0(N__23451),
            .in1(N__23423),
            .in2(N__25672),
            .in3(N__24660),
            .lcout(\b2v_inst9.fsm_state_ns_i_i_0_a2_2_2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_13_LC_11_12_6 .C_ON=1'b0;
    defparam \b2v_inst.state_13_LC_11_12_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.state_13_LC_11_12_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \b2v_inst.state_13_LC_11_12_6  (
            .in0(_gnd_net_),
            .in1(N__30420),
            .in2(_gnd_net_),
            .in3(N__25829),
            .lcout(b2v_inst_state_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34439),
            .ce(),
            .sr(N__38075));
    defparam \b2v_inst.state_RNIB4B9_16_LC_11_13_0 .C_ON=1'b0;
    defparam \b2v_inst.state_RNIB4B9_16_LC_11_13_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNIB4B9_16_LC_11_13_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \b2v_inst.state_RNIB4B9_16_LC_11_13_0  (
            .in0(_gnd_net_),
            .in1(N__21018),
            .in2(_gnd_net_),
            .in3(N__19728),
            .lcout(\b2v_inst.N_514 ),
            .ltout(\b2v_inst.N_514_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNICSQN_4_LC_11_13_1 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNICSQN_4_LC_11_13_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNICSQN_4_LC_11_13_1 .LUT_INIT=16'b0101111100000000;
    LogicCell40 \b2v_inst.data_a_escribir_RNICSQN_4_LC_11_13_1  (
            .in0(N__37680),
            .in1(_gnd_net_),
            .in2(N__19757),
            .in3(N__33325),
            .lcout(N_116_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNI72PL_16_LC_11_13_3 .C_ON=1'b0;
    defparam \b2v_inst.state_RNI72PL_16_LC_11_13_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNI72PL_16_LC_11_13_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \b2v_inst.state_RNI72PL_16_LC_11_13_3  (
            .in0(N__19729),
            .in1(N__26934),
            .in2(N__21023),
            .in3(N__34694),
            .lcout(\b2v_inst.N_477 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_16_LC_11_13_4 .C_ON=1'b0;
    defparam \b2v_inst.state_16_LC_11_13_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.state_16_LC_11_13_4 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \b2v_inst.state_16_LC_11_13_4  (
            .in0(_gnd_net_),
            .in1(N__21022),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst.stateZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34448),
            .ce(),
            .sr(N__38077));
    defparam \b2v_inst.data_a_escribir_RNI3R2E1_4_LC_11_13_5 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNI3R2E1_4_LC_11_13_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNI3R2E1_4_LC_11_13_5 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \b2v_inst.data_a_escribir_RNI3R2E1_4_LC_11_13_5  (
            .in0(N__37679),
            .in1(N__24806),
            .in2(N__33336),
            .in3(N__37404),
            .lcout(N_548_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_fast_19_LC_11_13_7 .C_ON=1'b0;
    defparam \b2v_inst.state_fast_19_LC_11_13_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.state_fast_19_LC_11_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.state_fast_19_LC_11_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30874),
            .lcout(\b2v_inst.state_fastZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34448),
            .ce(),
            .sr(N__38077));
    defparam \b2v_inst.state_RNICIL71_0_LC_11_14_4 .C_ON=1'b0;
    defparam \b2v_inst.state_RNICIL71_0_LC_11_14_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNICIL71_0_LC_11_14_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst.state_RNICIL71_0_LC_11_14_4  (
            .in0(N__28297),
            .in1(N__21864),
            .in2(N__19700),
            .in3(N__20212),
            .lcout(),
            .ltout(\b2v_inst.N_692_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_32_rep1_RNI0G5H1_LC_11_14_5 .C_ON=1'b0;
    defparam \b2v_inst.state_32_rep1_RNI0G5H1_LC_11_14_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_32_rep1_RNI0G5H1_LC_11_14_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \b2v_inst.state_32_rep1_RNI0G5H1_LC_11_14_5  (
            .in0(N__27910),
            .in1(N__25524),
            .in2(N__19664),
            .in3(N__21254),
            .lcout(\b2v_inst.N_247 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNIH20J1_31_LC_11_14_6 .C_ON=1'b0;
    defparam \b2v_inst.state_RNIH20J1_31_LC_11_14_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNIH20J1_31_LC_11_14_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \b2v_inst.state_RNIH20J1_31_LC_11_14_6  (
            .in0(N__21253),
            .in1(N__21827),
            .in2(N__25531),
            .in3(N__20213),
            .lcout(\b2v_inst.N_494 ),
            .ltout(\b2v_inst.N_494_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_energia_RNITFMB2_1_LC_11_14_7 .C_ON=1'b0;
    defparam \b2v_inst.dir_energia_RNITFMB2_1_LC_11_14_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_energia_RNITFMB2_1_LC_11_14_7 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \b2v_inst.dir_energia_RNITFMB2_1_LC_11_14_7  (
            .in0(N__20195),
            .in1(_gnd_net_),
            .in2(N__20171),
            .in3(N__38697),
            .lcout(\b2v_inst.addr_ram_energia_m0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_RNIIBV05_10_LC_11_15_0 .C_ON=1'b0;
    defparam \b2v_inst.indice_RNIIBV05_10_LC_11_15_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_RNIIBV05_10_LC_11_15_0 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \b2v_inst.indice_RNIIBV05_10_LC_11_15_0  (
            .in0(N__21634),
            .in1(N__19778),
            .in2(N__36738),
            .in3(N__35189),
            .lcout(SYNTHESIZED_WIRE_12_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_energia_RNIVHMB2_2_LC_11_15_1 .C_ON=1'b0;
    defparam \b2v_inst.dir_energia_RNIVHMB2_2_LC_11_15_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_energia_RNIVHMB2_2_LC_11_15_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst.dir_energia_RNIVHMB2_2_LC_11_15_1  (
            .in0(N__21707),
            .in1(N__20042),
            .in2(_gnd_net_),
            .in3(N__36146),
            .lcout(),
            .ltout(\b2v_inst.addr_ram_energia_m0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_RNI5RT15_2_LC_11_15_2 .C_ON=1'b0;
    defparam \b2v_inst.indice_RNI5RT15_2_LC_11_15_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_RNI5RT15_2_LC_11_15_2 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \b2v_inst.indice_RNI5RT15_2_LC_11_15_2  (
            .in0(N__21631),
            .in1(N__35186),
            .in2(N__20021),
            .in3(N__36114),
            .lcout(SYNTHESIZED_WIRE_12_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_energia_RNI5OMB2_5_LC_11_15_3 .C_ON=1'b0;
    defparam \b2v_inst.dir_energia_RNI5OMB2_5_LC_11_15_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_energia_RNI5OMB2_5_LC_11_15_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst.dir_energia_RNI5OMB2_5_LC_11_15_3  (
            .in0(N__21706),
            .in1(N__19916),
            .in2(_gnd_net_),
            .in3(N__35577),
            .lcout(),
            .ltout(\b2v_inst.addr_ram_energia_m0_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_RNIE4U15_5_LC_11_15_4 .C_ON=1'b0;
    defparam \b2v_inst.indice_RNIE4U15_5_LC_11_15_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_RNIE4U15_5_LC_11_15_4 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \b2v_inst.indice_RNIE4U15_5_LC_11_15_4  (
            .in0(N__21633),
            .in1(N__35706),
            .in2(N__19904),
            .in3(N__35188),
            .lcout(SYNTHESIZED_WIRE_12_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_energia_RNIT4122_10_LC_11_15_5 .C_ON=1'b0;
    defparam \b2v_inst.dir_energia_RNIT4122_10_LC_11_15_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_energia_RNIT4122_10_LC_11_15_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst.dir_energia_RNIT4122_10_LC_11_15_5  (
            .in0(N__21704),
            .in1(N__19799),
            .in2(_gnd_net_),
            .in3(N__36776),
            .lcout(\b2v_inst.addr_ram_energia_m0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_energia_RNI1KMB2_3_LC_11_15_6 .C_ON=1'b0;
    defparam \b2v_inst.dir_energia_RNI1KMB2_3_LC_11_15_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_energia_RNI1KMB2_3_LC_11_15_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst.dir_energia_RNI1KMB2_3_LC_11_15_6  (
            .in0(N__19772),
            .in1(N__36453),
            .in2(_gnd_net_),
            .in3(N__21705),
            .lcout(),
            .ltout(\b2v_inst.addr_ram_energia_m0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_RNI8UT15_3_LC_11_15_7 .C_ON=1'b0;
    defparam \b2v_inst.indice_RNI8UT15_3_LC_11_15_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_RNI8UT15_3_LC_11_15_7 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \b2v_inst.indice_RNI8UT15_3_LC_11_15_7  (
            .in0(N__35187),
            .in1(N__21632),
            .in2(N__20537),
            .in3(N__36580),
            .lcout(SYNTHESIZED_WIRE_12_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.energia_temp_6_LC_11_16_4 .C_ON=1'b0;
    defparam \b2v_inst.energia_temp_6_LC_11_16_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.energia_temp_6_LC_11_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.energia_temp_6_LC_11_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20425),
            .lcout(b2v_inst_energia_temp_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34475),
            .ce(N__26197),
            .sr(N__38095));
    defparam \b2v_inst.dir_energia_RNIRDMB2_0_LC_11_18_2 .C_ON=1'b0;
    defparam \b2v_inst.dir_energia_RNIRDMB2_0_LC_11_18_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_energia_RNIRDMB2_0_LC_11_18_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst.dir_energia_RNIRDMB2_0_LC_11_18_2  (
            .in0(N__20396),
            .in1(N__39376),
            .in2(_gnd_net_),
            .in3(N__21719),
            .lcout(\b2v_inst.addr_ram_energia_m0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNI9PQN_1_LC_12_4_0 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNI9PQN_1_LC_12_4_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNI9PQN_1_LC_12_4_0 .LUT_INIT=16'b0010001010101010;
    LogicCell40 \b2v_inst.data_a_escribir_RNI9PQN_1_LC_12_4_0  (
            .in0(N__34838),
            .in1(N__37732),
            .in2(_gnd_net_),
            .in3(N__37503),
            .lcout(N_120_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNI1TMA4_32_LC_12_5_0 .C_ON=1'b0;
    defparam \b2v_inst.state_RNI1TMA4_32_LC_12_5_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNI1TMA4_32_LC_12_5_0 .LUT_INIT=16'b1000111100000000;
    LogicCell40 \b2v_inst.state_RNI1TMA4_32_LC_12_5_0  (
            .in0(N__27997),
            .in1(N__27960),
            .in2(N__25951),
            .in3(N__20582),
            .lcout(\b2v_inst.N_432_1 ),
            .ltout(\b2v_inst.N_432_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_10_LC_12_5_1 .C_ON=1'b0;
    defparam \b2v_inst.indice_10_LC_12_5_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.indice_10_LC_12_5_1 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \b2v_inst.indice_10_LC_12_5_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20357),
            .in3(N__20354),
            .lcout(\b2v_inst.indiceZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34476),
            .ce(N__22056),
            .sr(N__38096));
    defparam \b2v_inst.indice_8_LC_12_5_7 .C_ON=1'b0;
    defparam \b2v_inst.indice_8_LC_12_5_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.indice_8_LC_12_5_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \b2v_inst.indice_8_LC_12_5_7  (
            .in0(_gnd_net_),
            .in1(N__20321),
            .in2(_gnd_net_),
            .in3(N__22085),
            .lcout(\b2v_inst.indiceZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34476),
            .ce(N__22056),
            .sr(N__38096));
    defparam \b2v_inst.dir_mem_2_0_LC_12_6_0 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_2_0_LC_12_6_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.dir_mem_2_0_LC_12_6_0 .LUT_INIT=16'b0101010101010110;
    LogicCell40 \b2v_inst.dir_mem_2_0_LC_12_6_0  (
            .in0(N__39227),
            .in1(N__20248),
            .in2(N__20270),
            .in3(N__20645),
            .lcout(\b2v_inst.dir_mem_2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34464),
            .ce(N__20606),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_2_10_LC_12_6_1 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_2_10_LC_12_6_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.dir_mem_2_10_LC_12_6_1 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \b2v_inst.dir_mem_2_10_LC_12_6_1  (
            .in0(N__20646),
            .in1(N__20269),
            .in2(N__22286),
            .in3(N__20249),
            .lcout(\b2v_inst.dir_mem_2Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34464),
            .ce(N__20606),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_2_7_LC_12_6_2 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_2_7_LC_12_6_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.dir_mem_2_7_LC_12_6_2 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \b2v_inst.dir_mem_2_7_LC_12_6_2  (
            .in0(N__20783),
            .in1(N__20685),
            .in2(N__22328),
            .in3(N__20644),
            .lcout(\b2v_inst.dir_mem_2Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34464),
            .ce(N__20606),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_2_8_LC_12_6_3 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_2_8_LC_12_6_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.dir_mem_2_8_LC_12_6_3 .LUT_INIT=16'b1101110010001100;
    LogicCell40 \b2v_inst.dir_mem_2_8_LC_12_6_3  (
            .in0(N__20647),
            .in1(N__22313),
            .in2(N__20690),
            .in3(N__20741),
            .lcout(\b2v_inst.dir_mem_2Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34464),
            .ce(N__20606),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_2_9_LC_12_6_4 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_2_9_LC_12_6_4 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.dir_mem_2_9_LC_12_6_4 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \b2v_inst.dir_mem_2_9_LC_12_6_4  (
            .in0(N__20708),
            .in1(N__20689),
            .in2(N__22301),
            .in3(N__20648),
            .lcout(\b2v_inst.dir_mem_2Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34464),
            .ce(N__20606),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_RNIPLHB_0_LC_12_6_5 .C_ON=1'b0;
    defparam \b2v_inst.indice_RNIPLHB_0_LC_12_6_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_RNIPLHB_0_LC_12_6_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \b2v_inst.indice_RNIPLHB_0_LC_12_6_5  (
            .in0(_gnd_net_),
            .in1(N__38793),
            .in2(_gnd_net_),
            .in3(N__39226),
            .lcout(\b2v_inst.N_648_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNIHQTC2_11_LC_12_6_7 .C_ON=1'b0;
    defparam \b2v_inst.state_RNIHQTC2_11_LC_12_6_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNIHQTC2_11_LC_12_6_7 .LUT_INIT=16'b1000111100001111;
    LogicCell40 \b2v_inst.state_RNIHQTC2_11_LC_12_6_7  (
            .in0(N__20591),
            .in1(N__20561),
            .in2(N__26031),
            .in3(N__23749),
            .lcout(\b2v_inst.N_432_1_tz ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNIP0281_0_LC_12_7_0 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNIP0281_0_LC_12_7_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNIP0281_0_LC_12_7_0 .LUT_INIT=16'b0101110100001000;
    LogicCell40 \b2v_inst.data_a_escribir_RNIP0281_0_LC_12_7_0  (
            .in0(N__37510),
            .in1(N__34974),
            .in2(N__37759),
            .in3(N__24404),
            .lcout(N_556_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_RNIBMAH_3_LC_12_7_2 .C_ON=1'b0;
    defparam \b2v_inst.indice_RNIBMAH_3_LC_12_7_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_RNIBMAH_3_LC_12_7_2 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \b2v_inst.indice_RNIBMAH_3_LC_12_7_2  (
            .in0(N__39027),
            .in1(N__35682),
            .in2(_gnd_net_),
            .in3(N__36571),
            .lcout(\b2v_inst.indice_4_i_a2_0_7_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNIBRQN_3_LC_12_7_5 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNIBRQN_3_LC_12_7_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNIBRQN_3_LC_12_7_5 .LUT_INIT=16'b0010001010101010;
    LogicCell40 \b2v_inst.data_a_escribir_RNIBRQN_3_LC_12_7_5  (
            .in0(N__33254),
            .in1(N__37728),
            .in2(_gnd_net_),
            .in3(N__37509),
            .lcout(N_117_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNIQFKA_5_LC_12_8_2 .C_ON=1'b0;
    defparam \b2v_inst.state_RNIQFKA_5_LC_12_8_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNIQFKA_5_LC_12_8_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \b2v_inst.state_RNIQFKA_5_LC_12_8_2  (
            .in0(_gnd_net_),
            .in1(N__21882),
            .in2(_gnd_net_),
            .in3(N__34741),
            .lcout(\b2v_inst.N_577_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_1_RNIMNIR_9_LC_12_8_6 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_1_RNIMNIR_9_LC_12_8_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_1_RNIMNIR_9_LC_12_8_6 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \b2v_inst.dir_mem_1_RNIMNIR_9_LC_12_8_6  (
            .in0(N__20888),
            .in1(N__25359),
            .in2(N__20876),
            .in3(N__25254),
            .lcout(\b2v_inst.addr_ram_iv_i_1_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNINBVD1_1_LC_12_9_0 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNINBVD1_1_LC_12_9_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNINBVD1_1_LC_12_9_0 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \b2v_inst.data_a_escribir_RNINBVD1_1_LC_12_9_0  (
            .in0(N__24371),
            .in1(N__37753),
            .in2(N__34839),
            .in3(N__37479),
            .lcout(N_554_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_2_RNIVME21_2_LC_12_9_3 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_2_RNIVME21_2_LC_12_9_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_2_RNIVME21_2_LC_12_9_3 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \b2v_inst.dir_mem_2_RNIVME21_2_LC_12_9_3  (
            .in0(N__22404),
            .in1(N__20843),
            .in2(N__20828),
            .in3(N__22524),
            .lcout(\b2v_inst.addr_ram_iv_i_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_2_RNID5F21_9_LC_12_9_4 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_2_RNID5F21_9_LC_12_9_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_2_RNID5F21_9_LC_12_9_4 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \b2v_inst.dir_mem_2_RNID5F21_9_LC_12_9_4  (
            .in0(N__21746),
            .in1(N__22523),
            .in2(N__20816),
            .in3(N__22405),
            .lcout(\b2v_inst.addr_ram_iv_i_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_1_RNI89IR_2_LC_12_9_5 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_1_RNI89IR_2_LC_12_9_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_1_RNI89IR_2_LC_12_9_5 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \b2v_inst.dir_mem_1_RNI89IR_2_LC_12_9_5  (
            .in0(N__20804),
            .in1(N__25348),
            .in2(N__20798),
            .in3(N__25253),
            .lcout(\b2v_inst.addr_ram_iv_i_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNO_2_31_LC_12_10_0 .C_ON=1'b0;
    defparam \b2v_inst.state_RNO_2_31_LC_12_10_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNO_2_31_LC_12_10_0 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \b2v_inst.state_RNO_2_31_LC_12_10_0  (
            .in0(N__21890),
            .in1(N__20986),
            .in2(_gnd_net_),
            .in3(N__28331),
            .lcout(\b2v_inst.state_ns_a3_i_0_a2_5_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNIG6QI_21_LC_12_10_1 .C_ON=1'b0;
    defparam \b2v_inst.state_RNIG6QI_21_LC_12_10_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNIG6QI_21_LC_12_10_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst.state_RNIG6QI_21_LC_12_10_1  (
            .in0(N__26450),
            .in1(N__32897),
            .in2(N__31667),
            .in3(N__32025),
            .lcout(\b2v_inst.N_829 ),
            .ltout(\b2v_inst.N_829_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNIHMD31_5_LC_12_10_2 .C_ON=1'b0;
    defparam \b2v_inst.state_RNIHMD31_5_LC_12_10_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNIHMD31_5_LC_12_10_2 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \b2v_inst.state_RNIHMD31_5_LC_12_10_2  (
            .in0(N__21888),
            .in1(N__34725),
            .in2(N__20786),
            .in3(N__34623),
            .lcout(\b2v_inst.un1_data_a_escribir_0_sqmuxa_3_i_i_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_32_rep1_RNIKPV5_LC_12_10_3 .C_ON=1'b0;
    defparam \b2v_inst.state_32_rep1_RNIKPV5_LC_12_10_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_32_rep1_RNIKPV5_LC_12_10_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \b2v_inst.state_32_rep1_RNIKPV5_LC_12_10_3  (
            .in0(_gnd_net_),
            .in1(N__27919),
            .in2(_gnd_net_),
            .in3(N__21889),
            .lcout(),
            .ltout(\b2v_inst.un1_state_23_i_a2_0_a2_0_a2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNI2KE31_9_LC_12_10_4 .C_ON=1'b0;
    defparam \b2v_inst.state_RNI2KE31_9_LC_12_10_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNI2KE31_9_LC_12_10_4 .LUT_INIT=16'b1111111111011111;
    LogicCell40 \b2v_inst.state_RNI2KE31_9_LC_12_10_4  (
            .in0(N__20987),
            .in1(N__34726),
            .in2(N__20975),
            .in3(N__34624),
            .lcout(\b2v_inst.N_547_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_21_LC_12_10_5 .C_ON=1'b0;
    defparam \b2v_inst.state_21_LC_12_10_5 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.state_21_LC_12_10_5 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \b2v_inst.state_21_LC_12_10_5  (
            .in0(N__20968),
            .in1(N__32026),
            .in2(_gnd_net_),
            .in3(N__22996),
            .lcout(\b2v_inst.stateZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34429),
            .ce(),
            .sr(N__38067));
    defparam \b2v_inst.state_23_LC_12_10_6 .C_ON=1'b0;
    defparam \b2v_inst.state_23_LC_12_10_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.state_23_LC_12_10_6 .LUT_INIT=16'b1111111110100000;
    LogicCell40 \b2v_inst.state_23_LC_12_10_6  (
            .in0(N__32898),
            .in1(_gnd_net_),
            .in2(N__23014),
            .in3(N__30233),
            .lcout(\b2v_inst.stateZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34429),
            .ce(),
            .sr(N__38067));
    defparam \b2v_inst.state_25_LC_12_10_7 .C_ON=1'b0;
    defparam \b2v_inst.state_25_LC_12_10_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.state_25_LC_12_10_7 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \b2v_inst.state_25_LC_12_10_7  (
            .in0(N__26451),
            .in1(N__20946),
            .in2(_gnd_net_),
            .in3(N__23000),
            .lcout(\b2v_inst.stateZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34429),
            .ce(),
            .sr(N__38067));
    defparam \b2v_inst.cuenta_RNI6BB31_6_LC_12_11_0 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_RNI6BB31_6_LC_12_11_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.cuenta_RNI6BB31_6_LC_12_11_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst.cuenta_RNI6BB31_6_LC_12_11_0  (
            .in0(N__23153),
            .in1(N__20918),
            .in2(N__23117),
            .in3(N__23297),
            .lcout(\b2v_inst.un2_cuentalto10_i_a2_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.cuenta_RNI2E6K_2_LC_12_11_2 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_RNI2E6K_2_LC_12_11_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.cuenta_RNI2E6K_2_LC_12_11_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst.cuenta_RNI2E6K_2_LC_12_11_2  (
            .in0(N__23185),
            .in1(N__23215),
            .in2(N__24209),
            .in3(N__23248),
            .lcout(\b2v_inst.un2_cuentalto10_i_a2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_SM_Main_ns_2_0__m16_0_a3_0_LC_12_11_3 .C_ON=1'b0;
    defparam \b2v_inst1.r_SM_Main_ns_2_0__m16_0_a3_0_LC_12_11_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_SM_Main_ns_2_0__m16_0_a3_0_LC_12_11_3 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \b2v_inst1.r_SM_Main_ns_2_0__m16_0_a3_0_LC_12_11_3  (
            .in0(N__22619),
            .in1(N__21190),
            .in2(N__21076),
            .in3(N__22786),
            .lcout(),
            .ltout(\b2v_inst1.m16_0_a3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_SM_Main_1_LC_12_11_4 .C_ON=1'b0;
    defparam \b2v_inst1.r_SM_Main_1_LC_12_11_4 .SEQ_MODE=4'b1000;
    defparam \b2v_inst1.r_SM_Main_1_LC_12_11_4 .LUT_INIT=16'b1111100011111010;
    LogicCell40 \b2v_inst1.r_SM_Main_1_LC_12_11_4  (
            .in0(N__22863),
            .in1(N__20912),
            .in2(N__20891),
            .in3(N__22620),
            .lcout(\b2v_inst1.r_SM_MainZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34420),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_Clk_Count_RNO_1_1_LC_12_11_5 .C_ON=1'b0;
    defparam \b2v_inst1.r_Clk_Count_RNO_1_1_LC_12_11_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_Clk_Count_RNO_1_1_LC_12_11_5 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \b2v_inst1.r_Clk_Count_RNO_1_1_LC_12_11_5  (
            .in0(N__22737),
            .in1(N__22862),
            .in2(_gnd_net_),
            .in3(N__22785),
            .lcout(),
            .ltout(\b2v_inst1.r_Clk_Count_6_iv_0_a3_1_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_Clk_Count_RNO_0_1_LC_12_11_6 .C_ON=1'b0;
    defparam \b2v_inst1.r_Clk_Count_RNO_0_1_LC_12_11_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_Clk_Count_RNO_0_1_LC_12_11_6 .LUT_INIT=16'b1010000010110011;
    LogicCell40 \b2v_inst1.r_Clk_Count_RNO_0_1_LC_12_11_6  (
            .in0(N__21191),
            .in1(N__22738),
            .in2(N__21170),
            .in3(N__21166),
            .lcout(),
            .ltout(\b2v_inst1.r_Clk_Count_6_iv_0_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_Clk_Count_1_LC_12_11_7 .C_ON=1'b0;
    defparam \b2v_inst1.r_Clk_Count_1_LC_12_11_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst1.r_Clk_Count_1_LC_12_11_7 .LUT_INIT=16'b0000011000001100;
    LogicCell40 \b2v_inst1.r_Clk_Count_1_LC_12_11_7  (
            .in0(N__21167),
            .in1(N__21067),
            .in2(N__21122),
            .in3(N__21119),
            .lcout(\b2v_inst1.r_Clk_CountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34420),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNO_0_17_LC_12_12_0 .C_ON=1'b0;
    defparam \b2v_inst.state_RNO_0_17_LC_12_12_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNO_0_17_LC_12_12_0 .LUT_INIT=16'b1010000000100000;
    LogicCell40 \b2v_inst.state_RNO_0_17_LC_12_12_0  (
            .in0(N__37405),
            .in1(N__21008),
            .in2(N__34727),
            .in3(N__20996),
            .lcout(),
            .ltout(\b2v_inst.N_653_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_17_LC_12_12_1 .C_ON=1'b0;
    defparam \b2v_inst.state_17_LC_12_12_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.state_17_LC_12_12_1 .LUT_INIT=16'b1111000011111000;
    LogicCell40 \b2v_inst.state_17_LC_12_12_1  (
            .in0(N__28553),
            .in1(N__37406),
            .in2(N__21026),
            .in3(N__28521),
            .lcout(\b2v_inst.stateZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34430),
            .ce(),
            .sr(N__38078));
    defparam \b2v_inst.state_RNO_1_17_LC_12_12_2 .C_ON=1'b0;
    defparam \b2v_inst.state_RNO_1_17_LC_12_12_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNO_1_17_LC_12_12_2 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \b2v_inst.state_RNO_1_17_LC_12_12_2  (
            .in0(N__23055),
            .in1(N__23496),
            .in2(_gnd_net_),
            .in3(N__23718),
            .lcout(\b2v_inst.state_ns_i_a2_1_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.cuenta_RNIKUJV_0_LC_12_12_3 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_RNIKUJV_0_LC_12_12_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.cuenta_RNIKUJV_0_LC_12_12_3 .LUT_INIT=16'b0000000000001101;
    LogicCell40 \b2v_inst.cuenta_RNIKUJV_0_LC_12_12_3  (
            .in0(N__22936),
            .in1(N__23300),
            .in2(N__24226),
            .in3(N__23170),
            .lcout(),
            .ltout(\b2v_inst.cuenta_RNIKUJVZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.cuenta_RNI5AT71_0_LC_12_12_4 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_RNI5AT71_0_LC_12_12_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.cuenta_RNI5AT71_0_LC_12_12_4 .LUT_INIT=16'b1101100011011000;
    LogicCell40 \b2v_inst.cuenta_RNI5AT71_0_LC_12_12_4  (
            .in0(N__23131),
            .in1(_gnd_net_),
            .in2(N__21002),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\b2v_inst.un20_cuentalto10_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un4_cuenta_cry_1_c_RNICQI02_LC_12_12_5 .C_ON=1'b0;
    defparam \b2v_inst.un4_cuenta_cry_1_c_RNICQI02_LC_12_12_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un4_cuenta_cry_1_c_RNICQI02_LC_12_12_5 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \b2v_inst.un4_cuenta_cry_1_c_RNICQI02_LC_12_12_5  (
            .in0(N__23234),
            .in1(N__23200),
            .in2(N__20999),
            .in3(N__23092),
            .lcout(\b2v_inst.un20_cuentalto10_sx ),
            .ltout(\b2v_inst.un20_cuentalto10_sx_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un4_cuenta_cry_7_c_RNIO18R2_LC_12_12_6 .C_ON=1'b0;
    defparam \b2v_inst.un4_cuenta_cry_7_c_RNIO18R2_LC_12_12_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un4_cuenta_cry_7_c_RNIO18R2_LC_12_12_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst.un4_cuenta_cry_7_c_RNIO18R2_LC_12_12_6  (
            .in0(N__23056),
            .in1(N__23497),
            .in2(N__20990),
            .in3(N__23719),
            .lcout(\b2v_inst.state18_li_0 ),
            .ltout(\b2v_inst.state18_li_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_18_LC_12_12_7 .C_ON=1'b0;
    defparam \b2v_inst.state_18_LC_12_12_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.state_18_LC_12_12_7 .LUT_INIT=16'b1111110011001100;
    LogicCell40 \b2v_inst.state_18_LC_12_12_7  (
            .in0(_gnd_net_),
            .in1(N__23966),
            .in2(N__21476),
            .in3(N__34706),
            .lcout(\b2v_inst.stateZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34430),
            .ce(),
            .sr(N__38078));
    defparam \b2v_inst.state_RNI1MHN_31_LC_12_13_0 .C_ON=1'b0;
    defparam \b2v_inst.state_RNI1MHN_31_LC_12_13_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNI1MHN_31_LC_12_13_0 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \b2v_inst.state_RNI1MHN_31_LC_12_13_0  (
            .in0(N__25529),
            .in1(N__21250),
            .in2(N__25899),
            .in3(N__37384),
            .lcout(N_130_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_30_LC_12_13_1 .C_ON=1'b0;
    defparam \b2v_inst.state_30_LC_12_13_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.state_30_LC_12_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.state_30_LC_12_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25530),
            .lcout(\b2v_inst.stateZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34440),
            .ce(),
            .sr(N__38084));
    defparam \b2v_inst.state_32_LC_12_13_2 .C_ON=1'b0;
    defparam \b2v_inst.state_32_LC_12_13_2 .SEQ_MODE=4'b1011;
    defparam \b2v_inst.state_32_LC_12_13_2 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \b2v_inst.state_32_LC_12_13_2  (
            .in0(_gnd_net_),
            .in1(N__21252),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst.stateZ0Z_32 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34440),
            .ce(),
            .sr(N__38084));
    defparam \b2v_inst.state_fast_32_LC_12_13_3 .C_ON=1'b0;
    defparam \b2v_inst.state_fast_32_LC_12_13_3 .SEQ_MODE=4'b1011;
    defparam \b2v_inst.state_fast_32_LC_12_13_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst.state_fast_32_LC_12_13_3  (
            .in0(N__21251),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst.state_fastZ0Z_32 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34440),
            .ce(),
            .sr(N__38084));
    defparam \b2v_inst.state_5_LC_12_13_5 .C_ON=1'b0;
    defparam \b2v_inst.state_5_LC_12_13_5 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.state_5_LC_12_13_5 .LUT_INIT=16'b1101100010001000;
    LogicCell40 \b2v_inst.state_5_LC_12_13_5  (
            .in0(N__28313),
            .in1(N__21312),
            .in2(N__21891),
            .in3(N__22992),
            .lcout(\b2v_inst.stateZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34440),
            .ce(),
            .sr(N__38084));
    defparam \b2v_inst.state_6_LC_12_13_6 .C_ON=1'b0;
    defparam \b2v_inst.state_6_LC_12_13_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.state_6_LC_12_13_6 .LUT_INIT=16'b0101000011011100;
    LogicCell40 \b2v_inst.state_6_LC_12_13_6  (
            .in0(N__21313),
            .in1(N__25437),
            .in2(N__28252),
            .in3(N__30426),
            .lcout(\b2v_inst.stateZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34440),
            .ce(),
            .sr(N__38084));
    defparam \b2v_inst.state_32_rep1_RNIKTF9_LC_12_14_0 .C_ON=1'b0;
    defparam \b2v_inst.state_32_rep1_RNIKTF9_LC_12_14_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_32_rep1_RNIKTF9_LC_12_14_0 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \b2v_inst.state_32_rep1_RNIKTF9_LC_12_14_0  (
            .in0(N__25528),
            .in1(N__21249),
            .in2(_gnd_net_),
            .in3(N__27886),
            .lcout(\b2v_inst.N_828 ),
            .ltout(\b2v_inst.N_828_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNIRG0E1_2_LC_12_14_1 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNIRG0E1_2_LC_12_14_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNIRG0E1_2_LC_12_14_1 .LUT_INIT=16'b0000101011001100;
    LogicCell40 \b2v_inst.data_a_escribir_RNIRG0E1_2_LC_12_14_1  (
            .in0(N__33135),
            .in1(N__24893),
            .in2(N__21209),
            .in3(N__37397),
            .lcout(N_552_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_energia_RNI13OT_11_LC_12_14_3 .C_ON=1'b0;
    defparam \b2v_inst.dir_energia_RNI13OT_11_LC_12_14_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_energia_RNI13OT_11_LC_12_14_3 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \b2v_inst.dir_energia_RNI13OT_11_LC_12_14_3  (
            .in0(N__36236),
            .in1(N__36780),
            .in2(N__23825),
            .in3(N__36147),
            .lcout(\b2v_inst.state_ns_0_i_o2_8_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNIVL1E1_3_LC_12_14_4 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNIVL1E1_3_LC_12_14_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNIVL1E1_3_LC_12_14_4 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \b2v_inst.data_a_escribir_RNIVL1E1_3_LC_12_14_4  (
            .in0(N__37396),
            .in1(N__37678),
            .in2(N__33255),
            .in3(N__24866),
            .lcout(N_550_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_fast_RNI70OJ_32_LC_12_14_5 .C_ON=1'b0;
    defparam \b2v_inst.state_fast_RNI70OJ_32_LC_12_14_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_fast_RNI70OJ_32_LC_12_14_5 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \b2v_inst.state_fast_RNI70OJ_32_LC_12_14_5  (
            .in0(N__21899),
            .in1(N__28293),
            .in2(_gnd_net_),
            .in3(N__21863),
            .lcout(\b2v_inst.addr_ram_energia_ss0_0_i_o2_i_o2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_6_LC_12_15_0 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_6_LC_12_15_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.dir_mem_6_LC_12_15_0 .LUT_INIT=16'b1110101010101010;
    LogicCell40 \b2v_inst.dir_mem_6_LC_12_15_0  (
            .in0(N__21821),
            .in1(N__22248),
            .in2(N__22271),
            .in3(N__23764),
            .lcout(\b2v_inst.dir_memZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34455),
            .ce(N__22196),
            .sr(N__38097));
    defparam \b2v_inst.dir_mem_8_LC_12_15_1 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_8_LC_12_15_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.dir_mem_8_LC_12_15_1 .LUT_INIT=16'b1111111110000000;
    LogicCell40 \b2v_inst.dir_mem_8_LC_12_15_1  (
            .in0(N__23763),
            .in1(N__22270),
            .in2(N__22250),
            .in3(N__21794),
            .lcout(\b2v_inst.dir_memZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34455),
            .ce(N__22196),
            .sr(N__38097));
    defparam \b2v_inst.dir_mem_9_LC_12_15_2 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_9_LC_12_15_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.dir_mem_9_LC_12_15_2 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \b2v_inst.dir_mem_9_LC_12_15_2  (
            .in0(N__22266),
            .in1(N__23765),
            .in2(N__21764),
            .in3(N__22249),
            .lcout(\b2v_inst.dir_memZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34455),
            .ce(N__22196),
            .sr(N__38097));
    defparam \b2v_inst.dir_energia_RNI3MMB2_4_LC_12_15_5 .C_ON=1'b0;
    defparam \b2v_inst.dir_energia_RNI3MMB2_4_LC_12_15_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_energia_RNI3MMB2_4_LC_12_15_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst.dir_energia_RNI3MMB2_4_LC_12_15_5  (
            .in0(N__21737),
            .in1(N__36247),
            .in2(_gnd_net_),
            .in3(N__21717),
            .lcout(),
            .ltout(\b2v_inst.addr_ram_energia_m0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_RNIB1U15_4_LC_12_15_6 .C_ON=1'b0;
    defparam \b2v_inst.indice_RNIB1U15_4_LC_12_15_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_RNIB1U15_4_LC_12_15_6 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \b2v_inst.indice_RNIB1U15_4_LC_12_15_6  (
            .in0(N__21635),
            .in1(N__35215),
            .in2(N__21599),
            .in3(N__36377),
            .lcout(SYNTHESIZED_WIRE_12_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_RX_Data_R_LC_12_16_1 .C_ON=1'b0;
    defparam \b2v_inst1.r_RX_Data_R_LC_12_16_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst1.r_RX_Data_R_LC_12_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst1.r_RX_Data_R_LC_12_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21494),
            .lcout(\b2v_inst1.r_RX_Data_RZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34465),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_RX_Data_LC_12_16_5 .C_ON=1'b0;
    defparam \b2v_inst1.r_RX_Data_LC_12_16_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst1.r_RX_Data_LC_12_16_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst1.r_RX_Data_LC_12_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22277),
            .lcout(\b2v_inst1.r_RX_DataZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34465),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_RNIEPAH_5_LC_13_5_3 .C_ON=1'b0;
    defparam \b2v_inst.indice_RNIEPAH_5_LC_13_5_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_RNIEPAH_5_LC_13_5_3 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \b2v_inst.indice_RNIEPAH_5_LC_13_5_3  (
            .in0(N__39026),
            .in1(N__38355),
            .in2(_gnd_net_),
            .in3(N__35683),
            .lcout(\b2v_inst.un9_indice_0_a2_2 ),
            .ltout(\b2v_inst.un9_indice_0_a2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_5_LC_13_5_4 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_5_LC_13_5_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.dir_mem_5_LC_13_5_4 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \b2v_inst.dir_mem_5_LC_13_5_4  (
            .in0(N__22237),
            .in1(N__22214),
            .in2(N__22199),
            .in3(N__23748),
            .lcout(\b2v_inst.dir_memZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34466),
            .ce(N__22195),
            .sr(N__38104));
    defparam \b2v_inst.indice_0_LC_13_6_0 .C_ON=1'b1;
    defparam \b2v_inst.indice_0_LC_13_6_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.indice_0_LC_13_6_0 .LUT_INIT=16'b1011101110111011;
    LogicCell40 \b2v_inst.indice_0_LC_13_6_0  (
            .in0(N__22095),
            .in1(N__39242),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst.indiceZ0Z_0 ),
            .ltout(),
            .carryin(bfn_13_6_0_),
            .carryout(\b2v_inst.un2_dir_mem_2_cry_0 ),
            .clk(N__34456),
            .ce(N__22058),
            .sr(N__38098));
    defparam \b2v_inst.un2_dir_mem_2_cry_0_THRU_LUT4_0_LC_13_6_1 .C_ON=1'b1;
    defparam \b2v_inst.un2_dir_mem_2_cry_0_THRU_LUT4_0_LC_13_6_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un2_dir_mem_2_cry_0_THRU_LUT4_0_LC_13_6_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.un2_dir_mem_2_cry_0_THRU_LUT4_0_LC_13_6_1  (
            .in0(_gnd_net_),
            .in1(N__38646),
            .in2(_gnd_net_),
            .in3(N__21986),
            .lcout(\b2v_inst.un2_dir_mem_2_cry_0_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst.un2_dir_mem_2_cry_0 ),
            .carryout(\b2v_inst.un2_dir_mem_2_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_2_RNO_0_2_LC_13_6_2 .C_ON=1'b1;
    defparam \b2v_inst.dir_mem_2_RNO_0_2_LC_13_6_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_2_RNO_0_2_LC_13_6_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst.dir_mem_2_RNO_0_2_LC_13_6_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__36113),
            .in3(N__21968),
            .lcout(\b2v_inst.dir_mem_2_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\b2v_inst.un2_dir_mem_2_cry_1 ),
            .carryout(\b2v_inst.un2_dir_mem_2_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_2_RNO_0_3_LC_13_6_3 .C_ON=1'b1;
    defparam \b2v_inst.dir_mem_2_RNO_0_3_LC_13_6_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_2_RNO_0_3_LC_13_6_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.dir_mem_2_RNO_0_3_LC_13_6_3  (
            .in0(_gnd_net_),
            .in1(N__36569),
            .in2(_gnd_net_),
            .in3(N__21953),
            .lcout(\b2v_inst.dir_mem_2_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(\b2v_inst.un2_dir_mem_2_cry_2 ),
            .carryout(\b2v_inst.un2_dir_mem_2_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_2_RNO_0_4_LC_13_6_4 .C_ON=1'b1;
    defparam \b2v_inst.dir_mem_2_RNO_0_4_LC_13_6_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_2_RNO_0_4_LC_13_6_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst.dir_mem_2_RNO_0_4_LC_13_6_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__36375),
            .in3(N__21938),
            .lcout(\b2v_inst.dir_mem_2_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\b2v_inst.un2_dir_mem_2_cry_3 ),
            .carryout(\b2v_inst.un2_dir_mem_2_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_2_RNO_0_5_LC_13_6_5 .C_ON=1'b1;
    defparam \b2v_inst.dir_mem_2_RNO_0_5_LC_13_6_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_2_RNO_0_5_LC_13_6_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst.dir_mem_2_RNO_0_5_LC_13_6_5  (
            .in0(_gnd_net_),
            .in1(N__35711),
            .in2(N__37307),
            .in3(N__22346),
            .lcout(\b2v_inst.dir_mem_2_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\b2v_inst.un2_dir_mem_2_cry_4 ),
            .carryout(\b2v_inst.un2_dir_mem_2_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_2_RNO_0_6_LC_13_6_6 .C_ON=1'b1;
    defparam \b2v_inst.dir_mem_2_RNO_0_6_LC_13_6_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_2_RNO_0_6_LC_13_6_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.dir_mem_2_RNO_0_6_LC_13_6_6  (
            .in0(_gnd_net_),
            .in1(N__38370),
            .in2(_gnd_net_),
            .in3(N__22331),
            .lcout(\b2v_inst.dir_mem_2_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\b2v_inst.un2_dir_mem_2_cry_5 ),
            .carryout(\b2v_inst.un2_dir_mem_2_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_2_RNO_0_7_LC_13_6_7 .C_ON=1'b1;
    defparam \b2v_inst.dir_mem_2_RNO_0_7_LC_13_6_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_2_RNO_0_7_LC_13_6_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst.dir_mem_2_RNO_0_7_LC_13_6_7  (
            .in0(_gnd_net_),
            .in1(N__37263),
            .in2(N__38862),
            .in3(N__22316),
            .lcout(\b2v_inst.dir_mem_2_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(\b2v_inst.un2_dir_mem_2_cry_6 ),
            .carryout(\b2v_inst.un2_dir_mem_2_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_2_RNO_0_8_LC_13_7_0 .C_ON=1'b1;
    defparam \b2v_inst.dir_mem_2_RNO_0_8_LC_13_7_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_2_RNO_0_8_LC_13_7_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.dir_mem_2_RNO_0_8_LC_13_7_0  (
            .in0(_gnd_net_),
            .in1(N__39049),
            .in2(_gnd_net_),
            .in3(N__22304),
            .lcout(\b2v_inst.dir_mem_2_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(bfn_13_7_0_),
            .carryout(\b2v_inst.un2_dir_mem_2_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_2_RNO_0_9_LC_13_7_1 .C_ON=1'b1;
    defparam \b2v_inst.dir_mem_2_RNO_0_9_LC_13_7_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_2_RNO_0_9_LC_13_7_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.dir_mem_2_RNO_0_9_LC_13_7_1  (
            .in0(_gnd_net_),
            .in1(N__35937),
            .in2(_gnd_net_),
            .in3(N__22292),
            .lcout(\b2v_inst.dir_mem_2_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(\b2v_inst.un2_dir_mem_2_cry_8 ),
            .carryout(\b2v_inst.un2_dir_mem_2_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_2_RNO_0_10_LC_13_7_2 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_2_RNO_0_10_LC_13_7_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_2_RNO_0_10_LC_13_7_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \b2v_inst.dir_mem_2_RNO_0_10_LC_13_7_2  (
            .in0(_gnd_net_),
            .in1(N__36697),
            .in2(_gnd_net_),
            .in3(N__22289),
            .lcout(\b2v_inst.dir_mem_2_RNO_0Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.cuenta_6_LC_13_8_1 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_6_LC_13_8_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.cuenta_6_LC_13_8_1 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \b2v_inst.cuenta_6_LC_13_8_1  (
            .in0(N__25955),
            .in1(N__24273),
            .in2(_gnd_net_),
            .in3(N__23135),
            .lcout(\b2v_inst.cuentaZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34441),
            .ce(N__24185),
            .sr(N__38085));
    defparam \b2v_inst.cuenta_7_LC_13_8_2 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_7_LC_13_8_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.cuenta_7_LC_13_8_2 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \b2v_inst.cuenta_7_LC_13_8_2  (
            .in0(N__24274),
            .in1(N__25957),
            .in2(_gnd_net_),
            .in3(N__23096),
            .lcout(\b2v_inst.cuentaZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34441),
            .ce(N__24185),
            .sr(N__38085));
    defparam \b2v_inst.cuenta_8_LC_13_8_3 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_8_LC_13_8_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.cuenta_8_LC_13_8_3 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \b2v_inst.cuenta_8_LC_13_8_3  (
            .in0(N__25956),
            .in1(N__24275),
            .in2(_gnd_net_),
            .in3(N__23060),
            .lcout(\b2v_inst.cuentaZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34441),
            .ce(N__24185),
            .sr(N__38085));
    defparam \b2v_inst.cuenta_9_LC_13_8_4 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_9_LC_13_8_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.cuenta_9_LC_13_8_4 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \b2v_inst.cuenta_9_LC_13_8_4  (
            .in0(N__24276),
            .in1(N__25958),
            .in2(_gnd_net_),
            .in3(N__23501),
            .lcout(\b2v_inst.cuentaZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34441),
            .ce(N__24185),
            .sr(N__38085));
    defparam \b2v_inst1.r_SM_Main_ns_2_0__m13_i_a3_1_LC_13_9_0 .C_ON=1'b0;
    defparam \b2v_inst1.r_SM_Main_ns_2_0__m13_i_a3_1_LC_13_9_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_SM_Main_ns_2_0__m13_i_a3_1_LC_13_9_0 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \b2v_inst1.r_SM_Main_ns_2_0__m13_i_a3_1_LC_13_9_0  (
            .in0(N__22907),
            .in1(N__22812),
            .in2(_gnd_net_),
            .in3(N__22573),
            .lcout(),
            .ltout(\b2v_inst1.N_95_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_SM_Main_0_LC_13_9_1 .C_ON=1'b0;
    defparam \b2v_inst1.r_SM_Main_0_LC_13_9_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst1.r_SM_Main_0_LC_13_9_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst1.r_SM_Main_0_LC_13_9_1  (
            .in0(N__22739),
            .in1(N__22676),
            .in2(N__22661),
            .in3(N__22658),
            .lcout(\b2v_inst1.r_SM_MainZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34431),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_2_RNI5TE21_5_LC_13_9_2 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_2_RNI5TE21_5_LC_13_9_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_2_RNI5TE21_5_LC_13_9_2 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \b2v_inst.dir_mem_2_RNI5TE21_5_LC_13_9_2  (
            .in0(N__22544),
            .in1(N__22526),
            .in2(N__22460),
            .in3(N__22429),
            .lcout(\b2v_inst.addr_ram_iv_i_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.cuenta_RNIN5ML_10_LC_13_9_3 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_RNIN5ML_10_LC_13_9_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.cuenta_RNIN5ML_10_LC_13_9_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst.cuenta_RNIN5ML_10_LC_13_9_3  (
            .in0(N__23512),
            .in1(N__23074),
            .in2(N__23704),
            .in3(N__23273),
            .lcout(\b2v_inst.un2_cuentalto10_i_a2_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst9.data_to_send_esr_RNO_0_5_LC_13_10_1 .C_ON=1'b0;
    defparam \b2v_inst9.data_to_send_esr_RNO_0_5_LC_13_10_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst9.data_to_send_esr_RNO_0_5_LC_13_10_1 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \b2v_inst9.data_to_send_esr_RNO_0_5_LC_13_10_1  (
            .in0(N__24560),
            .in1(N__25013),
            .in2(N__23036),
            .in3(N__30419),
            .lcout(),
            .ltout(\b2v_inst9.data_to_send_10_0_0_0_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst9.data_to_send_esr_5_LC_13_10_2 .C_ON=1'b0;
    defparam \b2v_inst9.data_to_send_esr_5_LC_13_10_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst9.data_to_send_esr_5_LC_13_10_2 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \b2v_inst9.data_to_send_esr_5_LC_13_10_2  (
            .in0(N__25634),
            .in1(N__37597),
            .in2(N__22370),
            .in3(N__24113),
            .lcout(\b2v_inst9.data_to_sendZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34421),
            .ce(N__24590),
            .sr(N__38073));
    defparam \b2v_inst9.data_to_send_esr_RNO_0_4_LC_13_10_3 .C_ON=1'b0;
    defparam \b2v_inst9.data_to_send_esr_RNO_0_4_LC_13_10_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst9.data_to_send_esr_RNO_0_4_LC_13_10_3 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \b2v_inst9.data_to_send_esr_RNO_0_4_LC_13_10_3  (
            .in0(N__24558),
            .in1(N__25061),
            .in2(N__22367),
            .in3(N__30417),
            .lcout(\b2v_inst9.data_to_send_10_0_0_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst9.data_to_send_esr_RNO_0_3_LC_13_10_4 .C_ON=1'b0;
    defparam \b2v_inst9.data_to_send_esr_RNO_0_3_LC_13_10_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst9.data_to_send_esr_RNO_0_3_LC_13_10_4 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \b2v_inst9.data_to_send_esr_RNO_0_3_LC_13_10_4  (
            .in0(N__30418),
            .in1(N__25109),
            .in2(N__24128),
            .in3(N__24559),
            .lcout(),
            .ltout(\b2v_inst9.data_to_send_10_0_0_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst9.data_to_send_esr_3_LC_13_10_5 .C_ON=1'b0;
    defparam \b2v_inst9.data_to_send_esr_3_LC_13_10_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst9.data_to_send_esr_3_LC_13_10_5 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \b2v_inst9.data_to_send_esr_3_LC_13_10_5  (
            .in0(N__33244),
            .in1(N__24437),
            .in2(N__23039),
            .in3(N__25633),
            .lcout(\b2v_inst9.data_to_sendZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34421),
            .ce(N__24590),
            .sr(N__38073));
    defparam \b2v_inst9.data_to_send_esr_6_LC_13_10_6 .C_ON=1'b0;
    defparam \b2v_inst9.data_to_send_esr_6_LC_13_10_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst9.data_to_send_esr_6_LC_13_10_6 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \b2v_inst9.data_to_send_esr_6_LC_13_10_6  (
            .in0(N__25635),
            .in1(N__35326),
            .in2(_gnd_net_),
            .in3(N__24353),
            .lcout(\b2v_inst9.data_to_sendZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34421),
            .ce(N__24590),
            .sr(N__38073));
    defparam \b2v_inst.cuenta_1_LC_13_11_0 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_1_LC_13_11_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.cuenta_1_LC_13_11_0 .LUT_INIT=16'b0100010001000000;
    LogicCell40 \b2v_inst.cuenta_1_LC_13_11_0  (
            .in0(N__24254),
            .in1(N__22937),
            .in2(N__25934),
            .in3(N__22994),
            .lcout(\b2v_inst.cuentaZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34411),
            .ce(N__24181),
            .sr(N__38079));
    defparam \b2v_inst.state_RNI1P613_32_LC_13_11_1 .C_ON=1'b0;
    defparam \b2v_inst.state_RNI1P613_32_LC_13_11_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNI1P613_32_LC_13_11_1 .LUT_INIT=16'b1000101000001010;
    LogicCell40 \b2v_inst.state_RNI1P613_32_LC_13_11_1  (
            .in0(N__23027),
            .in1(N__27983),
            .in2(N__25933),
            .in3(N__27950),
            .lcout(\b2v_inst.N_655 ),
            .ltout(\b2v_inst.N_655_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.cuenta_0_LC_13_11_2 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_0_LC_13_11_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.cuenta_0_LC_13_11_2 .LUT_INIT=16'b1111010111110111;
    LogicCell40 \b2v_inst.cuenta_0_LC_13_11_2  (
            .in0(N__23299),
            .in1(N__25912),
            .in2(N__23021),
            .in3(N__22993),
            .lcout(\b2v_inst.cuentaZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34411),
            .ce(N__24181),
            .sr(N__38079));
    defparam \b2v_inst.cuenta_RNIR03A_1_LC_13_11_3 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_RNIR03A_1_LC_13_11_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.cuenta_RNIR03A_1_LC_13_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst.cuenta_RNIR03A_1_LC_13_11_3  (
            .in0(_gnd_net_),
            .in1(N__23298),
            .in2(_gnd_net_),
            .in3(N__23268),
            .lcout(\b2v_inst.cuenta_RNIR03AZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.cuenta_2_LC_13_11_5 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_2_LC_13_11_5 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.cuenta_2_LC_13_11_5 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \b2v_inst.cuenta_2_LC_13_11_5  (
            .in0(N__25909),
            .in1(N__24255),
            .in2(_gnd_net_),
            .in3(N__23233),
            .lcout(\b2v_inst.cuentaZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34411),
            .ce(N__24181),
            .sr(N__38079));
    defparam \b2v_inst.cuenta_3_LC_13_11_6 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_3_LC_13_11_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.cuenta_3_LC_13_11_6 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \b2v_inst.cuenta_3_LC_13_11_6  (
            .in0(N__24256),
            .in1(N__25911),
            .in2(_gnd_net_),
            .in3(N__23201),
            .lcout(\b2v_inst.cuentaZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34411),
            .ce(N__24181),
            .sr(N__38079));
    defparam \b2v_inst.cuenta_4_LC_13_11_7 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_4_LC_13_11_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.cuenta_4_LC_13_11_7 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \b2v_inst.cuenta_4_LC_13_11_7  (
            .in0(N__25910),
            .in1(N__24257),
            .in2(_gnd_net_),
            .in3(N__23171),
            .lcout(\b2v_inst.cuentaZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34411),
            .ce(N__24181),
            .sr(N__38079));
    defparam \b2v_inst.un4_cuenta_cry_1_c_LC_13_12_0 .C_ON=1'b1;
    defparam \b2v_inst.un4_cuenta_cry_1_c_LC_13_12_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un4_cuenta_cry_1_c_LC_13_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.un4_cuenta_cry_1_c_LC_13_12_0  (
            .in0(_gnd_net_),
            .in1(N__23296),
            .in2(N__23272),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_13_12_0_),
            .carryout(\b2v_inst.un4_cuenta_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un4_cuenta_cry_1_c_RNI9V48_LC_13_12_1 .C_ON=1'b1;
    defparam \b2v_inst.un4_cuenta_cry_1_c_RNI9V48_LC_13_12_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un4_cuenta_cry_1_c_RNI9V48_LC_13_12_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst.un4_cuenta_cry_1_c_RNI9V48_LC_13_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23249),
            .in3(N__23219),
            .lcout(\b2v_inst.un4_cuenta_cry_1_c_RNI9VZ0Z48 ),
            .ltout(),
            .carryin(\b2v_inst.un4_cuenta_cry_1 ),
            .carryout(\b2v_inst.un4_cuenta_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un4_cuenta_cry_2_c_RNIB268_LC_13_12_2 .C_ON=1'b1;
    defparam \b2v_inst.un4_cuenta_cry_2_c_RNIB268_LC_13_12_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un4_cuenta_cry_2_c_RNIB268_LC_13_12_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst.un4_cuenta_cry_2_c_RNIB268_LC_13_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23216),
            .in3(N__23189),
            .lcout(\b2v_inst.un4_cuenta_cry_2_c_RNIBZ0Z268 ),
            .ltout(),
            .carryin(\b2v_inst.un4_cuenta_cry_2 ),
            .carryout(\b2v_inst.un4_cuenta_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un4_cuenta_cry_3_c_RNID578_LC_13_12_3 .C_ON=1'b1;
    defparam \b2v_inst.un4_cuenta_cry_3_c_RNID578_LC_13_12_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un4_cuenta_cry_3_c_RNID578_LC_13_12_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst.un4_cuenta_cry_3_c_RNID578_LC_13_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23186),
            .in3(N__23159),
            .lcout(\b2v_inst.un4_cuenta_cry_3_c_RNIDZ0Z578 ),
            .ltout(),
            .carryin(\b2v_inst.un4_cuenta_cry_3 ),
            .carryout(\b2v_inst.un4_cuenta_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un4_cuenta_cry_4_c_RNIF888_LC_13_12_4 .C_ON=1'b1;
    defparam \b2v_inst.un4_cuenta_cry_4_c_RNIF888_LC_13_12_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un4_cuenta_cry_4_c_RNIF888_LC_13_12_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.un4_cuenta_cry_4_c_RNIF888_LC_13_12_4  (
            .in0(_gnd_net_),
            .in1(N__24205),
            .in2(_gnd_net_),
            .in3(N__23156),
            .lcout(\b2v_inst.un4_cuenta_cry_4_c_RNIFZ0Z888 ),
            .ltout(),
            .carryin(\b2v_inst.un4_cuenta_cry_4 ),
            .carryout(\b2v_inst.un4_cuenta_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un4_cuenta_cry_5_c_RNIHB98_LC_13_12_5 .C_ON=1'b1;
    defparam \b2v_inst.un4_cuenta_cry_5_c_RNIHB98_LC_13_12_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un4_cuenta_cry_5_c_RNIHB98_LC_13_12_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.un4_cuenta_cry_5_c_RNIHB98_LC_13_12_5  (
            .in0(_gnd_net_),
            .in1(N__23152),
            .in2(_gnd_net_),
            .in3(N__23120),
            .lcout(\b2v_inst.un4_cuenta_cry_5_c_RNIHBZ0Z98 ),
            .ltout(),
            .carryin(\b2v_inst.un4_cuenta_cry_5 ),
            .carryout(\b2v_inst.un4_cuenta_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un4_cuenta_cry_6_c_RNIJEA8_LC_13_12_6 .C_ON=1'b1;
    defparam \b2v_inst.un4_cuenta_cry_6_c_RNIJEA8_LC_13_12_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un4_cuenta_cry_6_c_RNIJEA8_LC_13_12_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.un4_cuenta_cry_6_c_RNIJEA8_LC_13_12_6  (
            .in0(_gnd_net_),
            .in1(N__23116),
            .in2(_gnd_net_),
            .in3(N__23081),
            .lcout(\b2v_inst.un4_cuenta_cry_6_c_RNIJEAZ0Z8 ),
            .ltout(),
            .carryin(\b2v_inst.un4_cuenta_cry_6 ),
            .carryout(\b2v_inst.un4_cuenta_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un4_cuenta_cry_7_c_RNILHB8_LC_13_12_7 .C_ON=1'b1;
    defparam \b2v_inst.un4_cuenta_cry_7_c_RNILHB8_LC_13_12_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un4_cuenta_cry_7_c_RNILHB8_LC_13_12_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.un4_cuenta_cry_7_c_RNILHB8_LC_13_12_7  (
            .in0(_gnd_net_),
            .in1(N__23078),
            .in2(_gnd_net_),
            .in3(N__23042),
            .lcout(\b2v_inst.un4_cuenta_cry_7_c_RNILHBZ0Z8 ),
            .ltout(),
            .carryin(\b2v_inst.un4_cuenta_cry_7 ),
            .carryout(\b2v_inst.un4_cuenta_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un4_cuenta_cry_8_c_RNINKC8_LC_13_13_0 .C_ON=1'b1;
    defparam \b2v_inst.un4_cuenta_cry_8_c_RNINKC8_LC_13_13_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un4_cuenta_cry_8_c_RNINKC8_LC_13_13_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.un4_cuenta_cry_8_c_RNINKC8_LC_13_13_0  (
            .in0(_gnd_net_),
            .in1(N__23519),
            .in2(_gnd_net_),
            .in3(N__23483),
            .lcout(\b2v_inst.un4_cuenta_cry_8_c_RNINKCZ0Z8 ),
            .ltout(),
            .carryin(bfn_13_13_0_),
            .carryout(\b2v_inst.un4_cuenta_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un4_cuenta_cry_9_c_RNI01T9_LC_13_13_1 .C_ON=1'b0;
    defparam \b2v_inst.un4_cuenta_cry_9_c_RNI01T9_LC_13_13_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un4_cuenta_cry_9_c_RNI01T9_LC_13_13_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \b2v_inst.un4_cuenta_cry_9_c_RNI01T9_LC_13_13_1  (
            .in0(_gnd_net_),
            .in1(N__23705),
            .in2(_gnd_net_),
            .in3(N__23480),
            .lcout(\b2v_inst.un4_cuenta_cry_9_c_RNI01TZ0Z9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNIFA6E1_7_LC_13_13_2 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNIFA6E1_7_LC_13_13_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNIFA6E1_7_LC_13_13_2 .LUT_INIT=16'b0000110010101010;
    LogicCell40 \b2v_inst.data_a_escribir_RNIFA6E1_7_LC_13_13_2  (
            .in0(N__24701),
            .in1(N__35500),
            .in2(N__37709),
            .in3(N__37449),
            .lcout(N_458_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst9.data_to_send_esr_RNO_1_0_LC_13_13_5 .C_ON=1'b0;
    defparam \b2v_inst9.data_to_send_esr_RNO_1_0_LC_13_13_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst9.data_to_send_esr_RNO_1_0_LC_13_13_5 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \b2v_inst9.data_to_send_esr_RNO_1_0_LC_13_13_5  (
            .in0(N__24548),
            .in1(N__24947),
            .in2(N__24475),
            .in3(N__34910),
            .lcout(\b2v_inst9.data_to_send_10_0_0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst9.fsm_state_RNISRGO_0_LC_13_13_6 .C_ON=1'b0;
    defparam \b2v_inst9.fsm_state_RNISRGO_0_LC_13_13_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst9.fsm_state_RNISRGO_0_LC_13_13_6 .LUT_INIT=16'b0000010100000100;
    LogicCell40 \b2v_inst9.fsm_state_RNISRGO_0_LC_13_13_6  (
            .in0(N__26903),
            .in1(N__23462),
            .in2(N__27206),
            .in3(N__28066),
            .lcout(\b2v_inst9.N_740 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst9.fsm_state_RNI44HO_0_LC_13_13_7 .C_ON=1'b0;
    defparam \b2v_inst9.fsm_state_RNI44HO_0_LC_13_13_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst9.fsm_state_RNI44HO_0_LC_13_13_7 .LUT_INIT=16'b0000000001010100;
    LogicCell40 \b2v_inst9.fsm_state_RNI44HO_0_LC_13_13_7  (
            .in0(N__26902),
            .in1(N__23435),
            .in2(N__25483),
            .in3(N__27203),
            .lcout(\b2v_inst9.N_741 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.energia_temp_0_LC_13_14_0 .C_ON=1'b0;
    defparam \b2v_inst.energia_temp_0_LC_13_14_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.energia_temp_0_LC_13_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.energia_temp_0_LC_13_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23405),
            .lcout(b2v_inst_energia_temp_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34442),
            .ce(N__26180),
            .sr(N__38099));
    defparam \b2v_inst.energia_temp_1_LC_13_14_1 .C_ON=1'b0;
    defparam \b2v_inst.energia_temp_1_LC_13_14_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.energia_temp_1_LC_13_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.energia_temp_1_LC_13_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23371),
            .lcout(b2v_inst_energia_temp_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34442),
            .ce(N__26180),
            .sr(N__38099));
    defparam \b2v_inst.energia_temp_13_LC_13_14_5 .C_ON=1'b0;
    defparam \b2v_inst.energia_temp_13_LC_13_14_5 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.energia_temp_13_LC_13_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.energia_temp_13_LC_13_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23333),
            .lcout(b2v_inst_energia_temp_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34442),
            .ce(N__26180),
            .sr(N__38099));
    defparam \b2v_inst.energia_temp_2_LC_13_14_6 .C_ON=1'b0;
    defparam \b2v_inst.energia_temp_2_LC_13_14_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.energia_temp_2_LC_13_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.energia_temp_2_LC_13_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23681),
            .lcout(b2v_inst_energia_temp_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34442),
            .ce(N__26180),
            .sr(N__38099));
    defparam \b2v_inst.energia_temp_3_LC_13_14_7 .C_ON=1'b0;
    defparam \b2v_inst.energia_temp_3_LC_13_14_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.energia_temp_3_LC_13_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.energia_temp_3_LC_13_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23654),
            .lcout(b2v_inst_energia_temp_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34442),
            .ce(N__26180),
            .sr(N__38099));
    defparam \b2v_inst.data_a_escribir_RNI704E1_5_LC_13_15_1 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNI704E1_5_LC_13_15_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNI704E1_5_LC_13_15_1 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \b2v_inst.data_a_escribir_RNI704E1_5_LC_13_15_1  (
            .in0(N__37681),
            .in1(N__24773),
            .in2(N__37626),
            .in3(N__37465),
            .lcout(N_546_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_energia_cry_c_0_LC_13_16_0 .C_ON=1'b1;
    defparam \b2v_inst.dir_energia_cry_c_0_LC_13_16_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_energia_cry_c_0_LC_13_16_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.dir_energia_cry_c_0_LC_13_16_0  (
            .in0(_gnd_net_),
            .in1(N__39369),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_13_16_0_),
            .carryout(\b2v_inst.dir_energia_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_energia_RNO_0_1_LC_13_16_1 .C_ON=1'b1;
    defparam \b2v_inst.dir_energia_RNO_0_1_LC_13_16_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_energia_RNO_0_1_LC_13_16_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.dir_energia_RNO_0_1_LC_13_16_1  (
            .in0(_gnd_net_),
            .in1(N__38707),
            .in2(_gnd_net_),
            .in3(N__23591),
            .lcout(\b2v_inst.dir_energia_s_1 ),
            .ltout(),
            .carryin(\b2v_inst.dir_energia_cry_0 ),
            .carryout(\b2v_inst.dir_energia_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_energia_RNO_0_2_LC_13_16_2 .C_ON=1'b1;
    defparam \b2v_inst.dir_energia_RNO_0_2_LC_13_16_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_energia_RNO_0_2_LC_13_16_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.dir_energia_RNO_0_2_LC_13_16_2  (
            .in0(_gnd_net_),
            .in1(N__36154),
            .in2(_gnd_net_),
            .in3(N__23573),
            .lcout(\b2v_inst.dir_energia_s_2 ),
            .ltout(),
            .carryin(\b2v_inst.dir_energia_cry_1 ),
            .carryout(\b2v_inst.dir_energia_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_energia_RNO_0_3_LC_13_16_3 .C_ON=1'b1;
    defparam \b2v_inst.dir_energia_RNO_0_3_LC_13_16_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_energia_RNO_0_3_LC_13_16_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.dir_energia_RNO_0_3_LC_13_16_3  (
            .in0(_gnd_net_),
            .in1(N__36463),
            .in2(_gnd_net_),
            .in3(N__23558),
            .lcout(\b2v_inst.dir_energia_s_3 ),
            .ltout(),
            .carryin(\b2v_inst.dir_energia_cry_2 ),
            .carryout(\b2v_inst.dir_energia_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_energia_RNO_0_4_LC_13_16_4 .C_ON=1'b1;
    defparam \b2v_inst.dir_energia_RNO_0_4_LC_13_16_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_energia_RNO_0_4_LC_13_16_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.dir_energia_RNO_0_4_LC_13_16_4  (
            .in0(_gnd_net_),
            .in1(N__36246),
            .in2(_gnd_net_),
            .in3(N__23537),
            .lcout(\b2v_inst.dir_energia_s_4 ),
            .ltout(),
            .carryin(\b2v_inst.dir_energia_cry_3 ),
            .carryout(\b2v_inst.dir_energia_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_energia_RNO_0_5_LC_13_16_5 .C_ON=1'b1;
    defparam \b2v_inst.dir_energia_RNO_0_5_LC_13_16_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_energia_RNO_0_5_LC_13_16_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.dir_energia_RNO_0_5_LC_13_16_5  (
            .in0(_gnd_net_),
            .in1(N__35584),
            .in2(_gnd_net_),
            .in3(N__23522),
            .lcout(\b2v_inst.dir_energia_s_5 ),
            .ltout(),
            .carryin(\b2v_inst.dir_energia_cry_4 ),
            .carryout(\b2v_inst.dir_energia_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_energia_RNO_0_6_LC_13_16_6 .C_ON=1'b1;
    defparam \b2v_inst.dir_energia_RNO_0_6_LC_13_16_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_energia_RNO_0_6_LC_13_16_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.dir_energia_RNO_0_6_LC_13_16_6  (
            .in0(_gnd_net_),
            .in1(N__38422),
            .in2(_gnd_net_),
            .in3(N__24044),
            .lcout(\b2v_inst.dir_energia_s_6 ),
            .ltout(),
            .carryin(\b2v_inst.dir_energia_cry_5 ),
            .carryout(\b2v_inst.dir_energia_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_energia_RNO_0_7_LC_13_16_7 .C_ON=1'b1;
    defparam \b2v_inst.dir_energia_RNO_0_7_LC_13_16_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_energia_RNO_0_7_LC_13_16_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.dir_energia_RNO_0_7_LC_13_16_7  (
            .in0(_gnd_net_),
            .in1(N__38917),
            .in2(_gnd_net_),
            .in3(N__24029),
            .lcout(\b2v_inst.dir_energia_s_7 ),
            .ltout(),
            .carryin(\b2v_inst.dir_energia_cry_6 ),
            .carryout(\b2v_inst.dir_energia_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_energia_RNO_0_8_LC_13_17_0 .C_ON=1'b1;
    defparam \b2v_inst.dir_energia_RNO_0_8_LC_13_17_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_energia_RNO_0_8_LC_13_17_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.dir_energia_RNO_0_8_LC_13_17_0  (
            .in0(_gnd_net_),
            .in1(N__39139),
            .in2(_gnd_net_),
            .in3(N__24014),
            .lcout(\b2v_inst.dir_energia_s_8 ),
            .ltout(),
            .carryin(bfn_13_17_0_),
            .carryout(\b2v_inst.dir_energia_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_energia_RNO_0_9_LC_13_17_1 .C_ON=1'b1;
    defparam \b2v_inst.dir_energia_RNO_0_9_LC_13_17_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_energia_RNO_0_9_LC_13_17_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.dir_energia_RNO_0_9_LC_13_17_1  (
            .in0(_gnd_net_),
            .in1(N__35823),
            .in2(_gnd_net_),
            .in3(N__23999),
            .lcout(\b2v_inst.dir_energia_s_9 ),
            .ltout(),
            .carryin(\b2v_inst.dir_energia_cry_8 ),
            .carryout(\b2v_inst.dir_energia_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_energia_RNO_0_10_LC_13_17_2 .C_ON=1'b1;
    defparam \b2v_inst.dir_energia_RNO_0_10_LC_13_17_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_energia_RNO_0_10_LC_13_17_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.dir_energia_RNO_0_10_LC_13_17_2  (
            .in0(_gnd_net_),
            .in1(N__36787),
            .in2(_gnd_net_),
            .in3(N__23981),
            .lcout(\b2v_inst.dir_energia_s_10 ),
            .ltout(),
            .carryin(\b2v_inst.dir_energia_cry_9 ),
            .carryout(\b2v_inst.dir_energia_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_energia_11_LC_13_17_3 .C_ON=1'b0;
    defparam \b2v_inst.dir_energia_11_LC_13_17_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.dir_energia_11_LC_13_17_3 .LUT_INIT=16'b0101001101011100;
    LogicCell40 \b2v_inst.dir_energia_11_LC_13_17_3  (
            .in0(N__23978),
            .in1(N__23818),
            .in2(N__23882),
            .in3(N__23828),
            .lcout(\b2v_inst.dir_energiaZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34467),
            .ce(N__23804),
            .sr(N__38114));
    defparam \b2v_inst.indice_RNI8UI51_10_LC_14_6_2 .C_ON=1'b0;
    defparam \b2v_inst.indice_RNI8UI51_10_LC_14_6_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_RNI8UI51_10_LC_14_6_2 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \b2v_inst.indice_RNI8UI51_10_LC_14_6_2  (
            .in0(N__23774),
            .in1(N__36096),
            .in2(N__36726),
            .in3(N__38641),
            .lcout(\b2v_inst.un9_indice_0_a2_5_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.cuenta_10_LC_14_7_3 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_10_LC_14_7_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.cuenta_10_LC_14_7_3 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \b2v_inst.cuenta_10_LC_14_7_3  (
            .in0(N__25953),
            .in1(N__24281),
            .in2(_gnd_net_),
            .in3(N__23726),
            .lcout(\b2v_inst.cuentaZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34443),
            .ce(N__24180),
            .sr(N__38100));
    defparam \b2v_inst.cuenta_5_LC_14_8_6 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_5_LC_14_8_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.cuenta_5_LC_14_8_6 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \b2v_inst.cuenta_5_LC_14_8_6  (
            .in0(N__25954),
            .in1(N__24280),
            .in2(_gnd_net_),
            .in3(N__24230),
            .lcout(\b2v_inst.cuentaZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34432),
            .ce(N__24179),
            .sr(N__38091));
    defparam \b2v_inst9.data_to_send_esr_1_LC_14_9_1 .C_ON=1'b0;
    defparam \b2v_inst9.data_to_send_esr_1_LC_14_9_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst9.data_to_send_esr_1_LC_14_9_1 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \b2v_inst9.data_to_send_esr_1_LC_14_9_1  (
            .in0(N__24623),
            .in1(N__24311),
            .in2(_gnd_net_),
            .in3(N__24614),
            .lcout(\b2v_inst9.data_to_sendZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34422),
            .ce(N__24591),
            .sr(N__38086));
    defparam \b2v_inst9.data_to_send_esr_4_LC_14_9_6 .C_ON=1'b0;
    defparam \b2v_inst9.data_to_send_esr_4_LC_14_9_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst9.data_to_send_esr_4_LC_14_9_6 .LUT_INIT=16'b1111111111101010;
    LogicCell40 \b2v_inst9.data_to_send_esr_4_LC_14_9_6  (
            .in0(N__24119),
            .in1(N__25640),
            .in2(N__33341),
            .in3(N__24137),
            .lcout(\b2v_inst9.data_to_sendZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34422),
            .ce(N__24591),
            .sr(N__38086));
    defparam \b2v_inst9.data_to_send_esr_RNO_1_4_LC_14_10_0 .C_ON=1'b0;
    defparam \b2v_inst9.data_to_send_esr_RNO_1_4_LC_14_10_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst9.data_to_send_esr_RNO_1_4_LC_14_10_0 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \b2v_inst9.data_to_send_esr_RNO_1_4_LC_14_10_0  (
            .in0(N__24521),
            .in1(N__32630),
            .in2(N__24488),
            .in3(N__24835),
            .lcout(\b2v_inst9.data_to_send_10_0_0_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst9.data_to_send_esr_RNO_1_5_LC_14_10_3 .C_ON=1'b0;
    defparam \b2v_inst9.data_to_send_esr_RNO_1_5_LC_14_10_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst9.data_to_send_esr_RNO_1_5_LC_14_10_3 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \b2v_inst9.data_to_send_esr_RNO_1_5_LC_14_10_3  (
            .in0(N__24487),
            .in1(N__24522),
            .in2(N__32600),
            .in3(N__24791),
            .lcout(\b2v_inst9.data_to_send_10_0_0_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst9.data_to_send_esr_RNO_2_0_LC_14_10_4 .C_ON=1'b0;
    defparam \b2v_inst9.data_to_send_esr_RNO_2_0_LC_14_10_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst9.data_to_send_esr_RNO_2_0_LC_14_10_4 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \b2v_inst9.data_to_send_esr_RNO_2_0_LC_14_10_4  (
            .in0(N__25632),
            .in1(N__24513),
            .in2(N__34966),
            .in3(N__24425),
            .lcout(\b2v_inst9.data_to_send_10_0_0_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst9.fsm_state_RNI7PQ71_0_LC_14_10_5 .C_ON=1'b0;
    defparam \b2v_inst9.fsm_state_RNI7PQ71_0_LC_14_10_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst9.fsm_state_RNI7PQ71_0_LC_14_10_5 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \b2v_inst9.fsm_state_RNI7PQ71_0_LC_14_10_5  (
            .in0(N__26900),
            .in1(N__24104),
            .in2(N__27204),
            .in3(N__26067),
            .lcout(\b2v_inst9.N_583 ),
            .ltout(\b2v_inst9.N_583_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst9.fsm_state_RNIQAU12_0_LC_14_10_6 .C_ON=1'b0;
    defparam \b2v_inst9.fsm_state_RNIQAU12_0_LC_14_10_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst9.fsm_state_RNIQAU12_0_LC_14_10_6 .LUT_INIT=16'b0000000000000111;
    LogicCell40 \b2v_inst9.fsm_state_RNIQAU12_0_LC_14_10_6  (
            .in0(N__30473),
            .in1(N__27196),
            .in2(N__24092),
            .in3(N__26901),
            .lcout(),
            .ltout(\b2v_inst9.un2_n_fsm_state_0_sqmuxa_2_0_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst9.fsm_state_RNI2D372_0_LC_14_10_7 .C_ON=1'b0;
    defparam \b2v_inst9.fsm_state_RNI2D372_0_LC_14_10_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst9.fsm_state_RNI2D372_0_LC_14_10_7 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \b2v_inst9.fsm_state_RNI2D372_0_LC_14_10_7  (
            .in0(N__24089),
            .in1(_gnd_net_),
            .in2(N__24059),
            .in3(_gnd_net_),
            .lcout(\b2v_inst9.un2_n_fsm_state_0_sqmuxa_2_0_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst9.data_to_send_esr_RNO_0_6_LC_14_11_0 .C_ON=1'b0;
    defparam \b2v_inst9.data_to_send_esr_RNO_0_6_LC_14_11_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst9.data_to_send_esr_RNO_0_6_LC_14_11_0 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \b2v_inst9.data_to_send_esr_RNO_0_6_LC_14_11_0  (
            .in0(N__24514),
            .in1(N__30376),
            .in2(N__24344),
            .in3(N__24764),
            .lcout(\b2v_inst9.data_to_send_10_0_0_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst9.data_to_send_esr_RNO_0_7_LC_14_11_1 .C_ON=1'b0;
    defparam \b2v_inst9.data_to_send_esr_RNO_0_7_LC_14_11_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst9.data_to_send_esr_RNO_0_7_LC_14_11_1 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \b2v_inst9.data_to_send_esr_RNO_0_7_LC_14_11_1  (
            .in0(N__30377),
            .in1(N__35493),
            .in2(N__25639),
            .in3(N__24343),
            .lcout(),
            .ltout(\b2v_inst9.data_to_send_10_0_0_0_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst9.data_to_send_esr_7_LC_14_11_2 .C_ON=1'b0;
    defparam \b2v_inst9.data_to_send_esr_7_LC_14_11_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst9.data_to_send_esr_7_LC_14_11_2 .LUT_INIT=16'b1111101011110000;
    LogicCell40 \b2v_inst9.data_to_send_esr_7_LC_14_11_2  (
            .in0(N__24515),
            .in1(_gnd_net_),
            .in2(N__24347),
            .in3(N__24728),
            .lcout(\b2v_inst9.data_to_sendZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34404),
            .ce(N__24592),
            .sr(N__38087));
    defparam \b2v_inst9.data_to_send_esr_0_LC_14_11_3 .C_ON=1'b0;
    defparam \b2v_inst9.data_to_send_esr_0_LC_14_11_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst9.data_to_send_esr_0_LC_14_11_3 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \b2v_inst9.data_to_send_esr_0_LC_14_11_3  (
            .in0(N__24332),
            .in1(N__24326),
            .in2(_gnd_net_),
            .in3(N__24287),
            .lcout(\b2v_inst9.data_to_sendZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34404),
            .ce(N__24592),
            .sr(N__38087));
    defparam \b2v_inst9.fsm_state_RNIONGO_0_LC_14_11_5 .C_ON=1'b0;
    defparam \b2v_inst9.fsm_state_RNIONGO_0_LC_14_11_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst9.fsm_state_RNIONGO_0_LC_14_11_5 .LUT_INIT=16'b0000010100000100;
    LogicCell40 \b2v_inst9.fsm_state_RNIONGO_0_LC_14_11_5  (
            .in0(N__26899),
            .in1(N__26060),
            .in2(N__27205),
            .in3(N__25419),
            .lcout(\b2v_inst9.N_738 ),
            .ltout(\b2v_inst9.N_738_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst9.data_to_send_esr_RNO_2_1_LC_14_11_6 .C_ON=1'b0;
    defparam \b2v_inst9.data_to_send_esr_RNO_2_1_LC_14_11_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst9.data_to_send_esr_RNO_2_1_LC_14_11_6 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \b2v_inst9.data_to_send_esr_RNO_2_1_LC_14_11_6  (
            .in0(N__34825),
            .in1(N__25628),
            .in2(N__24314),
            .in3(N__24389),
            .lcout(\b2v_inst9.data_to_send_10_0_0_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_14_LC_14_12_1 .C_ON=1'b0;
    defparam \b2v_inst.state_14_LC_14_12_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.state_14_LC_14_12_1 .LUT_INIT=16'b1111101010101010;
    LogicCell40 \b2v_inst.state_14_LC_14_12_1  (
            .in0(N__24662),
            .in1(_gnd_net_),
            .in2(N__30411),
            .in3(N__25816),
            .lcout(b2v_inst_state_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34412),
            .ce(),
            .sr(N__38092));
    defparam \b2v_inst9.fsm_state_RNIP6JC_0_LC_14_12_3 .C_ON=1'b0;
    defparam \b2v_inst9.fsm_state_RNIP6JC_0_LC_14_12_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst9.fsm_state_RNIP6JC_0_LC_14_12_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \b2v_inst9.fsm_state_RNIP6JC_0_LC_14_12_3  (
            .in0(_gnd_net_),
            .in1(N__27146),
            .in2(_gnd_net_),
            .in3(N__26881),
            .lcout(N_478),
            .ltout(N_478_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst9.data_to_send_esr_RNO_0_0_LC_14_12_4 .C_ON=1'b0;
    defparam \b2v_inst9.data_to_send_esr_RNO_0_0_LC_14_12_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst9.data_to_send_esr_RNO_0_0_LC_14_12_4 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \b2v_inst9.data_to_send_esr_RNO_0_0_LC_14_12_4  (
            .in0(N__24302),
            .in1(N__33380),
            .in2(N__24290),
            .in3(N__25774),
            .lcout(\b2v_inst9.data_to_send_10_0_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst9.fsm_state_RNI07UL_0_LC_14_12_5 .C_ON=1'b0;
    defparam \b2v_inst9.fsm_state_RNI07UL_0_LC_14_12_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst9.fsm_state_RNI07UL_0_LC_14_12_5 .LUT_INIT=16'b0000001100000010;
    LogicCell40 \b2v_inst9.fsm_state_RNI07UL_0_LC_14_12_5  (
            .in0(N__24661),
            .in1(N__26882),
            .in2(N__27182),
            .in3(N__25815),
            .lcout(\b2v_inst9.N_832 ),
            .ltout(\b2v_inst9.N_832_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst9.data_to_send_esr_RNO_0_1_LC_14_12_6 .C_ON=1'b0;
    defparam \b2v_inst9.data_to_send_esr_RNO_0_1_LC_14_12_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst9.data_to_send_esr_RNO_0_1_LC_14_12_6 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \b2v_inst9.data_to_send_esr_RNO_0_1_LC_14_12_6  (
            .in0(N__32853),
            .in1(N__24602),
            .in2(N__24626),
            .in3(N__30371),
            .lcout(\b2v_inst9.data_to_send_10_0_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst9.data_to_send_esr_RNO_1_1_LC_14_13_1 .C_ON=1'b0;
    defparam \b2v_inst9.data_to_send_esr_RNO_1_1_LC_14_13_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst9.data_to_send_esr_RNO_1_1_LC_14_13_1 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \b2v_inst9.data_to_send_esr_RNO_1_1_LC_14_13_1  (
            .in0(N__24549),
            .in1(N__26225),
            .in2(N__24476),
            .in3(N__34874),
            .lcout(\b2v_inst9.data_to_send_10_0_0_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst9.data_to_send_esr_RNO_2_2_LC_14_13_2 .C_ON=1'b0;
    defparam \b2v_inst9.data_to_send_esr_RNO_2_2_LC_14_13_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst9.data_to_send_esr_RNO_2_2_LC_14_13_2 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \b2v_inst9.data_to_send_esr_RNO_2_2_LC_14_13_2  (
            .in0(N__24523),
            .in1(N__25624),
            .in2(N__33131),
            .in3(N__24907),
            .lcout(),
            .ltout(\b2v_inst9.data_to_send_10_0_0_2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst9.data_to_send_esr_2_LC_14_13_3 .C_ON=1'b0;
    defparam \b2v_inst9.data_to_send_esr_2_LC_14_13_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst9.data_to_send_esr_2_LC_14_13_3 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \b2v_inst9.data_to_send_esr_2_LC_14_13_3  (
            .in0(_gnd_net_),
            .in1(N__24530),
            .in2(N__24605),
            .in3(N__25748),
            .lcout(\b2v_inst9.data_to_sendZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34423),
            .ce(N__24593),
            .sr(N__38101));
    defparam \b2v_inst9.data_to_send_esr_RNO_1_2_LC_14_13_4 .C_ON=1'b0;
    defparam \b2v_inst9.data_to_send_esr_RNO_1_2_LC_14_13_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst9.data_to_send_esr_RNO_1_2_LC_14_13_4 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \b2v_inst9.data_to_send_esr_RNO_1_2_LC_14_13_4  (
            .in0(N__24466),
            .in1(N__24550),
            .in2(N__25145),
            .in3(N__32660),
            .lcout(\b2v_inst9.data_to_send_10_0_0_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst9.data_to_send_esr_RNO_1_3_LC_14_13_6 .C_ON=1'b0;
    defparam \b2v_inst9.data_to_send_esr_RNO_1_3_LC_14_13_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst9.data_to_send_esr_RNO_1_3_LC_14_13_6 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \b2v_inst9.data_to_send_esr_RNO_1_3_LC_14_13_6  (
            .in0(N__24524),
            .in1(N__34556),
            .in2(N__24477),
            .in3(N__24880),
            .lcout(\b2v_inst9.data_to_send_10_0_0_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.pix_data_reg_RNIH87G_0_LC_14_14_0 .C_ON=1'b1;
    defparam \b2v_inst.pix_data_reg_RNIH87G_0_LC_14_14_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.pix_data_reg_RNIH87G_0_LC_14_14_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \b2v_inst.pix_data_reg_RNIH87G_0_LC_14_14_0  (
            .in0(_gnd_net_),
            .in1(N__25577),
            .in2(N__24421),
            .in3(_gnd_net_),
            .lcout(\b2v_inst.un14_data_ram_energia_o_axb_0 ),
            .ltout(),
            .carryin(bfn_14_14_0_),
            .carryout(\b2v_inst.un14_data_ram_energia_o_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un14_data_ram_energia_o_cry_0_c_RNIEI4M_LC_14_14_1 .C_ON=1'b1;
    defparam \b2v_inst.un14_data_ram_energia_o_cry_0_c_RNIEI4M_LC_14_14_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un14_data_ram_energia_o_cry_0_c_RNIEI4M_LC_14_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst.un14_data_ram_energia_o_cry_0_c_RNIEI4M_LC_14_14_1  (
            .in0(_gnd_net_),
            .in1(N__25571),
            .in2(N__24388),
            .in3(N__24356),
            .lcout(\b2v_inst.un14_data_ram_energia_o_cry_0_c_RNIEI4MZ0 ),
            .ltout(),
            .carryin(\b2v_inst.un14_data_ram_energia_o_cry_0 ),
            .carryout(\b2v_inst.un14_data_ram_energia_o_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un14_data_ram_energia_o_cry_1_c_RNIHM5M_LC_14_14_2 .C_ON=1'b1;
    defparam \b2v_inst.un14_data_ram_energia_o_cry_1_c_RNIHM5M_LC_14_14_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un14_data_ram_energia_o_cry_1_c_RNIHM5M_LC_14_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst.un14_data_ram_energia_o_cry_1_c_RNIHM5M_LC_14_14_2  (
            .in0(_gnd_net_),
            .in1(N__26300),
            .in2(N__24908),
            .in3(N__24884),
            .lcout(\b2v_inst.un14_data_ram_energia_o_cry_1_c_RNIHM5MZ0 ),
            .ltout(),
            .carryin(\b2v_inst.un14_data_ram_energia_o_cry_1 ),
            .carryout(\b2v_inst.un14_data_ram_energia_o_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un14_data_ram_energia_o_cry_2_c_RNIKQ6M_LC_14_14_3 .C_ON=1'b1;
    defparam \b2v_inst.un14_data_ram_energia_o_cry_2_c_RNIKQ6M_LC_14_14_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un14_data_ram_energia_o_cry_2_c_RNIKQ6M_LC_14_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst.un14_data_ram_energia_o_cry_2_c_RNIKQ6M_LC_14_14_3  (
            .in0(_gnd_net_),
            .in1(N__30260),
            .in2(N__24881),
            .in3(N__24857),
            .lcout(\b2v_inst.un14_data_ram_energia_o_cry_2_c_RNIKQ6MZ0 ),
            .ltout(),
            .carryin(\b2v_inst.un14_data_ram_energia_o_cry_2 ),
            .carryout(\b2v_inst.un14_data_ram_energia_o_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un14_data_ram_energia_o_cry_3_c_RNINU7M_LC_14_14_4 .C_ON=1'b1;
    defparam \b2v_inst.un14_data_ram_energia_o_cry_3_c_RNINU7M_LC_14_14_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un14_data_ram_energia_o_cry_3_c_RNINU7M_LC_14_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst.un14_data_ram_energia_o_cry_3_c_RNINU7M_LC_14_14_4  (
            .in0(_gnd_net_),
            .in1(N__24854),
            .in2(N__24836),
            .in3(N__24794),
            .lcout(\b2v_inst.un14_data_ram_energia_o_cry_3_c_RNINU7MZ0 ),
            .ltout(),
            .carryin(\b2v_inst.un14_data_ram_energia_o_cry_3 ),
            .carryout(\b2v_inst.un14_data_ram_energia_o_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un14_data_ram_energia_o_cry_4_c_RNIQ29M_LC_14_14_5 .C_ON=1'b1;
    defparam \b2v_inst.un14_data_ram_energia_o_cry_4_c_RNIQ29M_LC_14_14_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un14_data_ram_energia_o_cry_4_c_RNIQ29M_LC_14_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst.un14_data_ram_energia_o_cry_4_c_RNIQ29M_LC_14_14_5  (
            .in0(_gnd_net_),
            .in1(N__24790),
            .in2(N__26294),
            .in3(N__24767),
            .lcout(\b2v_inst.un14_data_ram_energia_o_cry_4_c_RNIQ29MZ0 ),
            .ltout(),
            .carryin(\b2v_inst.un14_data_ram_energia_o_cry_4 ),
            .carryout(\b2v_inst.un14_data_ram_energia_o_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un14_data_ram_energia_o_cry_5_c_RNIT6AM_LC_14_14_6 .C_ON=1'b1;
    defparam \b2v_inst.un14_data_ram_energia_o_cry_5_c_RNIT6AM_LC_14_14_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un14_data_ram_energia_o_cry_5_c_RNIT6AM_LC_14_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst.un14_data_ram_energia_o_cry_5_c_RNIT6AM_LC_14_14_6  (
            .in0(_gnd_net_),
            .in1(N__26285),
            .in2(N__24763),
            .in3(N__24731),
            .lcout(\b2v_inst.un14_data_ram_energia_o_cry_5_c_RNIT6AMZ0 ),
            .ltout(),
            .carryin(\b2v_inst.un14_data_ram_energia_o_cry_5 ),
            .carryout(\b2v_inst.un14_data_ram_energia_o_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un14_data_ram_energia_o_cry_6_c_RNI0BBM_LC_14_14_7 .C_ON=1'b1;
    defparam \b2v_inst.un14_data_ram_energia_o_cry_6_c_RNI0BBM_LC_14_14_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un14_data_ram_energia_o_cry_6_c_RNI0BBM_LC_14_14_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst.un14_data_ram_energia_o_cry_6_c_RNI0BBM_LC_14_14_7  (
            .in0(_gnd_net_),
            .in1(N__26279),
            .in2(N__24727),
            .in3(N__24695),
            .lcout(\b2v_inst.un14_data_ram_energia_o_cry_6_c_RNI0BBMZ0 ),
            .ltout(),
            .carryin(\b2v_inst.un14_data_ram_energia_o_cry_6 ),
            .carryout(\b2v_inst.un14_data_ram_energia_o_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un14_data_ram_energia_o_cry_7_c_RNIN84C_LC_14_15_0 .C_ON=1'b1;
    defparam \b2v_inst.un14_data_ram_energia_o_cry_7_c_RNIN84C_LC_14_15_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un14_data_ram_energia_o_cry_7_c_RNIN84C_LC_14_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.un14_data_ram_energia_o_cry_7_c_RNIN84C_LC_14_15_0  (
            .in0(_gnd_net_),
            .in1(N__24943),
            .in2(_gnd_net_),
            .in3(N__24680),
            .lcout(\b2v_inst.un14_data_ram_energia_o_cry_7_c_RNIN84CZ0 ),
            .ltout(),
            .carryin(bfn_14_15_0_),
            .carryout(\b2v_inst.un14_data_ram_energia_o_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un14_data_ram_energia_o_cry_8_c_RNIPB5C_LC_14_15_1 .C_ON=1'b1;
    defparam \b2v_inst.un14_data_ram_energia_o_cry_8_c_RNIPB5C_LC_14_15_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un14_data_ram_energia_o_cry_8_c_RNIPB5C_LC_14_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.un14_data_ram_energia_o_cry_8_c_RNIPB5C_LC_14_15_1  (
            .in0(_gnd_net_),
            .in1(N__26221),
            .in2(_gnd_net_),
            .in3(N__24665),
            .lcout(\b2v_inst.un14_data_ram_energia_o_cry_8_c_RNIPB5CZ0 ),
            .ltout(),
            .carryin(\b2v_inst.un14_data_ram_energia_o_cry_8 ),
            .carryout(\b2v_inst.un14_data_ram_energia_o_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un14_data_ram_energia_o_cry_9_c_RNI28GB_LC_14_15_2 .C_ON=1'b1;
    defparam \b2v_inst.un14_data_ram_energia_o_cry_9_c_RNI28GB_LC_14_15_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un14_data_ram_energia_o_cry_9_c_RNI28GB_LC_14_15_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.un14_data_ram_energia_o_cry_9_c_RNI28GB_LC_14_15_2  (
            .in0(_gnd_net_),
            .in1(N__25141),
            .in2(_gnd_net_),
            .in3(N__25112),
            .lcout(\b2v_inst.un14_data_ram_energia_o_cry_9_c_RNI28GBZ0 ),
            .ltout(),
            .carryin(\b2v_inst.un14_data_ram_energia_o_cry_9 ),
            .carryout(\b2v_inst.un14_data_ram_energia_o_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un14_data_ram_energia_o_cry_10_c_RNIMOAH_LC_14_15_3 .C_ON=1'b1;
    defparam \b2v_inst.un14_data_ram_energia_o_cry_10_c_RNIMOAH_LC_14_15_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un14_data_ram_energia_o_cry_10_c_RNIMOAH_LC_14_15_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst.un14_data_ram_energia_o_cry_10_c_RNIMOAH_LC_14_15_3  (
            .in0(N__37460),
            .in1(N__25105),
            .in2(_gnd_net_),
            .in3(N__25064),
            .lcout(SYNTHESIZED_WIRE_13_11),
            .ltout(),
            .carryin(\b2v_inst.un14_data_ram_energia_o_cry_10 ),
            .carryout(\b2v_inst.un14_data_ram_energia_o_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un14_data_ram_energia_o_cry_11_c_RNIORBH_LC_14_15_4 .C_ON=1'b1;
    defparam \b2v_inst.un14_data_ram_energia_o_cry_11_c_RNIORBH_LC_14_15_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un14_data_ram_energia_o_cry_11_c_RNIORBH_LC_14_15_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst.un14_data_ram_energia_o_cry_11_c_RNIORBH_LC_14_15_4  (
            .in0(N__37459),
            .in1(N__25057),
            .in2(_gnd_net_),
            .in3(N__25016),
            .lcout(SYNTHESIZED_WIRE_13_12),
            .ltout(),
            .carryin(\b2v_inst.un14_data_ram_energia_o_cry_11 ),
            .carryout(\b2v_inst.un14_data_ram_energia_o_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un14_data_ram_energia_o_cry_12_c_RNIQUCH_LC_14_15_5 .C_ON=1'b0;
    defparam \b2v_inst.un14_data_ram_energia_o_cry_12_c_RNIQUCH_LC_14_15_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un14_data_ram_energia_o_cry_12_c_RNIQUCH_LC_14_15_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst.un14_data_ram_energia_o_cry_12_c_RNIQUCH_LC_14_15_5  (
            .in0(N__37461),
            .in1(N__25009),
            .in2(_gnd_net_),
            .in3(N__24995),
            .lcout(SYNTHESIZED_WIRE_13_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.energia_temp_8_LC_14_15_6 .C_ON=1'b0;
    defparam \b2v_inst.energia_temp_8_LC_14_15_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.energia_temp_8_LC_14_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.energia_temp_8_LC_14_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24976),
            .lcout(b2v_inst_energia_temp_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34444),
            .ce(N__26190),
            .sr(N__38109));
    defparam \b2v_inst.data_a_escribir_RNIRV031_10_LC_14_16_0 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNIRV031_10_LC_14_16_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNIRV031_10_LC_14_16_0 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \b2v_inst.data_a_escribir_RNIRV031_10_LC_14_16_0  (
            .in0(N__37733),
            .in1(N__24932),
            .in2(N__33682),
            .in3(N__37502),
            .lcout(N_461_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.reg_ancho_2_5_LC_15_5_3 .C_ON=1'b0;
    defparam \b2v_inst.reg_ancho_2_5_LC_15_5_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_ancho_2_5_LC_15_5_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.reg_ancho_2_5_LC_15_5_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32124),
            .lcout(\b2v_inst.reg_ancho_2Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34449),
            .ce(N__32964),
            .sr(N__38115));
    defparam \b2v_inst.reg_anterior_2_LC_15_6_3 .C_ON=1'b0;
    defparam \b2v_inst.reg_anterior_2_LC_15_6_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_anterior_2_LC_15_6_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \b2v_inst.reg_anterior_2_LC_15_6_3  (
            .in0(_gnd_net_),
            .in1(N__31894),
            .in2(_gnd_net_),
            .in3(N__32210),
            .lcout(\b2v_inst.reg_anteriorZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34445),
            .ce(N__31686),
            .sr(N__38110));
    defparam \b2v_inst.reg_anterior_3_LC_15_6_4 .C_ON=1'b0;
    defparam \b2v_inst.reg_anterior_3_LC_15_6_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_anterior_3_LC_15_6_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \b2v_inst.reg_anterior_3_LC_15_6_4  (
            .in0(N__31895),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32285),
            .lcout(\b2v_inst.reg_anteriorZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34445),
            .ce(N__31686),
            .sr(N__38110));
    defparam \b2v_inst.data_a_escribir11_2_c_RNO_LC_15_7_0 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir11_2_c_RNO_LC_15_7_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir11_2_c_RNO_LC_15_7_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst.data_a_escribir11_2_c_RNO_LC_15_7_0  (
            .in0(N__29246),
            .in1(N__29988),
            .in2(N__27441),
            .in3(N__29949),
            .lcout(\b2v_inst.data_a_escribir11_2_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.reg_ancho_2_8_LC_15_7_3 .C_ON=1'b0;
    defparam \b2v_inst.reg_ancho_2_8_LC_15_7_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_ancho_2_8_LC_15_7_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.reg_ancho_2_8_LC_15_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27251),
            .lcout(\b2v_inst.reg_ancho_2Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34433),
            .ce(N__32930),
            .sr(N__38105));
    defparam \b2v_inst.data_a_escribir11_4_c_RNO_LC_15_7_4 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir11_4_c_RNO_LC_15_7_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir11_4_c_RNO_LC_15_7_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst.data_a_escribir11_4_c_RNO_LC_15_7_4  (
            .in0(N__27562),
            .in1(N__27319),
            .in2(N__29909),
            .in3(N__27383),
            .lcout(\b2v_inst.data_a_escribir11_4_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.reg_ancho_2_6_LC_15_7_6 .C_ON=1'b0;
    defparam \b2v_inst.reg_ancho_2_6_LC_15_7_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_ancho_2_6_LC_15_7_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.reg_ancho_2_6_LC_15_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31571),
            .lcout(\b2v_inst.reg_ancho_2Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34433),
            .ce(N__32930),
            .sr(N__38105));
    defparam \b2v_inst.reg_ancho_2_7_LC_15_7_7 .C_ON=1'b0;
    defparam \b2v_inst.reg_ancho_2_7_LC_15_7_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_ancho_2_7_LC_15_7_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.reg_ancho_2_7_LC_15_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27276),
            .lcout(\b2v_inst.reg_ancho_2Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34433),
            .ce(N__32930),
            .sr(N__38105));
    defparam \b2v_inst.data_a_escribir11_0_c_LC_15_8_0 .C_ON=1'b1;
    defparam \b2v_inst.data_a_escribir11_0_c_LC_15_8_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir11_0_c_LC_15_8_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.data_a_escribir11_0_c_LC_15_8_0  (
            .in0(_gnd_net_),
            .in1(N__26408),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_8_0_),
            .carryout(\b2v_inst.data_a_escribir11_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir11_1_c_LC_15_8_1 .C_ON=1'b1;
    defparam \b2v_inst.data_a_escribir11_1_c_LC_15_8_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir11_1_c_LC_15_8_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.data_a_escribir11_1_c_LC_15_8_1  (
            .in0(_gnd_net_),
            .in1(N__26630),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.data_a_escribir11_0 ),
            .carryout(\b2v_inst.data_a_escribir11_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir11_2_c_LC_15_8_2 .C_ON=1'b1;
    defparam \b2v_inst.data_a_escribir11_2_c_LC_15_8_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir11_2_c_LC_15_8_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.data_a_escribir11_2_c_LC_15_8_2  (
            .in0(_gnd_net_),
            .in1(N__25151),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.data_a_escribir11_1 ),
            .carryout(\b2v_inst.data_a_escribir11_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir11_3_c_LC_15_8_3 .C_ON=1'b1;
    defparam \b2v_inst.data_a_escribir11_3_c_LC_15_8_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir11_3_c_LC_15_8_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.data_a_escribir11_3_c_LC_15_8_3  (
            .in0(_gnd_net_),
            .in1(N__31415),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.data_a_escribir11_2 ),
            .carryout(\b2v_inst.data_a_escribir11_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir11_4_c_LC_15_8_4 .C_ON=1'b1;
    defparam \b2v_inst.data_a_escribir11_4_c_LC_15_8_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir11_4_c_LC_15_8_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.data_a_escribir11_4_c_LC_15_8_4  (
            .in0(_gnd_net_),
            .in1(N__25166),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.data_a_escribir11_3 ),
            .carryout(\b2v_inst.data_a_escribir11_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir11_5_c_LC_15_8_5 .C_ON=1'b1;
    defparam \b2v_inst.data_a_escribir11_5_c_LC_15_8_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir11_5_c_LC_15_8_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.data_a_escribir11_5_c_LC_15_8_5  (
            .in0(_gnd_net_),
            .in1(N__29648),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.data_a_escribir11_4 ),
            .carryout(\b2v_inst.data_a_escribir11_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir11_6_c_LC_15_8_6 .C_ON=1'b1;
    defparam \b2v_inst.data_a_escribir11_6_c_LC_15_8_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir11_6_c_LC_15_8_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.data_a_escribir11_6_c_LC_15_8_6  (
            .in0(_gnd_net_),
            .in1(N__29801),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.data_a_escribir11_5 ),
            .carryout(\b2v_inst.data_a_escribir11_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir11_7_c_LC_15_8_7 .C_ON=1'b1;
    defparam \b2v_inst.data_a_escribir11_7_c_LC_15_8_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir11_7_c_LC_15_8_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.data_a_escribir11_7_c_LC_15_8_7  (
            .in0(_gnd_net_),
            .in1(N__27296),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.data_a_escribir11_6 ),
            .carryout(\b2v_inst.data_a_escribir11_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir11_8_c_LC_15_9_0 .C_ON=1'b1;
    defparam \b2v_inst.data_a_escribir11_8_c_LC_15_9_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir11_8_c_LC_15_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.data_a_escribir11_8_c_LC_15_9_0  (
            .in0(_gnd_net_),
            .in1(N__25388),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_9_0_),
            .carryout(\b2v_inst.data_a_escribir11_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir11_9_c_LC_15_9_1 .C_ON=1'b1;
    defparam \b2v_inst.data_a_escribir11_9_c_LC_15_9_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir11_9_c_LC_15_9_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.data_a_escribir11_9_c_LC_15_9_1  (
            .in0(_gnd_net_),
            .in1(N__25157),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.data_a_escribir11_8 ),
            .carryout(\b2v_inst.data_a_escribir11_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir11_10_c_LC_15_9_2 .C_ON=1'b1;
    defparam \b2v_inst.data_a_escribir11_10_c_LC_15_9_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir11_10_c_LC_15_9_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.data_a_escribir11_10_c_LC_15_9_2  (
            .in0(_gnd_net_),
            .in1(N__30050),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.data_a_escribir11_9 ),
            .carryout(\b2v_inst.data_a_escribir12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir12_THRU_LUT4_0_LC_15_9_3 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir12_THRU_LUT4_0_LC_15_9_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir12_THRU_LUT4_0_LC_15_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.data_a_escribir12_THRU_LUT4_0_LC_15_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25160),
            .lcout(\b2v_inst.data_a_escribir12_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir11_9_c_RNO_LC_15_9_4 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir11_9_c_RNO_LC_15_9_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir11_9_c_RNO_LC_15_9_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst.data_a_escribir11_9_c_RNO_LC_15_9_4  (
            .in0(N__29105),
            .in1(N__30175),
            .in2(N__31529),
            .in3(N__29157),
            .lcout(\b2v_inst.data_a_escribir11_9_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir11_8_c_RNO_LC_15_9_5 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir11_8_c_RNO_LC_15_9_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir11_8_c_RNO_LC_15_9_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst.data_a_escribir11_8_c_RNO_LC_15_9_5  (
            .in0(N__28588),
            .in1(N__28614),
            .in2(N__29840),
            .in3(N__32309),
            .lcout(\b2v_inst.data_a_escribir11_8_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_3_RNI68I31_10_LC_15_9_7 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_3_RNI68I31_10_LC_15_9_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_3_RNI68I31_10_LC_15_9_7 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \b2v_inst.dir_mem_3_RNI68I31_10_LC_15_9_7  (
            .in0(N__25382),
            .in1(N__25367),
            .in2(N__25286),
            .in3(N__25268),
            .lcout(\b2v_inst.addr_ram_iv_i_1_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.eventos_0_LC_15_10_0 .C_ON=1'b1;
    defparam \b2v_inst.eventos_0_LC_15_10_0 .SEQ_MODE=4'b1011;
    defparam \b2v_inst.eventos_0_LC_15_10_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.eventos_0_LC_15_10_0  (
            .in0(_gnd_net_),
            .in1(N__26590),
            .in2(_gnd_net_),
            .in3(N__25187),
            .lcout(\b2v_inst.eventosZ0Z_0 ),
            .ltout(),
            .carryin(bfn_15_10_0_),
            .carryout(\b2v_inst.eventos_cry_0 ),
            .clk(N__34405),
            .ce(N__26651),
            .sr(N__38080));
    defparam \b2v_inst.eventos_1_LC_15_10_1 .C_ON=1'b1;
    defparam \b2v_inst.eventos_1_LC_15_10_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.eventos_1_LC_15_10_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.eventos_1_LC_15_10_1  (
            .in0(_gnd_net_),
            .in1(N__26569),
            .in2(_gnd_net_),
            .in3(N__25184),
            .lcout(\b2v_inst.eventosZ0Z_1 ),
            .ltout(),
            .carryin(\b2v_inst.eventos_cry_0 ),
            .carryout(\b2v_inst.eventos_cry_1 ),
            .clk(N__34405),
            .ce(N__26651),
            .sr(N__38080));
    defparam \b2v_inst.eventos_2_LC_15_10_2 .C_ON=1'b1;
    defparam \b2v_inst.eventos_2_LC_15_10_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.eventos_2_LC_15_10_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.eventos_2_LC_15_10_2  (
            .in0(_gnd_net_),
            .in1(N__31195),
            .in2(_gnd_net_),
            .in3(N__25181),
            .lcout(\b2v_inst.eventosZ0Z_2 ),
            .ltout(),
            .carryin(\b2v_inst.eventos_cry_1 ),
            .carryout(\b2v_inst.eventos_cry_2 ),
            .clk(N__34405),
            .ce(N__26651),
            .sr(N__38080));
    defparam \b2v_inst.eventos_3_LC_15_10_3 .C_ON=1'b1;
    defparam \b2v_inst.eventos_3_LC_15_10_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.eventos_3_LC_15_10_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.eventos_3_LC_15_10_3  (
            .in0(_gnd_net_),
            .in1(N__29863),
            .in2(_gnd_net_),
            .in3(N__25178),
            .lcout(\b2v_inst.eventosZ0Z_3 ),
            .ltout(),
            .carryin(\b2v_inst.eventos_cry_2 ),
            .carryout(\b2v_inst.eventos_cry_3 ),
            .clk(N__34405),
            .ce(N__26651),
            .sr(N__38080));
    defparam \b2v_inst.eventos_4_LC_15_10_4 .C_ON=1'b1;
    defparam \b2v_inst.eventos_4_LC_15_10_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.eventos_4_LC_15_10_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.eventos_4_LC_15_10_4  (
            .in0(_gnd_net_),
            .in1(N__26617),
            .in2(_gnd_net_),
            .in3(N__25175),
            .lcout(\b2v_inst.eventosZ0Z_4 ),
            .ltout(),
            .carryin(\b2v_inst.eventos_cry_3 ),
            .carryout(\b2v_inst.eventos_cry_4 ),
            .clk(N__34405),
            .ce(N__26651),
            .sr(N__38080));
    defparam \b2v_inst.eventos_5_LC_15_10_5 .C_ON=1'b1;
    defparam \b2v_inst.eventos_5_LC_15_10_5 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.eventos_5_LC_15_10_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.eventos_5_LC_15_10_5  (
            .in0(_gnd_net_),
            .in1(N__27520),
            .in2(_gnd_net_),
            .in3(N__25172),
            .lcout(\b2v_inst.eventosZ0Z_5 ),
            .ltout(),
            .carryin(\b2v_inst.eventos_cry_4 ),
            .carryout(\b2v_inst.eventos_cry_5 ),
            .clk(N__34405),
            .ce(N__26651),
            .sr(N__38080));
    defparam \b2v_inst.eventos_6_LC_15_10_6 .C_ON=1'b1;
    defparam \b2v_inst.eventos_6_LC_15_10_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.eventos_6_LC_15_10_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.eventos_6_LC_15_10_6  (
            .in0(_gnd_net_),
            .in1(N__26674),
            .in2(_gnd_net_),
            .in3(N__25169),
            .lcout(\b2v_inst.eventosZ0Z_6 ),
            .ltout(),
            .carryin(\b2v_inst.eventos_cry_5 ),
            .carryout(\b2v_inst.eventos_cry_6 ),
            .clk(N__34405),
            .ce(N__26651),
            .sr(N__38080));
    defparam \b2v_inst.eventos_7_LC_15_10_7 .C_ON=1'b1;
    defparam \b2v_inst.eventos_7_LC_15_10_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.eventos_7_LC_15_10_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.eventos_7_LC_15_10_7  (
            .in0(_gnd_net_),
            .in1(N__28480),
            .in2(_gnd_net_),
            .in3(N__25565),
            .lcout(\b2v_inst.eventosZ0Z_7 ),
            .ltout(),
            .carryin(\b2v_inst.eventos_cry_6 ),
            .carryout(\b2v_inst.eventos_cry_7 ),
            .clk(N__34405),
            .ce(N__26651),
            .sr(N__38080));
    defparam \b2v_inst.eventos_8_LC_15_11_0 .C_ON=1'b1;
    defparam \b2v_inst.eventos_8_LC_15_11_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.eventos_8_LC_15_11_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.eventos_8_LC_15_11_0  (
            .in0(_gnd_net_),
            .in1(N__30034),
            .in2(_gnd_net_),
            .in3(N__25562),
            .lcout(\b2v_inst.eventosZ0Z_8 ),
            .ltout(),
            .carryin(bfn_15_11_0_),
            .carryout(\b2v_inst.eventos_cry_8 ),
            .clk(N__34394),
            .ce(N__26647),
            .sr(N__38093));
    defparam \b2v_inst.eventos_9_LC_15_11_1 .C_ON=1'b1;
    defparam \b2v_inst.eventos_9_LC_15_11_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.eventos_9_LC_15_11_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.eventos_9_LC_15_11_1  (
            .in0(_gnd_net_),
            .in1(N__30109),
            .in2(_gnd_net_),
            .in3(N__25559),
            .lcout(\b2v_inst.eventosZ0Z_9 ),
            .ltout(),
            .carryin(\b2v_inst.eventos_cry_8 ),
            .carryout(\b2v_inst.eventos_cry_9 ),
            .clk(N__34394),
            .ce(N__26647),
            .sr(N__38093));
    defparam \b2v_inst.eventos_10_LC_15_11_2 .C_ON=1'b0;
    defparam \b2v_inst.eventos_10_LC_15_11_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.eventos_10_LC_15_11_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \b2v_inst.eventos_10_LC_15_11_2  (
            .in0(_gnd_net_),
            .in1(N__26552),
            .in2(_gnd_net_),
            .in3(N__25556),
            .lcout(\b2v_inst.eventosZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34394),
            .ce(N__26647),
            .sr(N__38093));
    defparam \b2v_inst.state_RNO_1_31_LC_15_12_0 .C_ON=1'b0;
    defparam \b2v_inst.state_RNO_1_31_LC_15_12_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNO_1_31_LC_15_12_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst.state_RNO_1_31_LC_15_12_0  (
            .in0(N__25417),
            .in1(N__25470),
            .in2(N__34746),
            .in3(N__28064),
            .lcout(),
            .ltout(\b2v_inst.state_ns_a3_i_0_a2_4_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_31_LC_15_12_1 .C_ON=1'b0;
    defparam \b2v_inst.state_31_LC_15_12_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.state_31_LC_15_12_1 .LUT_INIT=16'b0000000001111111;
    LogicCell40 \b2v_inst.state_31_LC_15_12_1  (
            .in0(N__25784),
            .in1(N__25553),
            .in2(N__25541),
            .in3(N__28016),
            .lcout(\b2v_inst.stateZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34406),
            .ce(),
            .sr(N__38102));
    defparam \b2v_inst.state_RNO_6_31_LC_15_12_3 .C_ON=1'b0;
    defparam \b2v_inst.state_RNO_6_31_LC_15_12_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNO_6_31_LC_15_12_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst.state_RNO_6_31_LC_15_12_3  (
            .in0(N__25469),
            .in1(N__25416),
            .in2(N__25731),
            .in3(N__25814),
            .lcout(\b2v_inst.state_ns_a3_i_0_a2_1_4_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_1_LC_15_12_4 .C_ON=1'b0;
    defparam \b2v_inst.state_1_LC_15_12_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.state_1_LC_15_12_4 .LUT_INIT=16'b1111111110100000;
    LogicCell40 \b2v_inst.state_1_LC_15_12_4  (
            .in0(N__25418),
            .in1(_gnd_net_),
            .in2(N__30412),
            .in3(N__26061),
            .lcout(b2v_inst_state_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34406),
            .ce(),
            .sr(N__38102));
    defparam \b2v_inst.state_12_LC_15_12_5 .C_ON=1'b0;
    defparam \b2v_inst.state_12_LC_15_12_5 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.state_12_LC_15_12_5 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \b2v_inst.state_12_LC_15_12_5  (
            .in0(N__25722),
            .in1(N__30379),
            .in2(_gnd_net_),
            .in3(N__25691),
            .lcout(b2v_inst_state_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34406),
            .ce(),
            .sr(N__38102));
    defparam \b2v_inst.state_2_LC_15_12_6 .C_ON=1'b0;
    defparam \b2v_inst.state_2_LC_15_12_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.state_2_LC_15_12_6 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \b2v_inst.state_2_LC_15_12_6  (
            .in0(N__30383),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28065),
            .lcout(b2v_inst_state_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34406),
            .ce(),
            .sr(N__38102));
    defparam \b2v_inst.state_11_LC_15_12_7 .C_ON=1'b0;
    defparam \b2v_inst.state_11_LC_15_12_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.state_11_LC_15_12_7 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \b2v_inst.state_11_LC_15_12_7  (
            .in0(N__25721),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30378),
            .lcout(\b2v_inst.stateZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34406),
            .ce(),
            .sr(N__38102));
    defparam \b2v_inst.state_RNO_3_31_LC_15_13_0 .C_ON=1'b0;
    defparam \b2v_inst.state_RNO_3_31_LC_15_13_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNO_3_31_LC_15_13_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst.state_RNO_3_31_LC_15_13_0  (
            .in0(N__25724),
            .in1(N__33180),
            .in2(N__25935),
            .in3(N__25817),
            .lcout(\b2v_inst.state_ns_a3_i_0_a2_6_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst9.fsm_state_RNO_0_1_LC_15_13_4 .C_ON=1'b0;
    defparam \b2v_inst9.fsm_state_RNO_0_1_LC_15_13_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst9.fsm_state_RNO_0_1_LC_15_13_4 .LUT_INIT=16'b0010001000110011;
    LogicCell40 \b2v_inst9.fsm_state_RNO_0_1_LC_15_13_4  (
            .in0(N__30472),
            .in1(N__27162),
            .in2(_gnd_net_),
            .in3(N__26884),
            .lcout(),
            .ltout(\b2v_inst9.fsm_state_ns_i_0_i_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst9.fsm_state_1_LC_15_13_5 .C_ON=1'b0;
    defparam \b2v_inst9.fsm_state_1_LC_15_13_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst9.fsm_state_1_LC_15_13_5 .LUT_INIT=16'b0000010000001100;
    LogicCell40 \b2v_inst9.fsm_state_1_LC_15_13_5  (
            .in0(N__26885),
            .in1(N__27840),
            .in2(N__25778),
            .in3(N__27101),
            .lcout(\b2v_inst9.fsm_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34413),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst9.data_to_send_esr_RNO_0_2_LC_15_13_6 .C_ON=1'b0;
    defparam \b2v_inst9.data_to_send_esr_RNO_0_2_LC_15_13_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst9.data_to_send_esr_RNO_0_2_LC_15_13_6 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \b2v_inst9.data_to_send_esr_RNO_0_2_LC_15_13_6  (
            .in0(N__25775),
            .in1(N__33648),
            .in2(N__25763),
            .in3(N__30375),
            .lcout(\b2v_inst9.data_to_send_10_0_0_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst9.fsm_state_RNIS2UL_0_LC_15_13_7 .C_ON=1'b0;
    defparam \b2v_inst9.fsm_state_RNIS2UL_0_LC_15_13_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst9.fsm_state_RNIS2UL_0_LC_15_13_7 .LUT_INIT=16'b0000010100000100;
    LogicCell40 \b2v_inst9.fsm_state_RNIS2UL_0_LC_15_13_7  (
            .in0(N__26883),
            .in1(N__25723),
            .in2(N__27188),
            .in3(N__25687),
            .lcout(\b2v_inst9.N_739 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.pix_data_reg_0_LC_15_14_0 .C_ON=1'b0;
    defparam \b2v_inst.pix_data_reg_0_LC_15_14_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.pix_data_reg_0_LC_15_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.pix_data_reg_0_LC_15_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26690),
            .lcout(\b2v_inst.pix_data_regZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34424),
            .ce(N__30244),
            .sr(N__38111));
    defparam \b2v_inst.pix_data_reg_1_LC_15_14_1 .C_ON=1'b0;
    defparam \b2v_inst.pix_data_reg_1_LC_15_14_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.pix_data_reg_1_LC_15_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.pix_data_reg_1_LC_15_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26999),
            .lcout(\b2v_inst.pix_data_regZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34424),
            .ce(N__30244),
            .sr(N__38111));
    defparam \b2v_inst.pix_data_reg_2_LC_15_14_2 .C_ON=1'b0;
    defparam \b2v_inst.pix_data_reg_2_LC_15_14_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.pix_data_reg_2_LC_15_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.pix_data_reg_2_LC_15_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26966),
            .lcout(\b2v_inst.pix_data_regZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34424),
            .ce(N__30244),
            .sr(N__38111));
    defparam \b2v_inst.pix_data_reg_5_LC_15_14_4 .C_ON=1'b0;
    defparam \b2v_inst.pix_data_reg_5_LC_15_14_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.pix_data_reg_5_LC_15_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.pix_data_reg_5_LC_15_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28802),
            .lcout(\b2v_inst.pix_data_regZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34424),
            .ce(N__30244),
            .sr(N__38111));
    defparam \b2v_inst.pix_data_reg_6_LC_15_14_6 .C_ON=1'b0;
    defparam \b2v_inst.pix_data_reg_6_LC_15_14_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.pix_data_reg_6_LC_15_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.pix_data_reg_6_LC_15_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28841),
            .lcout(\b2v_inst.pix_data_regZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34424),
            .ce(N__30244),
            .sr(N__38111));
    defparam \b2v_inst.pix_data_reg_7_LC_15_14_7 .C_ON=1'b0;
    defparam \b2v_inst.pix_data_reg_7_LC_15_14_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.pix_data_reg_7_LC_15_14_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst.pix_data_reg_7_LC_15_14_7  (
            .in0(N__28853),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst.pix_data_regZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34424),
            .ce(N__30244),
            .sr(N__38111));
    defparam \b2v_inst9.fsm_state_0_LC_15_15_3 .C_ON=1'b0;
    defparam \b2v_inst9.fsm_state_0_LC_15_15_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst9.fsm_state_0_LC_15_15_3 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \b2v_inst9.fsm_state_0_LC_15_15_3  (
            .in0(N__26921),
            .in1(N__26273),
            .in2(N__27845),
            .in3(N__27097),
            .lcout(\b2v_inst9.fsm_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34434),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.energia_temp_9_LC_15_17_5 .C_ON=1'b0;
    defparam \b2v_inst.energia_temp_9_LC_15_17_5 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.energia_temp_9_LC_15_17_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.energia_temp_9_LC_15_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26260),
            .lcout(b2v_inst_energia_temp_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34450),
            .ce(N__26205),
            .sr(N__38128));
    defparam \b2v_inst9.txd_reg_LC_15_18_2 .C_ON=1'b0;
    defparam \b2v_inst9.txd_reg_LC_15_18_2 .SEQ_MODE=4'b1001;
    defparam \b2v_inst9.txd_reg_LC_15_18_2 .LUT_INIT=16'b1100110010111011;
    LogicCell40 \b2v_inst9.txd_reg_LC_15_18_2  (
            .in0(N__26111),
            .in1(N__27192),
            .in2(_gnd_net_),
            .in3(N__26898),
            .lcout(uart_tx_o_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34457),
            .ce(),
            .sr(N__38135));
    defparam \b2v_inst.reg_ancho_2_0_LC_16_4_2 .C_ON=1'b0;
    defparam \b2v_inst.reg_ancho_2_0_LC_16_4_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_ancho_2_0_LC_16_4_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst.reg_ancho_2_0_LC_16_4_2  (
            .in0(N__27486),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst.reg_ancho_2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34451),
            .ce(N__32958),
            .sr(N__38129));
    defparam \b2v_inst.reg_ancho_1_0_LC_16_5_0 .C_ON=1'b0;
    defparam \b2v_inst.reg_ancho_1_0_LC_16_5_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_ancho_1_0_LC_16_5_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \b2v_inst.reg_ancho_1_0_LC_16_5_0  (
            .in0(_gnd_net_),
            .in1(N__26522),
            .in2(_gnd_net_),
            .in3(N__27479),
            .lcout(\b2v_inst.reg_ancho_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34446),
            .ce(N__26462),
            .sr(N__38123));
    defparam \b2v_inst.reg_ancho_1_1_LC_16_5_1 .C_ON=1'b0;
    defparam \b2v_inst.reg_ancho_1_1_LC_16_5_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_ancho_1_1_LC_16_5_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \b2v_inst.reg_ancho_1_1_LC_16_5_1  (
            .in0(N__26524),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31394),
            .lcout(\b2v_inst.reg_ancho_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34446),
            .ce(N__26462),
            .sr(N__38123));
    defparam \b2v_inst.reg_ancho_1_10_LC_16_5_2 .C_ON=1'b0;
    defparam \b2v_inst.reg_ancho_1_10_LC_16_5_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_ancho_1_10_LC_16_5_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \b2v_inst.reg_ancho_1_10_LC_16_5_2  (
            .in0(_gnd_net_),
            .in1(N__26523),
            .in2(_gnd_net_),
            .in3(N__31781),
            .lcout(\b2v_inst.reg_ancho_1Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34446),
            .ce(N__26462),
            .sr(N__38123));
    defparam \b2v_inst.reg_ancho_1_2_LC_16_5_3 .C_ON=1'b0;
    defparam \b2v_inst.reg_ancho_1_2_LC_16_5_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_ancho_1_2_LC_16_5_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \b2v_inst.reg_ancho_1_2_LC_16_5_3  (
            .in0(N__26525),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32204),
            .lcout(\b2v_inst.reg_ancho_1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34446),
            .ce(N__26462),
            .sr(N__38123));
    defparam \b2v_inst.reg_ancho_1_3_LC_16_5_4 .C_ON=1'b0;
    defparam \b2v_inst.reg_ancho_1_3_LC_16_5_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_ancho_1_3_LC_16_5_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \b2v_inst.reg_ancho_1_3_LC_16_5_4  (
            .in0(_gnd_net_),
            .in1(N__26526),
            .in2(_gnd_net_),
            .in3(N__32282),
            .lcout(\b2v_inst.reg_ancho_1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34446),
            .ce(N__26462),
            .sr(N__38123));
    defparam \b2v_inst.reg_ancho_1_4_LC_16_5_5 .C_ON=1'b0;
    defparam \b2v_inst.reg_ancho_1_4_LC_16_5_5 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_ancho_1_4_LC_16_5_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \b2v_inst.reg_ancho_1_4_LC_16_5_5  (
            .in0(N__26527),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33062),
            .lcout(\b2v_inst.reg_ancho_1Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34446),
            .ce(N__26462),
            .sr(N__38123));
    defparam \b2v_inst.reg_ancho_1_6_LC_16_5_7 .C_ON=1'b0;
    defparam \b2v_inst.reg_ancho_1_6_LC_16_5_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_ancho_1_6_LC_16_5_7 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \b2v_inst.reg_ancho_1_6_LC_16_5_7  (
            .in0(N__26528),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31570),
            .lcout(\b2v_inst.reg_ancho_1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34446),
            .ce(N__26462),
            .sr(N__38123));
    defparam \b2v_inst.encontrar_maximo_un2_valor_max1_cry_0_c_inv_LC_16_6_0 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_un2_valor_max1_cry_0_c_inv_LC_16_6_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_un2_valor_max1_cry_0_c_inv_LC_16_6_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst.encontrar_maximo_un2_valor_max1_cry_0_c_inv_LC_16_6_0  (
            .in0(_gnd_net_),
            .in1(N__27430),
            .in2(N__26327),
            .in3(N__29045),
            .lcout(\b2v_inst.reg_ancho_1_i_0 ),
            .ltout(),
            .carryin(bfn_16_6_0_),
            .carryout(\b2v_inst.un2_valor_max1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_un2_valor_max1_cry_1_c_inv_LC_16_6_1 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_un2_valor_max1_cry_1_c_inv_LC_16_6_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_un2_valor_max1_cry_1_c_inv_LC_16_6_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst.encontrar_maximo_un2_valor_max1_cry_1_c_inv_LC_16_6_1  (
            .in0(_gnd_net_),
            .in1(N__31346),
            .in2(N__26318),
            .in3(N__28971),
            .lcout(\b2v_inst.reg_ancho_1_i_1 ),
            .ltout(),
            .carryin(\b2v_inst.un2_valor_max1_cry_0 ),
            .carryout(\b2v_inst.un2_valor_max1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_un2_valor_max1_cry_2_c_inv_LC_16_6_2 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_un2_valor_max1_cry_2_c_inv_LC_16_6_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_un2_valor_max1_cry_2_c_inv_LC_16_6_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst.encontrar_maximo_un2_valor_max1_cry_2_c_inv_LC_16_6_2  (
            .in0(_gnd_net_),
            .in1(N__31299),
            .in2(N__26309),
            .in3(N__31223),
            .lcout(\b2v_inst.reg_ancho_1_i_2 ),
            .ltout(),
            .carryin(\b2v_inst.un2_valor_max1_cry_1 ),
            .carryout(\b2v_inst.un2_valor_max1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_un2_valor_max1_cry_3_c_inv_LC_16_6_3 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_un2_valor_max1_cry_3_c_inv_LC_16_6_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_un2_valor_max1_cry_3_c_inv_LC_16_6_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst.encontrar_maximo_un2_valor_max1_cry_3_c_inv_LC_16_6_3  (
            .in0(_gnd_net_),
            .in1(N__32448),
            .in2(N__26399),
            .in3(N__31010),
            .lcout(\b2v_inst.reg_ancho_1_i_3 ),
            .ltout(),
            .carryin(\b2v_inst.un2_valor_max1_cry_2 ),
            .carryout(\b2v_inst.un2_valor_max1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_un2_valor_max1_cry_4_c_inv_LC_16_6_4 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_un2_valor_max1_cry_4_c_inv_LC_16_6_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_un2_valor_max1_cry_4_c_inv_LC_16_6_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst.encontrar_maximo_un2_valor_max1_cry_4_c_inv_LC_16_6_4  (
            .in0(_gnd_net_),
            .in1(N__33015),
            .in2(N__26390),
            .in3(N__29615),
            .lcout(\b2v_inst.reg_ancho_1_i_4 ),
            .ltout(),
            .carryin(\b2v_inst.un2_valor_max1_cry_3 ),
            .carryout(\b2v_inst.un2_valor_max1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_un2_valor_max1_cry_5_c_inv_LC_16_6_5 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_un2_valor_max1_cry_5_c_inv_LC_16_6_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_un2_valor_max1_cry_5_c_inv_LC_16_6_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst.encontrar_maximo_un2_valor_max1_cry_5_c_inv_LC_16_6_5  (
            .in0(_gnd_net_),
            .in1(N__27370),
            .in2(N__26381),
            .in3(N__29551),
            .lcout(\b2v_inst.reg_ancho_1_i_5 ),
            .ltout(),
            .carryin(\b2v_inst.un2_valor_max1_cry_4 ),
            .carryout(\b2v_inst.un2_valor_max1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_un2_valor_max1_cry_6_c_inv_LC_16_6_6 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_un2_valor_max1_cry_6_c_inv_LC_16_6_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_un2_valor_max1_cry_6_c_inv_LC_16_6_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst.encontrar_maximo_un2_valor_max1_cry_6_c_inv_LC_16_6_6  (
            .in0(_gnd_net_),
            .in1(N__27320),
            .in2(N__26372),
            .in3(N__29465),
            .lcout(\b2v_inst.reg_ancho_1_i_6 ),
            .ltout(),
            .carryin(\b2v_inst.un2_valor_max1_cry_5 ),
            .carryout(\b2v_inst.un2_valor_max1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_un2_valor_max1_cry_7_c_inv_LC_16_6_7 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_un2_valor_max1_cry_7_c_inv_LC_16_6_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_un2_valor_max1_cry_7_c_inv_LC_16_6_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst.encontrar_maximo_un2_valor_max1_cry_7_c_inv_LC_16_6_7  (
            .in0(_gnd_net_),
            .in1(N__27575),
            .in2(N__26363),
            .in3(N__29386),
            .lcout(\b2v_inst.reg_ancho_1_i_7 ),
            .ltout(),
            .carryin(\b2v_inst.un2_valor_max1_cry_6 ),
            .carryout(\b2v_inst.un2_valor_max1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_un2_valor_max1_cry_8_c_inv_LC_16_7_0 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_un2_valor_max1_cry_8_c_inv_LC_16_7_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_un2_valor_max1_cry_8_c_inv_LC_16_7_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst.encontrar_maximo_un2_valor_max1_cry_8_c_inv_LC_16_7_0  (
            .in0(N__29948),
            .in1(N__29899),
            .in2(N__26354),
            .in3(_gnd_net_),
            .lcout(\b2v_inst.reg_ancho_1_i_8 ),
            .ltout(),
            .carryin(bfn_16_7_0_),
            .carryout(\b2v_inst.un2_valor_max1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_un2_valor_max1_cry_9_c_inv_LC_16_7_1 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_un2_valor_max1_cry_9_c_inv_LC_16_7_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_un2_valor_max1_cry_9_c_inv_LC_16_7_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst.encontrar_maximo_un2_valor_max1_cry_9_c_inv_LC_16_7_1  (
            .in0(_gnd_net_),
            .in1(N__29725),
            .in2(N__26345),
            .in3(N__29987),
            .lcout(\b2v_inst.reg_ancho_1_i_9 ),
            .ltout(),
            .carryin(\b2v_inst.un2_valor_max1_cry_8 ),
            .carryout(\b2v_inst.un2_valor_max1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_un2_valor_max1_cry_10_c_inv_LC_16_7_2 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_un2_valor_max1_cry_10_c_inv_LC_16_7_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_un2_valor_max1_cry_10_c_inv_LC_16_7_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst.encontrar_maximo_un2_valor_max1_cry_10_c_inv_LC_16_7_2  (
            .in0(_gnd_net_),
            .in1(N__31487),
            .in2(N__26336),
            .in3(N__29245),
            .lcout(\b2v_inst.reg_ancho_1_i_10 ),
            .ltout(),
            .carryin(\b2v_inst.un2_valor_max1_cry_9 ),
            .carryout(\b2v_inst.un2_valor_max1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un2_valor_max1_THRU_LUT4_0_LC_16_7_3 .C_ON=1'b0;
    defparam \b2v_inst.un2_valor_max1_THRU_LUT4_0_LC_16_7_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un2_valor_max1_THRU_LUT4_0_LC_16_7_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.un2_valor_max1_THRU_LUT4_0_LC_16_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26531),
            .lcout(\b2v_inst.un2_valor_max1_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.reg_ancho_2_9_LC_16_7_4 .C_ON=1'b0;
    defparam \b2v_inst.reg_ancho_2_9_LC_16_7_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_ancho_2_9_LC_16_7_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.reg_ancho_2_9_LC_16_7_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31994),
            .lcout(\b2v_inst.reg_ancho_2Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34425),
            .ce(N__32963),
            .sr(N__38112));
    defparam \b2v_inst.reg_ancho_1_7_LC_16_8_0 .C_ON=1'b0;
    defparam \b2v_inst.reg_ancho_1_7_LC_16_8_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_ancho_1_7_LC_16_8_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \b2v_inst.reg_ancho_1_7_LC_16_8_0  (
            .in0(N__26519),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27283),
            .lcout(\b2v_inst.reg_ancho_1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34414),
            .ce(N__26458),
            .sr(N__38106));
    defparam \b2v_inst.reg_ancho_1_8_LC_16_8_1 .C_ON=1'b0;
    defparam \b2v_inst.reg_ancho_1_8_LC_16_8_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_ancho_1_8_LC_16_8_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \b2v_inst.reg_ancho_1_8_LC_16_8_1  (
            .in0(_gnd_net_),
            .in1(N__26520),
            .in2(_gnd_net_),
            .in3(N__27249),
            .lcout(\b2v_inst.reg_ancho_1Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34414),
            .ce(N__26458),
            .sr(N__38106));
    defparam \b2v_inst.reg_ancho_1_9_LC_16_8_2 .C_ON=1'b0;
    defparam \b2v_inst.reg_ancho_1_9_LC_16_8_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_ancho_1_9_LC_16_8_2 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \b2v_inst.reg_ancho_1_9_LC_16_8_2  (
            .in0(N__31993),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26521),
            .lcout(\b2v_inst.reg_ancho_1Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34414),
            .ce(N__26458),
            .sr(N__38106));
    defparam \b2v_inst.reg_ancho_1_5_LC_16_8_3 .C_ON=1'b0;
    defparam \b2v_inst.reg_ancho_1_5_LC_16_8_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_ancho_1_5_LC_16_8_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \b2v_inst.reg_ancho_1_5_LC_16_8_3  (
            .in0(_gnd_net_),
            .in1(N__26518),
            .in2(_gnd_net_),
            .in3(N__32132),
            .lcout(\b2v_inst.reg_ancho_1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34414),
            .ce(N__26458),
            .sr(N__38106));
    defparam \b2v_inst.reg_anterior_0_LC_16_9_0 .C_ON=1'b0;
    defparam \b2v_inst.reg_anterior_0_LC_16_9_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_anterior_0_LC_16_9_0 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \b2v_inst.reg_anterior_0_LC_16_9_0  (
            .in0(N__27488),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31831),
            .lcout(\b2v_inst.reg_anteriorZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34407),
            .ce(N__31671),
            .sr(N__38103));
    defparam \b2v_inst.reg_anterior_8_LC_16_9_3 .C_ON=1'b0;
    defparam \b2v_inst.reg_anterior_8_LC_16_9_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_anterior_8_LC_16_9_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \b2v_inst.reg_anterior_8_LC_16_9_3  (
            .in0(_gnd_net_),
            .in1(N__31833),
            .in2(_gnd_net_),
            .in3(N__27248),
            .lcout(\b2v_inst.reg_anteriorZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34407),
            .ce(N__31671),
            .sr(N__38103));
    defparam \b2v_inst.reg_anterior_7_LC_16_9_6 .C_ON=1'b0;
    defparam \b2v_inst.reg_anterior_7_LC_16_9_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_anterior_7_LC_16_9_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \b2v_inst.reg_anterior_7_LC_16_9_6  (
            .in0(_gnd_net_),
            .in1(N__31832),
            .in2(_gnd_net_),
            .in3(N__27284),
            .lcout(\b2v_inst.reg_anteriorZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34407),
            .ce(N__31671),
            .sr(N__38103));
    defparam \b2v_inst.data_a_escribir11_0_c_RNO_LC_16_10_0 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir11_0_c_RNO_LC_16_10_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir11_0_c_RNO_LC_16_10_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst.data_a_escribir11_0_c_RNO_LC_16_10_0  (
            .in0(N__31241),
            .in1(N__28982),
            .in2(N__31042),
            .in3(N__29060),
            .lcout(\b2v_inst.data_a_escribir11_0_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_2_0_LC_16_10_1 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_2_0_LC_16_10_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_2_0_LC_16_10_1 .LUT_INIT=16'b0011111101011111;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_2_0_LC_16_10_1  (
            .in0(N__29061),
            .in1(N__27449),
            .in2(N__30910),
            .in3(N__32540),
            .lcout(),
            .ltout(\b2v_inst.data_a_escribir_RNO_2Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_1_0_LC_16_10_2 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_1_0_LC_16_10_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_1_0_LC_16_10_2 .LUT_INIT=16'b0111011100001111;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_1_0_LC_16_10_2  (
            .in0(N__26591),
            .in1(N__30860),
            .in2(N__26579),
            .in3(N__31110),
            .lcout(),
            .ltout(\b2v_inst.un1_reg_anterior_0_i_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_0_LC_16_10_3 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_0_LC_16_10_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.data_a_escribir_0_LC_16_10_3 .LUT_INIT=16'b0001101101011010;
    LogicCell40 \b2v_inst.data_a_escribir_0_LC_16_10_3  (
            .in0(N__31112),
            .in1(N__27539),
            .in2(N__26576),
            .in3(N__30625),
            .lcout(b2v_inst_data_a_escribir_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34395),
            .ce(N__30553),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_2_1_LC_16_10_5 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_2_1_LC_16_10_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_2_1_LC_16_10_5 .LUT_INIT=16'b0011111101011111;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_2_1_LC_16_10_5  (
            .in0(N__28983),
            .in1(N__31350),
            .in2(N__30911),
            .in3(N__32541),
            .lcout(),
            .ltout(\b2v_inst.data_a_escribir_RNO_2Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_1_1_LC_16_10_6 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_1_1_LC_16_10_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_1_1_LC_16_10_6 .LUT_INIT=16'b0111011100001111;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_1_1_LC_16_10_6  (
            .in0(N__26573),
            .in1(N__30861),
            .in2(N__26558),
            .in3(N__31111),
            .lcout(),
            .ltout(\b2v_inst.un1_reg_anterior_0_i_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_1_LC_16_10_7 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_1_LC_16_10_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.data_a_escribir_1_LC_16_10_7 .LUT_INIT=16'b0001101101011010;
    LogicCell40 \b2v_inst.data_a_escribir_1_LC_16_10_7  (
            .in0(N__31113),
            .in1(N__27533),
            .in2(N__26555),
            .in3(N__30626),
            .lcout(b2v_inst_data_a_escribir_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34395),
            .ce(N__30553),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_2_10_LC_16_11_0 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_2_10_LC_16_11_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_2_10_LC_16_11_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_2_10_LC_16_11_0  (
            .in0(N__29258),
            .in1(N__31490),
            .in2(_gnd_net_),
            .in3(N__32537),
            .lcout(\b2v_inst.N_269 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_3_10_LC_16_11_1 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_3_10_LC_16_11_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_3_10_LC_16_11_1 .LUT_INIT=16'b0011111100001111;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_3_10_LC_16_11_1  (
            .in0(_gnd_net_),
            .in1(N__26551),
            .in2(N__30982),
            .in3(N__31114),
            .lcout(),
            .ltout(\b2v_inst.un1_reg_anterior_iv_0_0_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_1_10_LC_16_11_2 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_1_10_LC_16_11_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_1_10_LC_16_11_2 .LUT_INIT=16'b1111000011110001;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_1_10_LC_16_11_2  (
            .in0(N__31116),
            .in1(N__26540),
            .in2(N__26534),
            .in3(N__30607),
            .lcout(\b2v_inst.un1_reg_anterior_iv_0_1_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_3_6_LC_16_11_3 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_3_6_LC_16_11_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_3_6_LC_16_11_3 .LUT_INIT=16'b0101111100001111;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_3_6_LC_16_11_3  (
            .in0(N__26678),
            .in1(_gnd_net_),
            .in2(N__30981),
            .in3(N__31115),
            .lcout(),
            .ltout(\b2v_inst.un1_reg_anterior_iv_0_0_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_1_6_LC_16_11_4 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_1_6_LC_16_11_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_1_6_LC_16_11_4 .LUT_INIT=16'b1111000011110001;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_1_6_LC_16_11_4  (
            .in0(N__31117),
            .in1(N__26657),
            .in2(N__26660),
            .in3(N__30606),
            .lcout(\b2v_inst.un1_reg_anterior_iv_0_1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_2_6_LC_16_11_5 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_2_6_LC_16_11_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_2_6_LC_16_11_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_2_6_LC_16_11_5  (
            .in0(N__32536),
            .in1(N__27350),
            .in2(_gnd_net_),
            .in3(N__29486),
            .lcout(\b2v_inst.N_272 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNILIBG_20_LC_16_11_6 .C_ON=1'b0;
    defparam \b2v_inst.state_RNILIBG_20_LC_16_11_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNILIBG_20_LC_16_11_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \b2v_inst.state_RNILIBG_20_LC_16_11_6  (
            .in0(N__31118),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30946),
            .lcout(\b2v_inst.data_a_escribir_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_3_LC_16_11_7 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_3_LC_16_11_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.data_a_escribir_3_LC_16_11_7 .LUT_INIT=16'b0001001111001110;
    LogicCell40 \b2v_inst.data_a_escribir_3_LC_16_11_7  (
            .in0(N__30608),
            .in1(N__31119),
            .in2(N__29120),
            .in3(N__29852),
            .lcout(b2v_inst_data_a_escribir_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34391),
            .ce(N__30556),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir11_1_c_RNO_LC_16_12_0 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir11_1_c_RNO_LC_16_12_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir11_1_c_RNO_LC_16_12_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst.data_a_escribir11_1_c_RNO_LC_16_12_0  (
            .in0(N__29552),
            .in1(N__29474),
            .in2(N__29395),
            .in3(N__29633),
            .lcout(\b2v_inst.data_a_escribir11_1_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_3_4_LC_16_12_1 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_3_4_LC_16_12_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_3_4_LC_16_12_1 .LUT_INIT=16'b0101010111011101;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_3_4_LC_16_12_1  (
            .in0(N__30945),
            .in1(N__31164),
            .in2(_gnd_net_),
            .in3(N__26618),
            .lcout(),
            .ltout(\b2v_inst.un1_reg_anterior_iv_0_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_1_4_LC_16_12_2 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_1_4_LC_16_12_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_1_4_LC_16_12_2 .LUT_INIT=16'b1111000011110001;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_1_4_LC_16_12_2  (
            .in0(N__31165),
            .in1(N__26597),
            .in2(N__26603),
            .in3(N__30612),
            .lcout(),
            .ltout(\b2v_inst.un1_reg_anterior_iv_0_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_4_LC_16_12_3 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_4_LC_16_12_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.data_a_escribir_4_LC_16_12_3 .LUT_INIT=16'b0000111100001101;
    LogicCell40 \b2v_inst.data_a_escribir_4_LC_16_12_3  (
            .in0(N__30614),
            .in1(N__31167),
            .in2(N__26600),
            .in3(N__26819),
            .lcout(b2v_inst_data_a_escribir_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34396),
            .ce(N__30552),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_2_4_LC_16_12_4 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_2_4_LC_16_12_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_2_4_LC_16_12_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_2_4_LC_16_12_4  (
            .in0(N__33020),
            .in1(N__29634),
            .in2(_gnd_net_),
            .in3(N__32539),
            .lcout(\b2v_inst.N_274 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_2_7_LC_16_12_5 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_2_7_LC_16_12_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_2_7_LC_16_12_5 .LUT_INIT=16'b0101111100111111;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_2_7_LC_16_12_5  (
            .in0(N__27586),
            .in1(N__29390),
            .in2(N__30980),
            .in3(N__32538),
            .lcout(\b2v_inst.data_a_escribir_RNO_2Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_0_4_LC_16_12_6 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_0_4_LC_16_12_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_0_4_LC_16_12_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_0_4_LC_16_12_6  (
            .in0(N__30176),
            .in1(N__31442),
            .in2(_gnd_net_),
            .in3(N__32408),
            .lcout(\b2v_inst.N_268 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_10_LC_16_12_7 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_10_LC_16_12_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.data_a_escribir_10_LC_16_12_7 .LUT_INIT=16'b0000000011111101;
    LogicCell40 \b2v_inst.data_a_escribir_10_LC_16_12_7  (
            .in0(N__30613),
            .in1(N__31166),
            .in2(N__32324),
            .in3(N__26813),
            .lcout(b2v_inst_data_a_escribir_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34396),
            .ce(N__30552),
            .sr(_gnd_net_));
    defparam \b2v_inst4.reg_data_3_LC_16_13_0 .C_ON=1'b0;
    defparam \b2v_inst4.reg_data_3_LC_16_13_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst4.reg_data_3_LC_16_13_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst4.reg_data_3_LC_16_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26807),
            .lcout(SYNTHESIZED_WIRE_5_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34408),
            .ce(N__28783),
            .sr(N__38113));
    defparam \b2v_inst4.reg_data_4_LC_16_13_1 .C_ON=1'b0;
    defparam \b2v_inst4.reg_data_4_LC_16_13_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst4.reg_data_4_LC_16_13_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst4.reg_data_4_LC_16_13_1  (
            .in0(N__26780),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(SYNTHESIZED_WIRE_5_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34408),
            .ce(N__28783),
            .sr(N__38113));
    defparam \b2v_inst4.reg_data_6_LC_16_13_2 .C_ON=1'b0;
    defparam \b2v_inst4.reg_data_6_LC_16_13_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst4.reg_data_6_LC_16_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst4.reg_data_6_LC_16_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26762),
            .lcout(SYNTHESIZED_WIRE_5_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34408),
            .ce(N__28783),
            .sr(N__38113));
    defparam \b2v_inst4.reg_data_7_LC_16_13_3 .C_ON=1'b0;
    defparam \b2v_inst4.reg_data_7_LC_16_13_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst4.reg_data_7_LC_16_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst4.reg_data_7_LC_16_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26744),
            .lcout(SYNTHESIZED_WIRE_5_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34408),
            .ce(N__28783),
            .sr(N__38113));
    defparam \b2v_inst4.reg_data_0_LC_16_13_5 .C_ON=1'b0;
    defparam \b2v_inst4.reg_data_0_LC_16_13_5 .SEQ_MODE=4'b1010;
    defparam \b2v_inst4.reg_data_0_LC_16_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst4.reg_data_0_LC_16_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26720),
            .lcout(SYNTHESIZED_WIRE_5_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34408),
            .ce(N__28783),
            .sr(N__38113));
    defparam \b2v_inst.un12_pix_count_intlto7_N_2L1_LC_16_14_1 .C_ON=1'b0;
    defparam \b2v_inst.un12_pix_count_intlto7_N_2L1_LC_16_14_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un12_pix_count_intlto7_N_2L1_LC_16_14_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst.un12_pix_count_intlto7_N_2L1_LC_16_14_1  (
            .in0(N__26965),
            .in1(N__26998),
            .in2(N__30277),
            .in3(N__26689),
            .lcout(),
            .ltout(\b2v_inst.un12_pix_count_intlto7_N_2LZ0Z1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un12_pix_count_intlto7_LC_16_14_2 .C_ON=1'b0;
    defparam \b2v_inst.un12_pix_count_intlto7_LC_16_14_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un12_pix_count_intlto7_LC_16_14_2 .LUT_INIT=16'b1111011100000000;
    LogicCell40 \b2v_inst.un12_pix_count_intlto7_LC_16_14_2  (
            .in0(N__27073),
            .in1(N__28840),
            .in2(N__27062),
            .in3(N__28823),
            .lcout(\b2v_inst.un13_pix_count_int_li_0 ),
            .ltout(\b2v_inst.un13_pix_count_int_li_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNI3K574_29_LC_16_14_3 .C_ON=1'b0;
    defparam \b2v_inst.state_RNI3K574_29_LC_16_14_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNI3K574_29_LC_16_14_3 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \b2v_inst.state_RNI3K574_29_LC_16_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27032),
            .in3(N__28208),
            .lcout(\b2v_inst.N_654_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst4.reg_data_1_LC_16_14_5 .C_ON=1'b0;
    defparam \b2v_inst4.reg_data_1_LC_16_14_5 .SEQ_MODE=4'b1010;
    defparam \b2v_inst4.reg_data_1_LC_16_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst4.reg_data_1_LC_16_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27029),
            .lcout(SYNTHESIZED_WIRE_5_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34415),
            .ce(N__28779),
            .sr(N__38116));
    defparam \b2v_inst4.reg_data_2_LC_16_14_7 .C_ON=1'b0;
    defparam \b2v_inst4.reg_data_2_LC_16_14_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst4.reg_data_2_LC_16_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst4.reg_data_2_LC_16_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26987),
            .lcout(SYNTHESIZED_WIRE_5_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34415),
            .ce(N__28779),
            .sr(N__38116));
    defparam \b2v_inst.state_fast_RNITDD01_19_LC_16_15_1 .C_ON=1'b0;
    defparam \b2v_inst.state_fast_RNITDD01_19_LC_16_15_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_fast_RNITDD01_19_LC_16_15_1 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \b2v_inst.state_fast_RNITDD01_19_LC_16_15_1  (
            .in0(N__34745),
            .in1(N__37498),
            .in2(N__26954),
            .in3(N__33187),
            .lcout(\b2v_inst.N_484 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst9.fsm_state_RNO_0_0_LC_16_15_5 .C_ON=1'b0;
    defparam \b2v_inst9.fsm_state_RNO_0_0_LC_16_15_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst9.fsm_state_RNO_0_0_LC_16_15_5 .LUT_INIT=16'b0001000111000000;
    LogicCell40 \b2v_inst9.fsm_state_RNO_0_0_LC_16_15_5  (
            .in0(N__30471),
            .in1(N__27191),
            .in2(N__26915),
            .in3(N__26897),
            .lcout(\b2v_inst9.fsm_state_srsts_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst9.bit_counter_RNIM4971_3_LC_16_16_1 .C_ON=1'b0;
    defparam \b2v_inst9.bit_counter_RNIM4971_3_LC_16_16_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst9.bit_counter_RNIM4971_3_LC_16_16_1 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \b2v_inst9.bit_counter_RNIM4971_3_LC_16_16_1  (
            .in0(N__28693),
            .in1(N__28632),
            .in2(N__28676),
            .in3(N__28707),
            .lcout(\b2v_inst9.N_522 ),
            .ltout(\b2v_inst9.N_522_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst9.fsm_state_RNIND1P1_0_LC_16_16_2 .C_ON=1'b0;
    defparam \b2v_inst9.fsm_state_RNIND1P1_0_LC_16_16_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst9.fsm_state_RNIND1P1_0_LC_16_16_2 .LUT_INIT=16'b0111011101111111;
    LogicCell40 \b2v_inst9.fsm_state_RNIND1P1_0_LC_16_16_2  (
            .in0(N__27844),
            .in1(N__27189),
            .in2(N__26906),
            .in3(N__26874),
            .lcout(\b2v_inst9.fsm_state_RNIND1P1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst9.bit_counter_RNIBIKJ_1_LC_16_16_4 .C_ON=1'b0;
    defparam \b2v_inst9.bit_counter_RNIBIKJ_1_LC_16_16_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst9.bit_counter_RNIBIKJ_1_LC_16_16_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \b2v_inst9.bit_counter_RNIBIKJ_1_LC_16_16_4  (
            .in0(_gnd_net_),
            .in1(N__28671),
            .in2(_gnd_net_),
            .in3(N__28692),
            .lcout(),
            .ltout(\b2v_inst9.N_84_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst9.bit_counter_RNIJOID1_3_LC_16_16_5 .C_ON=1'b0;
    defparam \b2v_inst9.bit_counter_RNIJOID1_3_LC_16_16_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst9.bit_counter_RNIJOID1_3_LC_16_16_5 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \b2v_inst9.bit_counter_RNIJOID1_3_LC_16_16_5  (
            .in0(N__27190),
            .in1(N__28633),
            .in2(N__27104),
            .in3(N__28708),
            .lcout(\b2v_inst9.N_582 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_2_cry_0_c_LC_17_5_0 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_2_cry_0_c_LC_17_5_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_2_cry_0_c_LC_17_5_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final4_2_cry_0_c_LC_17_5_0  (
            .in0(_gnd_net_),
            .in1(N__29023),
            .in2(N__27434),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_17_5_0_),
            .carryout(\b2v_inst.valor_max_final4_2_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_2_cry_1_c_LC_17_5_1 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_2_cry_1_c_LC_17_5_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_2_cry_1_c_LC_17_5_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final4_2_cry_1_c_LC_17_5_1  (
            .in0(_gnd_net_),
            .in1(N__31351),
            .in2(N__28951),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.valor_max_final4_2_cry_0 ),
            .carryout(\b2v_inst.valor_max_final4_2_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_2_cry_2_c_LC_17_5_2 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_2_cry_2_c_LC_17_5_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_2_cry_2_c_LC_17_5_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final4_2_cry_2_c_LC_17_5_2  (
            .in0(_gnd_net_),
            .in1(N__31300),
            .in2(N__28916),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.valor_max_final4_2_cry_1 ),
            .carryout(\b2v_inst.valor_max_final4_2_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_2_cry_3_c_LC_17_5_3 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_2_cry_3_c_LC_17_5_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_2_cry_3_c_LC_17_5_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final4_2_cry_3_c_LC_17_5_3  (
            .in0(_gnd_net_),
            .in1(N__28882),
            .in2(N__32459),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.valor_max_final4_2_cry_2 ),
            .carryout(\b2v_inst.valor_max_final4_2_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_2_cry_4_c_LC_17_5_4 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_2_cry_4_c_LC_17_5_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_2_cry_4_c_LC_17_5_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final4_2_cry_4_c_LC_17_5_4  (
            .in0(_gnd_net_),
            .in1(N__33019),
            .in2(N__29591),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.valor_max_final4_2_cry_3 ),
            .carryout(\b2v_inst.valor_max_final4_2_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_2_cry_5_c_LC_17_5_5 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_2_cry_5_c_LC_17_5_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_2_cry_5_c_LC_17_5_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final4_2_cry_5_c_LC_17_5_5  (
            .in0(_gnd_net_),
            .in1(N__29512),
            .in2(N__27394),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.valor_max_final4_2_cry_4 ),
            .carryout(\b2v_inst.valor_max_final4_2_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_2_cry_6_c_LC_17_5_6 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_2_cry_6_c_LC_17_5_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_2_cry_6_c_LC_17_5_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final4_2_cry_6_c_LC_17_5_6  (
            .in0(_gnd_net_),
            .in1(N__29426),
            .in2(N__27348),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.valor_max_final4_2_cry_5 ),
            .carryout(\b2v_inst.valor_max_final4_2_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_2_cry_7_c_LC_17_5_7 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_2_cry_7_c_LC_17_5_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_2_cry_7_c_LC_17_5_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final4_2_cry_7_c_LC_17_5_7  (
            .in0(_gnd_net_),
            .in1(N__29351),
            .in2(N__27590),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.valor_max_final4_2_cry_6 ),
            .carryout(\b2v_inst.valor_max_final4_2_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_2_cry_8_c_LC_17_6_0 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_2_cry_8_c_LC_17_6_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_2_cry_8_c_LC_17_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final4_2_cry_8_c_LC_17_6_0  (
            .in0(_gnd_net_),
            .in1(N__29320),
            .in2(N__29926),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_17_6_0_),
            .carryout(\b2v_inst.valor_max_final4_2_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_2_cry_9_c_LC_17_6_1 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_2_cry_9_c_LC_17_6_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_2_cry_9_c_LC_17_6_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final4_2_cry_9_c_LC_17_6_1  (
            .in0(_gnd_net_),
            .in1(N__29726),
            .in2(N__29291),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.valor_max_final4_2_cry_8 ),
            .carryout(\b2v_inst.valor_max_final4_2_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_2_cry_10_c_LC_17_6_2 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_2_cry_10_c_LC_17_6_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_2_cry_10_c_LC_17_6_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final4_2_cry_10_c_LC_17_6_2  (
            .in0(_gnd_net_),
            .in1(N__31489),
            .in2(N__29213),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.valor_max_final4_2_cry_9 ),
            .carryout(\b2v_inst.valor_max_final42 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_2_cry_10_c_RNI9G0Q_LC_17_6_3 .C_ON=1'b0;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_2_cry_10_c_RNI9G0Q_LC_17_6_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_2_cry_10_c_RNI9G0Q_LC_17_6_3 .LUT_INIT=16'b0000101101011011;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final4_2_cry_10_c_RNI9G0Q_LC_17_6_3  (
            .in0(N__32349),
            .in1(N__29177),
            .in2(N__32542),
            .in3(N__27299),
            .lcout(\b2v_inst.m54_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir11_7_c_RNO_LC_17_7_0 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir11_7_c_RNO_LC_17_7_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir11_7_c_RNO_LC_17_7_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst.data_a_escribir11_7_c_RNO_LC_17_7_0  (
            .in0(N__30723),
            .in1(N__30691),
            .in2(N__30136),
            .in3(N__29443),
            .lcout(\b2v_inst.data_a_escribir11_7_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.reg_ancho_3_6_LC_17_7_2 .C_ON=1'b0;
    defparam \b2v_inst.reg_ancho_3_6_LC_17_7_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_ancho_3_6_LC_17_7_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \b2v_inst.reg_ancho_3_6_LC_17_7_2  (
            .in0(N__31905),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31563),
            .lcout(\b2v_inst.reg_ancho_3Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34416),
            .ce(N__32060),
            .sr(N__38117));
    defparam \b2v_inst.reg_ancho_3_7_LC_17_7_3 .C_ON=1'b0;
    defparam \b2v_inst.reg_ancho_3_7_LC_17_7_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_ancho_3_7_LC_17_7_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \b2v_inst.reg_ancho_3_7_LC_17_7_3  (
            .in0(_gnd_net_),
            .in1(N__27270),
            .in2(_gnd_net_),
            .in3(N__31906),
            .lcout(\b2v_inst.reg_ancho_3Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34416),
            .ce(N__32060),
            .sr(N__38117));
    defparam \b2v_inst.reg_ancho_3_8_LC_17_7_4 .C_ON=1'b0;
    defparam \b2v_inst.reg_ancho_3_8_LC_17_7_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_ancho_3_8_LC_17_7_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \b2v_inst.reg_ancho_3_8_LC_17_7_4  (
            .in0(N__31907),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27250),
            .lcout(\b2v_inst.reg_ancho_3Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34416),
            .ce(N__32060),
            .sr(N__38117));
    defparam \b2v_inst.reg_ancho_3_9_LC_17_7_5 .C_ON=1'b0;
    defparam \b2v_inst.reg_ancho_3_9_LC_17_7_5 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_ancho_3_9_LC_17_7_5 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \b2v_inst.reg_ancho_3_9_LC_17_7_5  (
            .in0(N__31989),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31908),
            .lcout(\b2v_inst.reg_ancho_3Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34416),
            .ce(N__32060),
            .sr(N__38117));
    defparam \b2v_inst.reg_ancho_3_1_LC_17_7_6 .C_ON=1'b0;
    defparam \b2v_inst.reg_ancho_3_1_LC_17_7_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_ancho_3_1_LC_17_7_6 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \b2v_inst.reg_ancho_3_1_LC_17_7_6  (
            .in0(N__31904),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31396),
            .lcout(\b2v_inst.reg_ancho_3Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34416),
            .ce(N__32060),
            .sr(N__38117));
    defparam \b2v_inst.reg_ancho_3_0_LC_17_7_7 .C_ON=1'b0;
    defparam \b2v_inst.reg_ancho_3_0_LC_17_7_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_ancho_3_0_LC_17_7_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \b2v_inst.reg_ancho_3_0_LC_17_7_7  (
            .in0(_gnd_net_),
            .in1(N__31903),
            .in2(_gnd_net_),
            .in3(N__27487),
            .lcout(\b2v_inst.reg_ancho_3Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34416),
            .ce(N__32060),
            .sr(N__38117));
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_3_cry_0_c_LC_17_8_0 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_3_cry_0_c_LC_17_8_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_3_cry_0_c_LC_17_8_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final4_3_cry_0_c_LC_17_8_0  (
            .in0(_gnd_net_),
            .in1(N__27505),
            .in2(N__27448),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_17_8_0_),
            .carryout(\b2v_inst.valor_max_final4_3_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_3_cry_1_c_LC_17_8_1 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_3_cry_1_c_LC_17_8_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_3_cry_1_c_LC_17_8_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final4_3_cry_1_c_LC_17_8_1  (
            .in0(_gnd_net_),
            .in1(N__27745),
            .in2(N__31352),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.valor_max_final4_3_cry_0 ),
            .carryout(\b2v_inst.valor_max_final4_3_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_3_cry_2_c_LC_17_8_2 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_3_cry_2_c_LC_17_8_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_3_cry_2_c_LC_17_8_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final4_3_cry_2_c_LC_17_8_2  (
            .in0(_gnd_net_),
            .in1(N__27727),
            .in2(N__31304),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.valor_max_final4_3_cry_1 ),
            .carryout(\b2v_inst.valor_max_final4_3_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_3_cry_3_c_LC_17_8_3 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_3_cry_3_c_LC_17_8_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_3_cry_3_c_LC_17_8_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final4_3_cry_3_c_LC_17_8_3  (
            .in0(_gnd_net_),
            .in1(N__27709),
            .in2(N__32458),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.valor_max_final4_3_cry_2 ),
            .carryout(\b2v_inst.valor_max_final4_3_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_3_cry_4_c_LC_17_8_4 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_3_cry_4_c_LC_17_8_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_3_cry_4_c_LC_17_8_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final4_3_cry_4_c_LC_17_8_4  (
            .in0(_gnd_net_),
            .in1(N__33014),
            .in2(N__27692),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.valor_max_final4_3_cry_3 ),
            .carryout(\b2v_inst.valor_max_final4_3_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_3_cry_5_c_LC_17_8_5 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_3_cry_5_c_LC_17_8_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_3_cry_5_c_LC_17_8_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final4_3_cry_5_c_LC_17_8_5  (
            .in0(_gnd_net_),
            .in1(N__27393),
            .in2(N__27671),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.valor_max_final4_3_cry_4 ),
            .carryout(\b2v_inst.valor_max_final4_3_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_3_cry_6_c_LC_17_8_6 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_3_cry_6_c_LC_17_8_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_3_cry_6_c_LC_17_8_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final4_3_cry_6_c_LC_17_8_6  (
            .in0(_gnd_net_),
            .in1(N__27649),
            .in2(N__27349),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.valor_max_final4_3_cry_5 ),
            .carryout(\b2v_inst.valor_max_final4_3_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_3_cry_7_c_LC_17_8_7 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_3_cry_7_c_LC_17_8_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_3_cry_7_c_LC_17_8_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final4_3_cry_7_c_LC_17_8_7  (
            .in0(_gnd_net_),
            .in1(N__27585),
            .in2(N__27632),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.valor_max_final4_3_cry_6 ),
            .carryout(\b2v_inst.valor_max_final4_3_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_3_cry_8_c_LC_17_9_0 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_3_cry_8_c_LC_17_9_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_3_cry_8_c_LC_17_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final4_3_cry_8_c_LC_17_9_0  (
            .in0(_gnd_net_),
            .in1(N__29927),
            .in2(N__27611),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_17_9_0_),
            .carryout(\b2v_inst.valor_max_final4_3_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_3_cry_9_c_LC_17_9_1 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_3_cry_9_c_LC_17_9_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_3_cry_9_c_LC_17_9_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final4_3_cry_9_c_LC_17_9_1  (
            .in0(_gnd_net_),
            .in1(N__29737),
            .in2(N__28406),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.valor_max_final4_3_cry_8 ),
            .carryout(\b2v_inst.valor_max_final4_3_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_3_cry_10_c_LC_17_9_2 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_3_cry_10_c_LC_17_9_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_3_cry_10_c_LC_17_9_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final4_3_cry_10_c_LC_17_9_2  (
            .in0(_gnd_net_),
            .in1(N__31483),
            .in2(N__28385),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.valor_max_final4_3_cry_9 ),
            .carryout(\b2v_inst.valor_max_final43 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.valor_max_final43_THRU_LUT4_0_LC_17_9_3 .C_ON=1'b0;
    defparam \b2v_inst.valor_max_final43_THRU_LUT4_0_LC_17_9_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.valor_max_final43_THRU_LUT4_0_LC_17_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.valor_max_final43_THRU_LUT4_0_LC_17_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27542),
            .lcout(\b2v_inst.valor_max_final43_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_0_0_LC_17_9_4 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_0_0_LC_17_9_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_0_0_LC_17_9_4 .LUT_INIT=16'b0100111101111111;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_0_0_LC_17_9_4  (
            .in0(N__28615),
            .in1(N__32405),
            .in2(N__30987),
            .in3(N__29674),
            .lcout(\b2v_inst.data_a_escribir_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_0_1_LC_17_9_6 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_0_1_LC_17_9_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_0_1_LC_17_9_6 .LUT_INIT=16'b0101111100111111;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_0_1_LC_17_9_6  (
            .in0(N__28589),
            .in1(N__29701),
            .in2(N__30988),
            .in3(N__32406),
            .lcout(\b2v_inst.data_a_escribir_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_3_5_LC_17_9_7 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_3_5_LC_17_9_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_3_5_LC_17_9_7 .LUT_INIT=16'b0111011100110011;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_3_5_LC_17_9_7  (
            .in0(N__27527),
            .in1(N__30961),
            .in2(_gnd_net_),
            .in3(N__31129),
            .lcout(\b2v_inst.un1_reg_anterior_iv_0_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_1_cry_0_c_inv_LC_17_10_0 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_1_cry_0_c_inv_LC_17_10_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_1_cry_0_c_inv_LC_17_10_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final4_1_cry_0_c_inv_LC_17_10_0  (
            .in0(_gnd_net_),
            .in1(N__29066),
            .in2(N__27506),
            .in3(N__28610),
            .lcout(\b2v_inst.reg_anterior_i_0 ),
            .ltout(),
            .carryin(bfn_17_10_0_),
            .carryout(\b2v_inst.valor_max_final4_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_1_cry_1_c_inv_LC_17_10_1 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_1_cry_1_c_inv_LC_17_10_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_1_cry_1_c_inv_LC_17_10_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final4_1_cry_1_c_inv_LC_17_10_1  (
            .in0(N__28574),
            .in1(N__28994),
            .in2(N__27746),
            .in3(_gnd_net_),
            .lcout(\b2v_inst.reg_anterior_i_1 ),
            .ltout(),
            .carryin(\b2v_inst.valor_max_final4_1_cry_0 ),
            .carryout(\b2v_inst.valor_max_final4_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_1_cry_2_c_inv_LC_17_10_2 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_1_cry_2_c_inv_LC_17_10_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_1_cry_2_c_inv_LC_17_10_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final4_1_cry_2_c_inv_LC_17_10_2  (
            .in0(_gnd_net_),
            .in1(N__31256),
            .in2(N__27728),
            .in3(N__29837),
            .lcout(\b2v_inst.reg_anterior_i_2 ),
            .ltout(),
            .carryin(\b2v_inst.valor_max_final4_1_cry_1 ),
            .carryout(\b2v_inst.valor_max_final4_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_1_cry_3_c_inv_LC_17_10_3 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_1_cry_3_c_inv_LC_17_10_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_1_cry_3_c_inv_LC_17_10_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final4_1_cry_3_c_inv_LC_17_10_3  (
            .in0(N__29158),
            .in1(N__31041),
            .in2(N__27710),
            .in3(_gnd_net_),
            .lcout(\b2v_inst.reg_anterior_i_3 ),
            .ltout(),
            .carryin(\b2v_inst.valor_max_final4_1_cry_2 ),
            .carryout(\b2v_inst.valor_max_final4_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_1_cry_4_c_inv_LC_17_10_4 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_1_cry_4_c_inv_LC_17_10_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_1_cry_4_c_inv_LC_17_10_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final4_1_cry_4_c_inv_LC_17_10_4  (
            .in0(_gnd_net_),
            .in1(N__29636),
            .in2(N__27691),
            .in3(N__30171),
            .lcout(\b2v_inst.reg_anterior_i_4 ),
            .ltout(),
            .carryin(\b2v_inst.valor_max_final4_1_cry_3 ),
            .carryout(\b2v_inst.valor_max_final4_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_1_cry_5_c_inv_LC_17_10_5 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_1_cry_5_c_inv_LC_17_10_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_1_cry_5_c_inv_LC_17_10_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final4_1_cry_5_c_inv_LC_17_10_5  (
            .in0(_gnd_net_),
            .in1(N__29559),
            .in2(N__27670),
            .in3(N__29101),
            .lcout(\b2v_inst.reg_anterior_i_5 ),
            .ltout(),
            .carryin(\b2v_inst.valor_max_final4_1_cry_4 ),
            .carryout(\b2v_inst.valor_max_final4_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_1_cry_6_c_inv_LC_17_10_6 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_1_cry_6_c_inv_LC_17_10_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_1_cry_6_c_inv_LC_17_10_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final4_1_cry_6_c_inv_LC_17_10_6  (
            .in0(N__31525),
            .in1(N__29485),
            .in2(N__27650),
            .in3(_gnd_net_),
            .lcout(\b2v_inst.reg_anterior_i_6 ),
            .ltout(),
            .carryin(\b2v_inst.valor_max_final4_1_cry_5 ),
            .carryout(\b2v_inst.valor_max_final4_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_1_cry_7_c_inv_LC_17_10_7 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_1_cry_7_c_inv_LC_17_10_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_1_cry_7_c_inv_LC_17_10_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final4_1_cry_7_c_inv_LC_17_10_7  (
            .in0(_gnd_net_),
            .in1(N__29396),
            .in2(N__27631),
            .in3(N__30657),
            .lcout(\b2v_inst.reg_anterior_i_7 ),
            .ltout(),
            .carryin(\b2v_inst.valor_max_final4_1_cry_6 ),
            .carryout(\b2v_inst.valor_max_final4_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_1_cry_8_c_inv_LC_17_11_0 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_1_cry_8_c_inv_LC_17_11_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_1_cry_8_c_inv_LC_17_11_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final4_1_cry_8_c_inv_LC_17_11_0  (
            .in0(_gnd_net_),
            .in1(N__29966),
            .in2(N__27610),
            .in3(N__30761),
            .lcout(\b2v_inst.reg_anterior_i_8 ),
            .ltout(),
            .carryin(bfn_17_11_0_),
            .carryout(\b2v_inst.valor_max_final4_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_1_cry_9_c_inv_LC_17_11_1 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_1_cry_9_c_inv_LC_17_11_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_1_cry_9_c_inv_LC_17_11_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final4_1_cry_9_c_inv_LC_17_11_1  (
            .in0(N__31950),
            .in1(N__30003),
            .in2(N__28405),
            .in3(_gnd_net_),
            .lcout(\b2v_inst.reg_anterior_i_9 ),
            .ltout(),
            .carryin(\b2v_inst.valor_max_final4_1_cry_8 ),
            .carryout(\b2v_inst.valor_max_final4_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_1_cry_10_c_inv_LC_17_11_2 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_1_cry_10_c_inv_LC_17_11_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_1_cry_10_c_inv_LC_17_11_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final4_1_cry_10_c_inv_LC_17_11_2  (
            .in0(_gnd_net_),
            .in1(N__29257),
            .in2(N__28384),
            .in3(N__31719),
            .lcout(\b2v_inst.reg_anterior_i_10 ),
            .ltout(),
            .carryin(\b2v_inst.valor_max_final4_1_cry_9 ),
            .carryout(\b2v_inst.valor_max_final41 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_3_cry_10_c_RNIUCPE1_LC_17_11_3 .C_ON=1'b0;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_3_cry_10_c_RNIUCPE1_LC_17_11_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_3_cry_10_c_RNIUCPE1_LC_17_11_3 .LUT_INIT=16'b0011010011110100;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final4_3_cry_10_c_RNIUCPE1_LC_17_11_3  (
            .in0(N__28364),
            .in1(N__32398),
            .in2(N__28355),
            .in3(N__28343),
            .lcout(\b2v_inst.N_711 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.reg_anterior_1_LC_17_11_7 .C_ON=1'b0;
    defparam \b2v_inst.reg_anterior_1_LC_17_11_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_anterior_1_LC_17_11_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \b2v_inst.reg_anterior_1_LC_17_11_7  (
            .in0(_gnd_net_),
            .in1(N__31858),
            .in2(_gnd_net_),
            .in3(N__31400),
            .lcout(\b2v_inst.reg_anteriorZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34380),
            .ce(N__31672),
            .sr(N__38107));
    defparam \b2v_inst.state_RNO_4_31_LC_17_12_1 .C_ON=1'b0;
    defparam \b2v_inst.state_RNO_4_31_LC_17_12_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNO_4_31_LC_17_12_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst.state_RNO_4_31_LC_17_12_1  (
            .in0(N__28340),
            .in1(N__28206),
            .in2(N__27920),
            .in3(N__28253),
            .lcout(\b2v_inst.N_694 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNO_5_31_LC_17_12_2 .C_ON=1'b0;
    defparam \b2v_inst.state_RNO_5_31_LC_17_12_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNO_5_31_LC_17_12_2 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \b2v_inst.state_RNO_5_31_LC_17_12_2  (
            .in0(N__28207),
            .in1(N__28076),
            .in2(N__28067),
            .in3(N__27918),
            .lcout(),
            .ltout(\b2v_inst.N_695_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNO_0_31_LC_17_12_3 .C_ON=1'b0;
    defparam \b2v_inst.state_RNO_0_31_LC_17_12_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNO_0_31_LC_17_12_3 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \b2v_inst.state_RNO_0_31_LC_17_12_3  (
            .in0(N__27962),
            .in1(N__28025),
            .in2(N__28019),
            .in3(N__28004),
            .lcout(\b2v_inst.state_ns_a3_i_0_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_32_rep1_RNIUROT1_LC_17_12_4 .C_ON=1'b0;
    defparam \b2v_inst.state_32_rep1_RNIUROT1_LC_17_12_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_32_rep1_RNIUROT1_LC_17_12_4 .LUT_INIT=16'b1111011111110000;
    LogicCell40 \b2v_inst.state_32_rep1_RNIUROT1_LC_17_12_4  (
            .in0(N__28003),
            .in1(N__27961),
            .in2(N__30983),
            .in3(N__27917),
            .lcout(),
            .ltout(\b2v_inst.un1_reset_inv_0_0_tz_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_32_rep1_RNIP5K4F_LC_17_12_5 .C_ON=1'b0;
    defparam \b2v_inst.state_32_rep1_RNIP5K4F_LC_17_12_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_32_rep1_RNIP5K4F_LC_17_12_5 .LUT_INIT=16'b1010000010101000;
    LogicCell40 \b2v_inst.state_32_rep1_RNIP5K4F_LC_17_12_5  (
            .in0(N__27833),
            .in1(N__28546),
            .in2(N__28529),
            .in3(N__28525),
            .lcout(\b2v_inst.un1_reset_inv_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_1_7_LC_17_12_6 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_1_7_LC_17_12_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_1_7_LC_17_12_6 .LUT_INIT=16'b0010101001111111;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_1_7_LC_17_12_6  (
            .in0(N__31176),
            .in1(N__30956),
            .in2(N__28490),
            .in3(N__28469),
            .lcout(\b2v_inst.un1_reg_anterior_0_i_1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst9.un1_cycle_counter_2_cry_0_c_LC_17_13_0 .C_ON=1'b1;
    defparam \b2v_inst9.un1_cycle_counter_2_cry_0_c_LC_17_13_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst9.un1_cycle_counter_2_cry_0_c_LC_17_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst9.un1_cycle_counter_2_cry_0_c_LC_17_13_0  (
            .in0(_gnd_net_),
            .in1(N__30416),
            .in2(N__30308),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_17_13_0_),
            .carryout(\b2v_inst9.un1_cycle_counter_2_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst9.un1_cycle_counter_2_cry_0_THRU_LUT4_0_LC_17_13_1 .C_ON=1'b1;
    defparam \b2v_inst9.un1_cycle_counter_2_cry_0_THRU_LUT4_0_LC_17_13_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst9.un1_cycle_counter_2_cry_0_THRU_LUT4_0_LC_17_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst9.un1_cycle_counter_2_cry_0_THRU_LUT4_0_LC_17_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__28427),
            .in3(N__28463),
            .lcout(\b2v_inst9.un1_cycle_counter_2_cry_0_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst9.un1_cycle_counter_2_cry_0 ),
            .carryout(\b2v_inst9.un1_cycle_counter_2_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst9.un1_cycle_counter_2_cry_1_THRU_LUT4_0_LC_17_13_2 .C_ON=1'b1;
    defparam \b2v_inst9.un1_cycle_counter_2_cry_1_THRU_LUT4_0_LC_17_13_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst9.un1_cycle_counter_2_cry_1_THRU_LUT4_0_LC_17_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst9.un1_cycle_counter_2_cry_1_THRU_LUT4_0_LC_17_13_2  (
            .in0(_gnd_net_),
            .in1(N__30493),
            .in2(_gnd_net_),
            .in3(N__28460),
            .lcout(\b2v_inst9.un1_cycle_counter_2_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst9.un1_cycle_counter_2_cry_1 ),
            .carryout(\b2v_inst9.un1_cycle_counter_2_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst9.cycle_counter_3_LC_17_13_3 .C_ON=1'b0;
    defparam \b2v_inst9.cycle_counter_3_LC_17_13_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst9.cycle_counter_3_LC_17_13_3 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \b2v_inst9.cycle_counter_3_LC_17_13_3  (
            .in0(N__28453),
            .in1(N__38151),
            .in2(_gnd_net_),
            .in3(N__28457),
            .lcout(\b2v_inst9.cycle_counterZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34397),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst9.cycle_counter_RNIQAGD_0_3_LC_17_13_5 .C_ON=1'b0;
    defparam \b2v_inst9.cycle_counter_RNIQAGD_0_3_LC_17_13_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst9.cycle_counter_RNIQAGD_0_3_LC_17_13_5 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \b2v_inst9.cycle_counter_RNIQAGD_0_3_LC_17_13_5  (
            .in0(N__30304),
            .in1(N__28452),
            .in2(N__28426),
            .in3(N__30492),
            .lcout(\b2v_inst9.N_175_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst9.cycle_counter_RNIQAGD_3_LC_17_13_6 .C_ON=1'b0;
    defparam \b2v_inst9.cycle_counter_RNIQAGD_3_LC_17_13_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst9.cycle_counter_RNIQAGD_3_LC_17_13_6 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \b2v_inst9.cycle_counter_RNIQAGD_3_LC_17_13_6  (
            .in0(N__30491),
            .in1(N__28418),
            .in2(N__28454),
            .in3(N__30303),
            .lcout(\b2v_inst9.cycle_counter_RNIQAGDZ0Z_3 ),
            .ltout(\b2v_inst9.cycle_counter_RNIQAGDZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst9.cycle_counter_1_LC_17_13_7 .C_ON=1'b0;
    defparam \b2v_inst9.cycle_counter_1_LC_17_13_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst9.cycle_counter_1_LC_17_13_7 .LUT_INIT=16'b0001000000100000;
    LogicCell40 \b2v_inst9.cycle_counter_1_LC_17_13_7  (
            .in0(N__28425),
            .in1(N__38150),
            .in2(N__28436),
            .in3(N__28433),
            .lcout(\b2v_inst9.cycle_counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34397),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un12_pix_count_intlto7_N_3L3_LC_17_14_7 .C_ON=1'b0;
    defparam \b2v_inst.un12_pix_count_intlto7_N_3L3_LC_17_14_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un12_pix_count_intlto7_N_3L3_LC_17_14_7 .LUT_INIT=16'b0001000101010101;
    LogicCell40 \b2v_inst.un12_pix_count_intlto7_N_3L3_LC_17_14_7  (
            .in0(N__28852),
            .in1(N__28839),
            .in2(_gnd_net_),
            .in3(N__28795),
            .lcout(\b2v_inst.un12_pix_count_intlto7_N_3LZ0Z3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst4.reg_data_5_LC_17_15_7 .C_ON=1'b0;
    defparam \b2v_inst4.reg_data_5_LC_17_15_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst4.reg_data_5_LC_17_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst4.reg_data_5_LC_17_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28817),
            .lcout(SYNTHESIZED_WIRE_5_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34417),
            .ce(N__28784),
            .sr(N__38130));
    defparam \b2v_inst9.bit_counter_0_LC_17_16_0 .C_ON=1'b1;
    defparam \b2v_inst9.bit_counter_0_LC_17_16_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst9.bit_counter_0_LC_17_16_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst9.bit_counter_0_LC_17_16_0  (
            .in0(N__28654),
            .in1(N__28709),
            .in2(N__28727),
            .in3(N__28726),
            .lcout(\b2v_inst9.bit_counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_17_16_0_),
            .carryout(\b2v_inst9.un1_bit_counter_3_cry_0 ),
            .clk(N__34426),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst9.bit_counter_1_LC_17_16_1 .C_ON=1'b1;
    defparam \b2v_inst9.bit_counter_1_LC_17_16_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst9.bit_counter_1_LC_17_16_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst9.bit_counter_1_LC_17_16_1  (
            .in0(N__28652),
            .in1(N__28694),
            .in2(_gnd_net_),
            .in3(N__28679),
            .lcout(\b2v_inst9.bit_counterZ1Z_1 ),
            .ltout(),
            .carryin(\b2v_inst9.un1_bit_counter_3_cry_0 ),
            .carryout(\b2v_inst9.un1_bit_counter_3_cry_1 ),
            .clk(N__34426),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst9.bit_counter_2_LC_17_16_2 .C_ON=1'b1;
    defparam \b2v_inst9.bit_counter_2_LC_17_16_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst9.bit_counter_2_LC_17_16_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst9.bit_counter_2_LC_17_16_2  (
            .in0(N__28655),
            .in1(N__28675),
            .in2(_gnd_net_),
            .in3(N__28658),
            .lcout(\b2v_inst9.bit_counterZ0Z_2 ),
            .ltout(),
            .carryin(\b2v_inst9.un1_bit_counter_3_cry_1 ),
            .carryout(\b2v_inst9.un1_bit_counter_3_cry_2 ),
            .clk(N__34426),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst9.bit_counter_3_LC_17_16_3 .C_ON=1'b0;
    defparam \b2v_inst9.bit_counter_3_LC_17_16_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst9.bit_counter_3_LC_17_16_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst9.bit_counter_3_LC_17_16_3  (
            .in0(N__28653),
            .in1(N__28634),
            .in2(_gnd_net_),
            .in3(N__28637),
            .lcout(\b2v_inst9.bit_counterZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34426),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.reg_anterior_5_LC_18_5_0 .C_ON=1'b0;
    defparam \b2v_inst.reg_anterior_5_LC_18_5_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_anterior_5_LC_18_5_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \b2v_inst.reg_anterior_5_LC_18_5_0  (
            .in0(_gnd_net_),
            .in1(N__31919),
            .in2(_gnd_net_),
            .in3(N__32117),
            .lcout(\b2v_inst.reg_anteriorZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34427),
            .ce(N__31687),
            .sr(N__38136));
    defparam \b2v_inst.encontrar_maximo_un2_valor_max2_cry_0_c_LC_18_6_0 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_un2_valor_max2_cry_0_c_LC_18_6_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_un2_valor_max2_cry_0_c_LC_18_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.encontrar_maximo_un2_valor_max2_cry_0_c_LC_18_6_0  (
            .in0(_gnd_net_),
            .in1(N__28619),
            .in2(N__29024),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_18_6_0_),
            .carryout(\b2v_inst.un2_valor_max2_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_un2_valor_max2_cry_1_c_LC_18_6_1 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_un2_valor_max2_cry_1_c_LC_18_6_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_un2_valor_max2_cry_1_c_LC_18_6_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.encontrar_maximo_un2_valor_max2_cry_1_c_LC_18_6_1  (
            .in0(_gnd_net_),
            .in1(N__28584),
            .in2(N__28952),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.un2_valor_max2_cry_0 ),
            .carryout(\b2v_inst.un2_valor_max2_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_un2_valor_max2_cry_2_c_LC_18_6_2 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_un2_valor_max2_cry_2_c_LC_18_6_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_un2_valor_max2_cry_2_c_LC_18_6_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.encontrar_maximo_un2_valor_max2_cry_2_c_LC_18_6_2  (
            .in0(_gnd_net_),
            .in1(N__29839),
            .in2(N__28915),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.un2_valor_max2_cry_1 ),
            .carryout(\b2v_inst.un2_valor_max2_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_un2_valor_max2_cry_3_c_LC_18_6_3 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_un2_valor_max2_cry_3_c_LC_18_6_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_un2_valor_max2_cry_3_c_LC_18_6_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.encontrar_maximo_un2_valor_max2_cry_3_c_LC_18_6_3  (
            .in0(_gnd_net_),
            .in1(N__29153),
            .in2(N__28883),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.un2_valor_max2_cry_2 ),
            .carryout(\b2v_inst.un2_valor_max2_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_un2_valor_max2_cry_4_c_LC_18_6_4 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_un2_valor_max2_cry_4_c_LC_18_6_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_un2_valor_max2_cry_4_c_LC_18_6_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.encontrar_maximo_un2_valor_max2_cry_4_c_LC_18_6_4  (
            .in0(_gnd_net_),
            .in1(N__30158),
            .in2(N__29590),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.un2_valor_max2_cry_3 ),
            .carryout(\b2v_inst.un2_valor_max2_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_un2_valor_max2_cry_5_c_LC_18_6_5 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_un2_valor_max2_cry_5_c_LC_18_6_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_un2_valor_max2_cry_5_c_LC_18_6_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.encontrar_maximo_un2_valor_max2_cry_5_c_LC_18_6_5  (
            .in0(_gnd_net_),
            .in1(N__29090),
            .in2(N__29513),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.un2_valor_max2_cry_4 ),
            .carryout(\b2v_inst.un2_valor_max2_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_un2_valor_max2_cry_6_c_LC_18_6_6 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_un2_valor_max2_cry_6_c_LC_18_6_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_un2_valor_max2_cry_6_c_LC_18_6_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.encontrar_maximo_un2_valor_max2_cry_6_c_LC_18_6_6  (
            .in0(_gnd_net_),
            .in1(N__31514),
            .in2(N__29425),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.un2_valor_max2_cry_5 ),
            .carryout(\b2v_inst.un2_valor_max2_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_un2_valor_max2_cry_7_c_LC_18_6_7 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_un2_valor_max2_cry_7_c_LC_18_6_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_un2_valor_max2_cry_7_c_LC_18_6_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.encontrar_maximo_un2_valor_max2_cry_7_c_LC_18_6_7  (
            .in0(_gnd_net_),
            .in1(N__30669),
            .in2(N__29350),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.un2_valor_max2_cry_6 ),
            .carryout(\b2v_inst.un2_valor_max2_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_un2_valor_max2_cry_8_c_LC_18_7_0 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_un2_valor_max2_cry_8_c_LC_18_7_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_un2_valor_max2_cry_8_c_LC_18_7_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.encontrar_maximo_un2_valor_max2_cry_8_c_LC_18_7_0  (
            .in0(_gnd_net_),
            .in1(N__30770),
            .in2(N__29321),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_18_7_0_),
            .carryout(\b2v_inst.un2_valor_max2_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_un2_valor_max2_cry_9_c_LC_18_7_1 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_un2_valor_max2_cry_9_c_LC_18_7_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_un2_valor_max2_cry_9_c_LC_18_7_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.encontrar_maximo_un2_valor_max2_cry_9_c_LC_18_7_1  (
            .in0(_gnd_net_),
            .in1(N__31955),
            .in2(N__29290),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.un2_valor_max2_cry_8 ),
            .carryout(\b2v_inst.un2_valor_max2_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_un2_valor_max2_cry_10_c_LC_18_7_2 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_un2_valor_max2_cry_10_c_LC_18_7_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_un2_valor_max2_cry_10_c_LC_18_7_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.encontrar_maximo_un2_valor_max2_cry_10_c_LC_18_7_2  (
            .in0(_gnd_net_),
            .in1(N__31726),
            .in2(N__29212),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.un2_valor_max2_cry_9 ),
            .carryout(\b2v_inst.un2_valor_max2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un2_valor_max2_THRU_LUT4_0_LC_18_7_3 .C_ON=1'b0;
    defparam \b2v_inst.un2_valor_max2_THRU_LUT4_0_LC_18_7_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un2_valor_max2_THRU_LUT4_0_LC_18_7_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.un2_valor_max2_THRU_LUT4_0_LC_18_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29165),
            .lcout(\b2v_inst.un2_valor_max2_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_0_3_LC_18_7_4 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_0_3_LC_18_7_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_0_3_LC_18_7_4 .LUT_INIT=16'b0011111101011111;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_0_3_LC_18_7_4  (
            .in0(N__32231),
            .in1(N__29162),
            .in2(N__30992),
            .in3(N__32392),
            .lcout(\b2v_inst.data_a_escribir_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_0_6_LC_18_7_5 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_0_6_LC_18_7_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_0_6_LC_18_7_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_0_6_LC_18_7_5  (
            .in0(N__32393),
            .in1(N__31518),
            .in2(_gnd_net_),
            .in3(N__29444),
            .lcout(\b2v_inst.valor_max2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_0_5_LC_18_7_7 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_0_5_LC_18_7_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_0_5_LC_18_7_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_0_5_LC_18_7_7  (
            .in0(N__32391),
            .in1(N__29097),
            .in2(_gnd_net_),
            .in3(N__32083),
            .lcout(\b2v_inst.N_267 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_0_cry_0_c_inv_LC_18_8_0 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_0_cry_0_c_inv_LC_18_8_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_0_cry_0_c_inv_LC_18_8_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final4_0_cry_0_c_inv_LC_18_8_0  (
            .in0(N__29664),
            .in1(N__29065),
            .in2(N__29022),
            .in3(_gnd_net_),
            .lcout(\b2v_inst.reg_ancho_3_i_0 ),
            .ltout(),
            .carryin(bfn_18_8_0_),
            .carryout(\b2v_inst.valor_max_final4_0_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_0_cry_1_c_inv_LC_18_8_1 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_0_cry_1_c_inv_LC_18_8_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_0_cry_1_c_inv_LC_18_8_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final4_0_cry_1_c_inv_LC_18_8_1  (
            .in0(_gnd_net_),
            .in1(N__28990),
            .in2(N__28944),
            .in3(N__29691),
            .lcout(\b2v_inst.reg_ancho_3_i_1 ),
            .ltout(),
            .carryin(\b2v_inst.valor_max_final4_0_cry_0 ),
            .carryout(\b2v_inst.valor_max_final4_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_0_cry_2_c_inv_LC_18_8_2 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_0_cry_2_c_inv_LC_18_8_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_0_cry_2_c_inv_LC_18_8_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final4_0_cry_2_c_inv_LC_18_8_2  (
            .in0(_gnd_net_),
            .in1(N__31245),
            .in2(N__28911),
            .in3(N__32153),
            .lcout(\b2v_inst.reg_ancho_3_i_2 ),
            .ltout(),
            .carryin(\b2v_inst.valor_max_final4_0_cry_1 ),
            .carryout(\b2v_inst.valor_max_final4_0_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_0_cry_3_c_inv_LC_18_8_3 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_0_cry_3_c_inv_LC_18_8_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_0_cry_3_c_inv_LC_18_8_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final4_0_cry_3_c_inv_LC_18_8_3  (
            .in0(N__32230),
            .in1(N__31037),
            .in2(N__28881),
            .in3(_gnd_net_),
            .lcout(\b2v_inst.reg_ancho_3_i_3 ),
            .ltout(),
            .carryin(\b2v_inst.valor_max_final4_0_cry_2 ),
            .carryout(\b2v_inst.valor_max_final4_0_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_0_cry_4_c_inv_LC_18_8_4 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_0_cry_4_c_inv_LC_18_8_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_0_cry_4_c_inv_LC_18_8_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final4_0_cry_4_c_inv_LC_18_8_4  (
            .in0(_gnd_net_),
            .in1(N__29635),
            .in2(N__29589),
            .in3(N__31426),
            .lcout(\b2v_inst.reg_ancho_3_i_4 ),
            .ltout(),
            .carryin(\b2v_inst.valor_max_final4_0_cry_3 ),
            .carryout(\b2v_inst.valor_max_final4_0_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_0_cry_5_c_inv_LC_18_8_5 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_0_cry_5_c_inv_LC_18_8_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_0_cry_5_c_inv_LC_18_8_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final4_0_cry_5_c_inv_LC_18_8_5  (
            .in0(_gnd_net_),
            .in1(N__29505),
            .in2(N__29561),
            .in3(N__32082),
            .lcout(\b2v_inst.reg_ancho_3_i_5 ),
            .ltout(),
            .carryin(\b2v_inst.valor_max_final4_0_cry_4 ),
            .carryout(\b2v_inst.valor_max_final4_0_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_0_cry_6_c_inv_LC_18_8_6 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_0_cry_6_c_inv_LC_18_8_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_0_cry_6_c_inv_LC_18_8_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final4_0_cry_6_c_inv_LC_18_8_6  (
            .in0(_gnd_net_),
            .in1(N__29484),
            .in2(N__29424),
            .in3(N__29442),
            .lcout(\b2v_inst.reg_ancho_3_i_6 ),
            .ltout(),
            .carryin(\b2v_inst.valor_max_final4_0_cry_5 ),
            .carryout(\b2v_inst.valor_max_final4_0_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_0_cry_7_c_inv_LC_18_8_7 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_0_cry_7_c_inv_LC_18_8_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_0_cry_7_c_inv_LC_18_8_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final4_0_cry_7_c_inv_LC_18_8_7  (
            .in0(_gnd_net_),
            .in1(N__29391),
            .in2(N__29349),
            .in3(N__30690),
            .lcout(\b2v_inst.reg_ancho_3_i_7 ),
            .ltout(),
            .carryin(\b2v_inst.valor_max_final4_0_cry_6 ),
            .carryout(\b2v_inst.valor_max_final4_0_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_0_cry_8_c_inv_LC_18_9_0 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_0_cry_8_c_inv_LC_18_9_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_0_cry_8_c_inv_LC_18_9_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final4_0_cry_8_c_inv_LC_18_9_0  (
            .in0(N__30724),
            .in1(N__29964),
            .in2(N__29319),
            .in3(_gnd_net_),
            .lcout(\b2v_inst.reg_ancho_3_i_8 ),
            .ltout(),
            .carryin(bfn_18_9_0_),
            .carryout(\b2v_inst.valor_max_final4_0_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_0_cry_9_c_inv_LC_18_9_1 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_0_cry_9_c_inv_LC_18_9_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_0_cry_9_c_inv_LC_18_9_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final4_0_cry_9_c_inv_LC_18_9_1  (
            .in0(_gnd_net_),
            .in1(N__30004),
            .in2(N__29286),
            .in3(N__30132),
            .lcout(\b2v_inst.reg_ancho_3_i_9 ),
            .ltout(),
            .carryin(\b2v_inst.valor_max_final4_0_cry_8 ),
            .carryout(\b2v_inst.valor_max_final4_0_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_0_cry_10_c_inv_LC_18_9_2 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_0_cry_10_c_inv_LC_18_9_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final4_0_cry_10_c_inv_LC_18_9_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final4_0_cry_10_c_inv_LC_18_9_2  (
            .in0(_gnd_net_),
            .in1(N__29256),
            .in2(N__29208),
            .in3(N__32301),
            .lcout(\b2v_inst.reg_ancho_3_i_10 ),
            .ltout(),
            .carryin(\b2v_inst.valor_max_final4_0_cry_9 ),
            .carryout(\b2v_inst.valor_max_final40 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.valor_max_final40_THRU_LUT4_0_LC_18_9_3 .C_ON=1'b0;
    defparam \b2v_inst.valor_max_final40_THRU_LUT4_0_LC_18_9_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.valor_max_final40_THRU_LUT4_0_LC_18_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.valor_max_final40_THRU_LUT4_0_LC_18_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29180),
            .lcout(\b2v_inst.valor_max_final40_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_0_9_LC_18_9_4 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_0_9_LC_18_9_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_0_9_LC_18_9_4 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_0_9_LC_18_9_4  (
            .in0(N__32546),
            .in1(_gnd_net_),
            .in2(N__29741),
            .in3(N__30005),
            .lcout(\b2v_inst.N_543 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_0_8_LC_18_9_5 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_0_8_LC_18_9_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_0_8_LC_18_9_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_0_8_LC_18_9_5  (
            .in0(N__29965),
            .in1(N__29925),
            .in2(_gnd_net_),
            .in3(N__32545),
            .lcout(\b2v_inst.N_542 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_1_3_LC_18_9_6 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_1_3_LC_18_9_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_1_3_LC_18_9_6 .LUT_INIT=16'b0100110001111111;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_1_3_LC_18_9_6  (
            .in0(N__30971),
            .in1(N__31180),
            .in2(N__29873),
            .in3(N__32465),
            .lcout(\b2v_inst.un1_reg_anterior_0_i_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_0_2_LC_18_9_7 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_0_2_LC_18_9_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_0_2_LC_18_9_7 .LUT_INIT=16'b0101111100111111;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_0_2_LC_18_9_7  (
            .in0(N__29838),
            .in1(N__32152),
            .in2(N__30989),
            .in3(N__32397),
            .lcout(\b2v_inst.data_a_escribir_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir11_6_c_RNO_LC_18_10_0 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir11_6_c_RNO_LC_18_10_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir11_6_c_RNO_LC_18_10_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst.data_a_escribir11_6_c_RNO_LC_18_10_0  (
            .in0(N__31438),
            .in1(N__32229),
            .in2(N__32084),
            .in3(N__32151),
            .lcout(\b2v_inst.data_a_escribir11_6_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_1_5_LC_18_10_1 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_1_5_LC_18_10_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_1_5_LC_18_10_1 .LUT_INIT=16'b1111000011110001;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_1_5_LC_18_10_1  (
            .in0(N__31177),
            .in1(N__29789),
            .in2(N__29774),
            .in3(N__30627),
            .lcout(),
            .ltout(\b2v_inst.un1_reg_anterior_iv_0_1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_5_LC_18_10_2 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_5_LC_18_10_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.data_a_escribir_5_LC_18_10_2 .LUT_INIT=16'b0000111100001101;
    LogicCell40 \b2v_inst.data_a_escribir_5_LC_18_10_2  (
            .in0(N__30629),
            .in1(N__29765),
            .in2(N__29753),
            .in3(N__31179),
            .lcout(b2v_inst_data_a_escribir_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34381),
            .ce(N__30555),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_2_LC_18_10_6 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_2_LC_18_10_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.data_a_escribir_2_LC_18_10_6 .LUT_INIT=16'b0001001111001110;
    LogicCell40 \b2v_inst.data_a_escribir_2_LC_18_10_6  (
            .in0(N__30628),
            .in1(N__31178),
            .in2(N__29750),
            .in3(N__31049),
            .lcout(b2v_inst_data_a_escribir_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34381),
            .ce(N__30555),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir11_5_c_RNO_LC_18_11_0 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir11_5_c_RNO_LC_18_11_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir11_5_c_RNO_LC_18_11_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst.data_a_escribir11_5_c_RNO_LC_18_11_0  (
            .in0(N__29736),
            .in1(N__29702),
            .in2(N__31488),
            .in3(N__29675),
            .lcout(\b2v_inst.data_a_escribir11_5_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_2_9_LC_18_11_2 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_2_9_LC_18_11_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_2_9_LC_18_11_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_2_9_LC_18_11_2  (
            .in0(N__31954),
            .in1(N__30137),
            .in2(_gnd_net_),
            .in3(N__32407),
            .lcout(\b2v_inst.N_545 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_3_9_LC_18_11_3 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_3_9_LC_18_11_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_3_9_LC_18_11_3 .LUT_INIT=16'b0111011100110011;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_3_9_LC_18_11_3  (
            .in0(N__30110),
            .in1(N__30957),
            .in2(_gnd_net_),
            .in3(N__31168),
            .lcout(),
            .ltout(\b2v_inst.un1_reg_anterior_iv_0_0_0_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_1_9_LC_18_11_4 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_1_9_LC_18_11_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_1_9_LC_18_11_4 .LUT_INIT=16'b1111000111110000;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_1_9_LC_18_11_4  (
            .in0(N__31169),
            .in1(N__30095),
            .in2(N__30089),
            .in3(N__30609),
            .lcout(),
            .ltout(\b2v_inst.un1_reg_anterior_iv_0_0_1_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_9_LC_18_11_5 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_9_LC_18_11_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.data_a_escribir_9_LC_18_11_5 .LUT_INIT=16'b0000111100001110;
    LogicCell40 \b2v_inst.data_a_escribir_9_LC_18_11_5  (
            .in0(N__30611),
            .in1(N__30086),
            .in2(N__30077),
            .in3(N__31171),
            .lcout(b2v_inst_data_a_escribir_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34378),
            .ce(N__30557),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_6_LC_18_11_7 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_6_LC_18_11_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.data_a_escribir_6_LC_18_11_7 .LUT_INIT=16'b0000000011111101;
    LogicCell40 \b2v_inst.data_a_escribir_6_LC_18_11_7  (
            .in0(N__30610),
            .in1(N__31170),
            .in2(N__30074),
            .in3(N__30059),
            .lcout(b2v_inst_data_a_escribir_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34378),
            .ce(N__30557),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir11_10_c_RNO_LC_18_12_0 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir11_10_c_RNO_LC_18_12_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir11_10_c_RNO_LC_18_12_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst.data_a_escribir11_10_c_RNO_LC_18_12_0  (
            .in0(N__31946),
            .in1(N__30768),
            .in2(N__31730),
            .in3(N__30670),
            .lcout(\b2v_inst.data_a_escribir11_10_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_3_8_LC_18_12_1 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_3_8_LC_18_12_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_3_8_LC_18_12_1 .LUT_INIT=16'b0111011100110011;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_3_8_LC_18_12_1  (
            .in0(N__30038),
            .in1(N__30990),
            .in2(_gnd_net_),
            .in3(N__31172),
            .lcout(),
            .ltout(\b2v_inst.un1_reg_anterior_iv_0_0_0_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_1_8_LC_18_12_2 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_1_8_LC_18_12_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_1_8_LC_18_12_2 .LUT_INIT=16'b1111000111110000;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_1_8_LC_18_12_2  (
            .in0(N__31173),
            .in1(N__30704),
            .in2(N__30020),
            .in3(N__30622),
            .lcout(),
            .ltout(\b2v_inst.un1_reg_anterior_iv_0_0_1_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_8_LC_18_12_3 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_8_LC_18_12_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.data_a_escribir_8_LC_18_12_3 .LUT_INIT=16'b0000111100001110;
    LogicCell40 \b2v_inst.data_a_escribir_8_LC_18_12_3  (
            .in0(N__30623),
            .in1(N__30017),
            .in2(N__30008),
            .in3(N__31175),
            .lcout(b2v_inst_data_a_escribir_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34382),
            .ce(N__30554),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_2_8_LC_18_12_4 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_2_8_LC_18_12_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_2_8_LC_18_12_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_2_8_LC_18_12_4  (
            .in0(N__30769),
            .in1(N__30728),
            .in2(_gnd_net_),
            .in3(N__32395),
            .lcout(\b2v_inst.N_544 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_0_7_LC_18_12_5 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_0_7_LC_18_12_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_0_7_LC_18_12_5 .LUT_INIT=16'b0001101111111111;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_0_7_LC_18_12_5  (
            .in0(N__32396),
            .in1(N__30698),
            .in2(N__30674),
            .in3(N__30991),
            .lcout(),
            .ltout(\b2v_inst.data_a_escribir_RNO_0Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_7_LC_18_12_6 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_7_LC_18_12_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.data_a_escribir_7_LC_18_12_6 .LUT_INIT=16'b0010011101100110;
    LogicCell40 \b2v_inst.data_a_escribir_7_LC_18_12_6  (
            .in0(N__31174),
            .in1(N__30638),
            .in2(N__30632),
            .in3(N__30624),
            .lcout(b2v_inst_data_a_escribir_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34382),
            .ce(N__30554),
            .sr(_gnd_net_));
    defparam \b2v_inst9.cycle_counter_2_LC_18_13_0 .C_ON=1'b0;
    defparam \b2v_inst9.cycle_counter_2_LC_18_13_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst9.cycle_counter_2_LC_18_13_0 .LUT_INIT=16'b0000001000100000;
    LogicCell40 \b2v_inst9.cycle_counter_2_LC_18_13_0  (
            .in0(N__30467),
            .in1(N__38155),
            .in2(N__30497),
            .in3(N__30503),
            .lcout(\b2v_inst9.cycle_counterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34392),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst9.cycle_counter_0_LC_18_13_1 .C_ON=1'b0;
    defparam \b2v_inst9.cycle_counter_0_LC_18_13_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst9.cycle_counter_0_LC_18_13_1 .LUT_INIT=16'b0000010000001000;
    LogicCell40 \b2v_inst9.cycle_counter_0_LC_18_13_1  (
            .in0(N__30302),
            .in1(N__30466),
            .in2(N__38156),
            .in3(N__30433),
            .lcout(\b2v_inst9.cycle_counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34392),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.pix_data_reg_3_LC_18_14_5 .C_ON=1'b0;
    defparam \b2v_inst.pix_data_reg_3_LC_18_14_5 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.pix_data_reg_3_LC_18_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.pix_data_reg_3_LC_18_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30281),
            .lcout(\b2v_inst.pix_data_regZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34398),
            .ce(N__30248),
            .sr(N__38131));
    defparam \b2v_inst.cantidad_temp_2_LC_18_15_6 .C_ON=1'b0;
    defparam \b2v_inst.cantidad_temp_2_LC_18_15_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.cantidad_temp_2_LC_18_15_6 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \b2v_inst.cantidad_temp_2_LC_18_15_6  (
            .in0(N__34765),
            .in1(N__32656),
            .in2(N__30191),
            .in3(N__34642),
            .lcout(b2v_inst_cantidad_temp_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34409),
            .ce(),
            .sr(N__38137));
    defparam \b2v_inst.reg_anterior_4_LC_19_6_0 .C_ON=1'b0;
    defparam \b2v_inst.reg_anterior_4_LC_19_6_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_anterior_4_LC_19_6_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \b2v_inst.reg_anterior_4_LC_19_6_0  (
            .in0(_gnd_net_),
            .in1(N__31917),
            .in2(_gnd_net_),
            .in3(N__33050),
            .lcout(\b2v_inst.reg_anteriorZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34410),
            .ce(N__31673),
            .sr(N__38138));
    defparam \b2v_inst.reg_anterior_6_LC_19_6_7 .C_ON=1'b0;
    defparam \b2v_inst.reg_anterior_6_LC_19_6_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_anterior_6_LC_19_6_7 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \b2v_inst.reg_anterior_6_LC_19_6_7  (
            .in0(N__31918),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31562),
            .lcout(\b2v_inst.reg_anteriorZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34410),
            .ce(N__31673),
            .sr(N__38138));
    defparam \b2v_inst.reg_ancho_2_10_LC_19_7_7 .C_ON=1'b0;
    defparam \b2v_inst.reg_ancho_2_10_LC_19_7_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_ancho_2_10_LC_19_7_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.reg_ancho_2_10_LC_19_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31780),
            .lcout(\b2v_inst.reg_ancho_2Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34399),
            .ce(N__32959),
            .sr(N__38132));
    defparam \b2v_inst.reg_ancho_3_4_LC_19_8_7 .C_ON=1'b0;
    defparam \b2v_inst.reg_ancho_3_4_LC_19_8_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_ancho_3_4_LC_19_8_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \b2v_inst.reg_ancho_3_4_LC_19_8_7  (
            .in0(_gnd_net_),
            .in1(N__31902),
            .in2(_gnd_net_),
            .in3(N__33061),
            .lcout(\b2v_inst.reg_ancho_3Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34393),
            .ce(N__32059),
            .sr(N__38124));
    defparam \b2v_inst.data_a_escribir11_3_c_RNO_LC_19_9_0 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir11_3_c_RNO_LC_19_9_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir11_3_c_RNO_LC_19_9_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst.data_a_escribir11_3_c_RNO_LC_19_9_0  (
            .in0(N__32434),
            .in1(N__31282),
            .in2(N__33010),
            .in3(N__31330),
            .lcout(\b2v_inst.data_a_escribir11_3_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.reg_ancho_2_1_LC_19_9_1 .C_ON=1'b0;
    defparam \b2v_inst.reg_ancho_2_1_LC_19_9_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_ancho_2_1_LC_19_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.reg_ancho_2_1_LC_19_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31395),
            .lcout(\b2v_inst.reg_ancho_2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34383),
            .ce(N__32965),
            .sr(N__38118));
    defparam \b2v_inst.reg_ancho_2_2_LC_19_9_2 .C_ON=1'b0;
    defparam \b2v_inst.reg_ancho_2_2_LC_19_9_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_ancho_2_2_LC_19_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.reg_ancho_2_2_LC_19_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32209),
            .lcout(\b2v_inst.reg_ancho_2Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34383),
            .ce(N__32965),
            .sr(N__38118));
    defparam \b2v_inst.data_a_escribir_RNO_2_2_LC_19_9_3 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_2_2_LC_19_9_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_2_2_LC_19_9_3 .LUT_INIT=16'b0101111100111111;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_2_2_LC_19_9_3  (
            .in0(N__31283),
            .in1(N__31255),
            .in2(N__30979),
            .in3(N__32544),
            .lcout(),
            .ltout(\b2v_inst.data_a_escribir_RNO_2Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_1_2_LC_19_9_4 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_1_2_LC_19_9_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_1_2_LC_19_9_4 .LUT_INIT=16'b0111011100001111;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_1_2_LC_19_9_4  (
            .in0(N__31202),
            .in1(N__30941),
            .in2(N__31184),
            .in3(N__31181),
            .lcout(\b2v_inst.un1_reg_anterior_0_i_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_2_3_LC_19_9_5 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_2_3_LC_19_9_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_2_3_LC_19_9_5 .LUT_INIT=16'b0101111100111111;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_2_3_LC_19_9_5  (
            .in0(N__32438),
            .in1(N__31043),
            .in2(N__30978),
            .in3(N__32543),
            .lcout(\b2v_inst.data_a_escribir_RNO_2Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.reg_ancho_2_3_LC_19_9_7 .C_ON=1'b0;
    defparam \b2v_inst.reg_ancho_2_3_LC_19_9_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_ancho_2_3_LC_19_9_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.reg_ancho_2_3_LC_19_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32283),
            .lcout(\b2v_inst.reg_ancho_2Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34383),
            .ce(N__32965),
            .sr(N__38118));
    defparam \b2v_inst.data_a_escribir_RNO_0_10_LC_19_10_1 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_0_10_LC_19_10_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_0_10_LC_19_10_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_0_10_LC_19_10_1  (
            .in0(N__31718),
            .in1(N__32305),
            .in2(_gnd_net_),
            .in3(N__32394),
            .lcout(\b2v_inst.N_264 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.reg_ancho_3_10_LC_19_10_2 .C_ON=1'b0;
    defparam \b2v_inst.reg_ancho_3_10_LC_19_10_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_ancho_3_10_LC_19_10_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \b2v_inst.reg_ancho_3_10_LC_19_10_2  (
            .in0(_gnd_net_),
            .in1(N__31898),
            .in2(_gnd_net_),
            .in3(N__31776),
            .lcout(\b2v_inst.reg_ancho_3Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34379),
            .ce(N__32052),
            .sr(N__38108));
    defparam \b2v_inst.reg_ancho_3_3_LC_19_10_3 .C_ON=1'b0;
    defparam \b2v_inst.reg_ancho_3_3_LC_19_10_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_ancho_3_3_LC_19_10_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \b2v_inst.reg_ancho_3_3_LC_19_10_3  (
            .in0(N__31900),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32284),
            .lcout(\b2v_inst.reg_ancho_3Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34379),
            .ce(N__32052),
            .sr(N__38108));
    defparam \b2v_inst.reg_ancho_3_2_LC_19_10_4 .C_ON=1'b0;
    defparam \b2v_inst.reg_ancho_3_2_LC_19_10_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_ancho_3_2_LC_19_10_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \b2v_inst.reg_ancho_3_2_LC_19_10_4  (
            .in0(_gnd_net_),
            .in1(N__31899),
            .in2(_gnd_net_),
            .in3(N__32205),
            .lcout(\b2v_inst.reg_ancho_3Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34379),
            .ce(N__32052),
            .sr(N__38108));
    defparam \b2v_inst.reg_ancho_3_5_LC_19_10_5 .C_ON=1'b0;
    defparam \b2v_inst.reg_ancho_3_5_LC_19_10_5 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_ancho_3_5_LC_19_10_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \b2v_inst.reg_ancho_3_5_LC_19_10_5  (
            .in0(N__31901),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32131),
            .lcout(\b2v_inst.reg_ancho_3Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34379),
            .ce(N__32052),
            .sr(N__38108));
    defparam \b2v_inst.reg_anterior_9_LC_19_11_0 .C_ON=1'b0;
    defparam \b2v_inst.reg_anterior_9_LC_19_11_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_anterior_9_LC_19_11_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \b2v_inst.reg_anterior_9_LC_19_11_0  (
            .in0(N__31897),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31985),
            .lcout(\b2v_inst.reg_anteriorZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34373),
            .ce(N__31688),
            .sr(N__38119));
    defparam \b2v_inst.reg_anterior_10_LC_19_11_1 .C_ON=1'b0;
    defparam \b2v_inst.reg_anterior_10_LC_19_11_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_anterior_10_LC_19_11_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \b2v_inst.reg_anterior_10_LC_19_11_1  (
            .in0(_gnd_net_),
            .in1(N__31896),
            .in2(_gnd_net_),
            .in3(N__31772),
            .lcout(\b2v_inst.reg_anteriorZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34373),
            .ce(N__31688),
            .sr(N__38119));
    defparam \b2v_inst.cantidad_temp_0_LC_19_13_3 .C_ON=1'b0;
    defparam \b2v_inst.cantidad_temp_0_LC_19_13_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.cantidad_temp_0_LC_19_13_3 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \b2v_inst.cantidad_temp_0_LC_19_13_3  (
            .in0(N__34908),
            .in1(N__34627),
            .in2(N__32705),
            .in3(N__34762),
            .lcout(b2v_inst_cantidad_temp_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34384),
            .ce(),
            .sr(N__38133));
    defparam \b2v_inst.cantidad_temp_1_LC_19_13_4 .C_ON=1'b0;
    defparam \b2v_inst.cantidad_temp_1_LC_19_13_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.cantidad_temp_1_LC_19_13_4 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \b2v_inst.cantidad_temp_1_LC_19_13_4  (
            .in0(N__34628),
            .in1(N__34870),
            .in2(N__32690),
            .in3(N__34764),
            .lcout(b2v_inst_cantidad_temp_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34384),
            .ce(),
            .sr(N__38133));
    defparam \b2v_inst.cantidad_temp_4_LC_19_13_7 .C_ON=1'b0;
    defparam \b2v_inst.cantidad_temp_4_LC_19_13_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.cantidad_temp_4_LC_19_13_7 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \b2v_inst.cantidad_temp_4_LC_19_13_7  (
            .in0(N__32623),
            .in1(N__34629),
            .in2(N__32678),
            .in3(N__34763),
            .lcout(b2v_inst_cantidad_temp_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34384),
            .ce(),
            .sr(N__38133));
    defparam \b2v_inst.un16_data_ram_cantidad_o_cry_1_c_LC_19_14_0 .C_ON=1'b1;
    defparam \b2v_inst.un16_data_ram_cantidad_o_cry_1_c_LC_19_14_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un16_data_ram_cantidad_o_cry_1_c_LC_19_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.un16_data_ram_cantidad_o_cry_1_c_LC_19_14_0  (
            .in0(_gnd_net_),
            .in1(N__34865),
            .in2(N__34909),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_19_14_0_),
            .carryout(\b2v_inst.un16_data_ram_cantidad_o_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un16_data_ram_cantidad_o_cry_1_c_RNI77CO_LC_19_14_1 .C_ON=1'b1;
    defparam \b2v_inst.un16_data_ram_cantidad_o_cry_1_c_RNI77CO_LC_19_14_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un16_data_ram_cantidad_o_cry_1_c_RNI77CO_LC_19_14_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.un16_data_ram_cantidad_o_cry_1_c_RNI77CO_LC_19_14_1  (
            .in0(_gnd_net_),
            .in1(N__32652),
            .in2(_gnd_net_),
            .in3(N__32636),
            .lcout(\b2v_inst.un16_data_ram_cantidad_o_cry_1_c_RNI77COZ0 ),
            .ltout(),
            .carryin(\b2v_inst.un16_data_ram_cantidad_o_cry_1 ),
            .carryout(\b2v_inst.un16_data_ram_cantidad_o_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un16_data_ram_cantidad_o_cry_2_c_RNI9ADO_LC_19_14_2 .C_ON=1'b1;
    defparam \b2v_inst.un16_data_ram_cantidad_o_cry_2_c_RNI9ADO_LC_19_14_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un16_data_ram_cantidad_o_cry_2_c_RNI9ADO_LC_19_14_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.un16_data_ram_cantidad_o_cry_2_c_RNI9ADO_LC_19_14_2  (
            .in0(_gnd_net_),
            .in1(N__34545),
            .in2(_gnd_net_),
            .in3(N__32633),
            .lcout(\b2v_inst.un16_data_ram_cantidad_o_cry_2_c_RNI9ADOZ0 ),
            .ltout(),
            .carryin(\b2v_inst.un16_data_ram_cantidad_o_cry_2 ),
            .carryout(\b2v_inst.un16_data_ram_cantidad_o_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un16_data_ram_cantidad_o_cry_3_c_RNIBDEO_LC_19_14_3 .C_ON=1'b1;
    defparam \b2v_inst.un16_data_ram_cantidad_o_cry_3_c_RNIBDEO_LC_19_14_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un16_data_ram_cantidad_o_cry_3_c_RNIBDEO_LC_19_14_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.un16_data_ram_cantidad_o_cry_3_c_RNIBDEO_LC_19_14_3  (
            .in0(_gnd_net_),
            .in1(N__32619),
            .in2(_gnd_net_),
            .in3(N__32603),
            .lcout(\b2v_inst.un16_data_ram_cantidad_o_cry_3_c_RNIBDEOZ0 ),
            .ltout(),
            .carryin(\b2v_inst.un16_data_ram_cantidad_o_cry_3 ),
            .carryout(\b2v_inst.un16_data_ram_cantidad_o_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un16_data_ram_cantidad_o_cry_4_c_RNIDGFO_LC_19_14_4 .C_ON=1'b0;
    defparam \b2v_inst.un16_data_ram_cantidad_o_cry_4_c_RNIDGFO_LC_19_14_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un16_data_ram_cantidad_o_cry_4_c_RNIDGFO_LC_19_14_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \b2v_inst.un16_data_ram_cantidad_o_cry_4_c_RNIDGFO_LC_19_14_4  (
            .in0(_gnd_net_),
            .in1(N__32599),
            .in2(_gnd_net_),
            .in3(N__32567),
            .lcout(\b2v_inst.un16_data_ram_cantidad_o_cry_4_c_RNIDGFOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNIH17G1_2_LC_19_14_5 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNIH17G1_2_LC_19_14_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNIH17G1_2_LC_19_14_5 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \b2v_inst.data_a_escribir_RNIH17G1_2_LC_19_14_5  (
            .in0(N__37792),
            .in1(N__32564),
            .in2(N__33140),
            .in3(N__37547),
            .lcout(N_553_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNIN99G1_4_LC_19_15_4 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNIN99G1_4_LC_19_15_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNIN99G1_4_LC_19_15_4 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \b2v_inst.data_a_escribir_RNIN99G1_4_LC_19_15_4  (
            .in0(N__37808),
            .in1(N__33347),
            .in2(N__33329),
            .in3(N__37530),
            .lcout(N_549_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNIK58G1_3_LC_19_15_6 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNIK58G1_3_LC_19_15_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNIK58G1_3_LC_19_15_6 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \b2v_inst.data_a_escribir_RNIK58G1_3_LC_19_15_6  (
            .in0(N__37807),
            .in1(N__33263),
            .in2(N__33257),
            .in3(N__37531),
            .lcout(N_551_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNIHBT91_10_LC_19_16_1 .C_ON=1'b0;
    defparam \b2v_inst.state_RNIHBT91_10_LC_19_16_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNIHBT91_10_LC_19_16_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \b2v_inst.state_RNIHBT91_10_LC_19_16_1  (
            .in0(_gnd_net_),
            .in1(N__35196),
            .in2(_gnd_net_),
            .in3(N__33188),
            .lcout(\b2v_inst.N_645 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNI8OQN_0_LC_20_3_7 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNI8OQN_0_LC_20_3_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNI8OQN_0_LC_20_3_7 .LUT_INIT=16'b0010001010101010;
    LogicCell40 \b2v_inst.data_a_escribir_RNI8OQN_0_LC_20_3_7  (
            .in0(N__34976),
            .in1(N__37841),
            .in2(_gnd_net_),
            .in3(N__37561),
            .lcout(N_121_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNIAQQN_2_LC_20_6_3 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNIAQQN_2_LC_20_6_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNIAQQN_2_LC_20_6_3 .LUT_INIT=16'b0010001010101010;
    LogicCell40 \b2v_inst.data_a_escribir_RNIAQQN_2_LC_20_6_3  (
            .in0(N__33124),
            .in1(N__37836),
            .in2(_gnd_net_),
            .in3(N__37562),
            .lcout(N_118_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.reg_ancho_2_4_LC_20_8_0 .C_ON=1'b0;
    defparam \b2v_inst.reg_ancho_2_4_LC_20_8_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_ancho_2_4_LC_20_8_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.reg_ancho_2_4_LC_20_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33054),
            .lcout(\b2v_inst.reg_ancho_2Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34385),
            .ce(N__32966),
            .sr(N__38134));
    defparam \b2v_inst.data_a_escribir_RNIH1RN_9_LC_20_9_4 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNIH1RN_9_LC_20_9_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNIH1RN_9_LC_20_9_4 .LUT_INIT=16'b0010001010101010;
    LogicCell40 \b2v_inst.data_a_escribir_RNIH1RN_9_LC_20_9_4  (
            .in0(N__32859),
            .in1(N__37823),
            .in2(_gnd_net_),
            .in3(N__37497),
            .lcout(N_111_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_RNI1E333_6_LC_20_10_0 .C_ON=1'b0;
    defparam \b2v_inst.indice_RNI1E333_6_LC_20_10_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_RNI1E333_6_LC_20_10_0 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \b2v_inst.indice_RNI1E333_6_LC_20_10_0  (
            .in0(N__32819),
            .in1(N__38377),
            .in2(N__32801),
            .in3(N__35240),
            .lcout(N_298),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_RNIS8333_5_LC_20_10_1 .C_ON=1'b0;
    defparam \b2v_inst.indice_RNIS8333_5_LC_20_10_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_RNIS8333_5_LC_20_10_1 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \b2v_inst.indice_RNIS8333_5_LC_20_10_1  (
            .in0(N__35243),
            .in1(N__34046),
            .in2(N__34031),
            .in3(N__35726),
            .lcout(indice_RNIS8333_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_RNIBO333_8_LC_20_10_5 .C_ON=1'b0;
    defparam \b2v_inst.indice_RNIBO333_8_LC_20_10_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_RNIBO333_8_LC_20_10_5 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \b2v_inst.indice_RNIBO333_8_LC_20_10_5  (
            .in0(N__35241),
            .in1(N__33929),
            .in2(N__33911),
            .in3(N__39081),
            .lcout(indice_RNIBO333_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_RNIGT333_9_LC_20_10_6 .C_ON=1'b0;
    defparam \b2v_inst.indice_RNIGT333_9_LC_20_10_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_RNIGT333_9_LC_20_10_6 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \b2v_inst.indice_RNIGT333_9_LC_20_10_6  (
            .in0(N__33812),
            .in1(N__35953),
            .in2(N__33797),
            .in3(N__35242),
            .lcout(indice_RNIGT333_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNIDTQN_5_LC_20_11_1 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNIDTQN_5_LC_20_11_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNIDTQN_5_LC_20_11_1 .LUT_INIT=16'b0010101000101010;
    LogicCell40 \b2v_inst.data_a_escribir_RNIDTQN_5_LC_20_11_1  (
            .in0(N__37598),
            .in1(N__37819),
            .in2(N__37560),
            .in3(_gnd_net_),
            .lcout(N_115_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNIPNGN_10_LC_20_11_4 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNIPNGN_10_LC_20_11_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNIPNGN_10_LC_20_11_4 .LUT_INIT=16'b0011111100000000;
    LogicCell40 \b2v_inst.data_a_escribir_RNIPNGN_10_LC_20_11_4  (
            .in0(_gnd_net_),
            .in1(N__37550),
            .in2(N__37835),
            .in3(N__33669),
            .lcout(N_110_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_RNI3F233_0_LC_20_11_6 .C_ON=1'b0;
    defparam \b2v_inst.indice_RNI3F233_0_LC_20_11_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_RNI3F233_0_LC_20_11_6 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \b2v_inst.indice_RNI3F233_0_LC_20_11_6  (
            .in0(N__33620),
            .in1(N__35238),
            .in2(N__33605),
            .in3(N__39318),
            .lcout(indice_RNI3F233_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_RNIO3V73_10_LC_20_11_7 .C_ON=1'b0;
    defparam \b2v_inst.indice_RNIO3V73_10_LC_20_11_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_RNIO3V73_10_LC_20_11_7 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \b2v_inst.indice_RNIO3V73_10_LC_20_11_7  (
            .in0(N__35239),
            .in1(N__33512),
            .in2(N__33494),
            .in3(N__36751),
            .lcout(N_37),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNIG0RN_8_LC_20_12_0 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNIG0RN_8_LC_20_12_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNIG0RN_8_LC_20_12_0 .LUT_INIT=16'b0101111100000000;
    LogicCell40 \b2v_inst.data_a_escribir_RNIG0RN_8_LC_20_12_0  (
            .in0(N__37544),
            .in1(_gnd_net_),
            .in2(N__37840),
            .in3(N__33381),
            .lcout(N_112_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNIFVQN_7_LC_20_12_1 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNIFVQN_7_LC_20_12_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNIFVQN_7_LC_20_12_1 .LUT_INIT=16'b0010001010101010;
    LogicCell40 \b2v_inst.data_a_escribir_RNIFVQN_7_LC_20_12_1  (
            .in0(N__35484),
            .in1(N__37831),
            .in2(_gnd_net_),
            .in3(N__37543),
            .lcout(N_113_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_RNI8K233_1_LC_20_12_5 .C_ON=1'b0;
    defparam \b2v_inst.indice_RNI8K233_1_LC_20_12_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_RNI8K233_1_LC_20_12_5 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \b2v_inst.indice_RNI8K233_1_LC_20_12_5  (
            .in0(N__35450),
            .in1(N__35209),
            .in2(N__35432),
            .in3(N__38660),
            .lcout(indice_RNI8K233_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNIEUQN_6_LC_20_13_2 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNIEUQN_6_LC_20_13_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNIEUQN_6_LC_20_13_2 .LUT_INIT=16'b0010001010101010;
    LogicCell40 \b2v_inst.data_a_escribir_RNIEUQN_6_LC_20_13_2  (
            .in0(N__35315),
            .in1(N__37809),
            .in2(_gnd_net_),
            .in3(N__37545),
            .lcout(N_114_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_RNIDP233_2_LC_20_13_4 .C_ON=1'b0;
    defparam \b2v_inst.indice_RNIDP233_2_LC_20_13_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_RNIDP233_2_LC_20_13_4 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \b2v_inst.indice_RNIDP233_2_LC_20_13_4  (
            .in0(N__35258),
            .in1(N__35208),
            .in2(N__35075),
            .in3(N__36122),
            .lcout(indice_RNIDP233_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNIIIS11_0_LC_20_13_7 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNIIIS11_0_LC_20_13_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNIIIS11_0_LC_20_13_7 .LUT_INIT=16'b0000100001011101;
    LogicCell40 \b2v_inst.data_a_escribir_RNIIIS11_0_LC_20_13_7  (
            .in0(N__37546),
            .in1(N__34975),
            .in2(N__37830),
            .in3(N__34907),
            .lcout(N_557_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.cantidad_temp_RNILL3K_1_LC_20_14_0 .C_ON=1'b0;
    defparam \b2v_inst.cantidad_temp_RNILL3K_1_LC_20_14_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.cantidad_temp_RNILL3K_1_LC_20_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst.cantidad_temp_RNILL3K_1_LC_20_14_0  (
            .in0(_gnd_net_),
            .in1(N__34903),
            .in2(_gnd_net_),
            .in3(N__34866),
            .lcout(),
            .ltout(\b2v_inst.cantidad_temp_RNILL3KZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNIUEUB1_1_LC_20_14_1 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNIUEUB1_1_LC_20_14_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNIUEUB1_1_LC_20_14_1 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \b2v_inst.data_a_escribir_RNIUEUB1_1_LC_20_14_1  (
            .in0(N__34840),
            .in1(N__37549),
            .in2(N__34775),
            .in3(N__37793),
            .lcout(N_555_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.cantidad_temp_3_LC_20_14_6 .C_ON=1'b0;
    defparam \b2v_inst.cantidad_temp_3_LC_20_14_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.cantidad_temp_3_LC_20_14_6 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \b2v_inst.cantidad_temp_3_LC_20_14_6  (
            .in0(N__34549),
            .in1(N__34766),
            .in2(N__34652),
            .in3(N__34643),
            .lcout(b2v_inst_cantidad_temp_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34386),
            .ce(),
            .sr(N__38139));
    defparam \b2v_inst.data_a_escribir_RNIQDAG1_5_LC_20_15_4 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNIQDAG1_5_LC_20_15_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNIQDAG1_5_LC_20_15_4 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \b2v_inst.data_a_escribir_RNIQDAG1_5_LC_20_15_4  (
            .in0(N__37813),
            .in1(N__37637),
            .in2(N__37627),
            .in3(N__37548),
            .lcout(N_547_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_20_15_5.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_20_15_5.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_20_15_5.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_20_15_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_energia_RNIFL4P2_10_LC_20_16_0 .C_ON=1'b0;
    defparam \b2v_inst.dir_energia_RNIFL4P2_10_LC_20_16_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_energia_RNIFL4P2_10_LC_20_16_0 .LUT_INIT=16'b0100010001010000;
    LogicCell40 \b2v_inst.dir_energia_RNIFL4P2_10_LC_20_16_0  (
            .in0(N__38458),
            .in1(N__36788),
            .in2(N__36752),
            .in3(N__38242),
            .lcout(N_445_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_energia_RNIJFLU2_3_LC_20_16_1 .C_ON=1'b0;
    defparam \b2v_inst.dir_energia_RNIJFLU2_3_LC_20_16_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_energia_RNIJFLU2_3_LC_20_16_1 .LUT_INIT=16'b0011000000100010;
    LogicCell40 \b2v_inst.dir_energia_RNIJFLU2_3_LC_20_16_1  (
            .in0(N__36581),
            .in1(N__38460),
            .in2(N__36467),
            .in3(N__38246),
            .lcout(N_357_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_energia_RNILHLU2_4_LC_20_16_2 .C_ON=1'b0;
    defparam \b2v_inst.dir_energia_RNILHLU2_4_LC_20_16_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_energia_RNILHLU2_4_LC_20_16_2 .LUT_INIT=16'b0101000001000100;
    LogicCell40 \b2v_inst.dir_energia_RNILHLU2_4_LC_20_16_2  (
            .in0(N__38461),
            .in1(N__36376),
            .in2(N__36257),
            .in3(N__38244),
            .lcout(N_356_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_energia_RNIHDLU2_2_LC_20_16_4 .C_ON=1'b0;
    defparam \b2v_inst.dir_energia_RNIHDLU2_2_LC_20_16_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_energia_RNIHDLU2_2_LC_20_16_4 .LUT_INIT=16'b0101000101000000;
    LogicCell40 \b2v_inst.dir_energia_RNIHDLU2_2_LC_20_16_4  (
            .in0(N__38459),
            .in1(N__38243),
            .in2(N__36164),
            .in3(N__36121),
            .lcout(N_358_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_energia_RNIVRLU2_9_LC_20_16_6 .C_ON=1'b0;
    defparam \b2v_inst.dir_energia_RNIVRLU2_9_LC_20_16_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_energia_RNIVRLU2_9_LC_20_16_6 .LUT_INIT=16'b0101000001000100;
    LogicCell40 \b2v_inst.dir_energia_RNIVRLU2_9_LC_20_16_6  (
            .in0(N__38463),
            .in1(N__35933),
            .in2(N__35831),
            .in3(N__38245),
            .lcout(N_444_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_energia_RNINJLU2_5_LC_20_16_7 .C_ON=1'b0;
    defparam \b2v_inst.dir_energia_RNINJLU2_5_LC_20_16_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_energia_RNINJLU2_5_LC_20_16_7 .LUT_INIT=16'b0011000000100010;
    LogicCell40 \b2v_inst.dir_energia_RNINJLU2_5_LC_20_16_7  (
            .in0(N__35722),
            .in1(N__38462),
            .in2(N__35594),
            .in3(N__38247),
            .lcout(N_355_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_energia_RNID9LU2_0_LC_20_17_0 .C_ON=1'b0;
    defparam \b2v_inst.dir_energia_RNID9LU2_0_LC_20_17_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_energia_RNID9LU2_0_LC_20_17_0 .LUT_INIT=16'b0101000101000000;
    LogicCell40 \b2v_inst.dir_energia_RNID9LU2_0_LC_20_17_0  (
            .in0(N__38464),
            .in1(N__38260),
            .in2(N__39383),
            .in3(N__39323),
            .lcout(N_360_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_energia_RNITPLU2_8_LC_20_17_2 .C_ON=1'b0;
    defparam \b2v_inst.dir_energia_RNITPLU2_8_LC_20_17_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_energia_RNITPLU2_8_LC_20_17_2 .LUT_INIT=16'b0100010001010000;
    LogicCell40 \b2v_inst.dir_energia_RNITPLU2_8_LC_20_17_2  (
            .in0(N__38468),
            .in1(N__39146),
            .in2(N__39100),
            .in3(N__38264),
            .lcout(N_443_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_energia_RNIRNLU2_7_LC_20_17_3 .C_ON=1'b0;
    defparam \b2v_inst.dir_energia_RNIRNLU2_7_LC_20_17_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_energia_RNIRNLU2_7_LC_20_17_3 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \b2v_inst.dir_energia_RNIRNLU2_7_LC_20_17_3  (
            .in0(N__38263),
            .in1(N__38467),
            .in2(N__38927),
            .in3(N__38866),
            .lcout(N_353_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_energia_RNIFBLU2_1_LC_20_17_4 .C_ON=1'b0;
    defparam \b2v_inst.dir_energia_RNIFBLU2_1_LC_20_17_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_energia_RNIFBLU2_1_LC_20_17_4 .LUT_INIT=16'b0101000101000000;
    LogicCell40 \b2v_inst.dir_energia_RNIFBLU2_1_LC_20_17_4  (
            .in0(N__38465),
            .in1(N__38261),
            .in2(N__38714),
            .in3(N__38666),
            .lcout(N_359_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_energia_RNIPLLU2_6_LC_20_17_6 .C_ON=1'b0;
    defparam \b2v_inst.dir_energia_RNIPLLU2_6_LC_20_17_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_energia_RNIPLLU2_6_LC_20_17_6 .LUT_INIT=16'b0100010001010000;
    LogicCell40 \b2v_inst.dir_energia_RNIPLLU2_6_LC_20_17_6  (
            .in0(N__38466),
            .in1(N__38429),
            .in2(N__38381),
            .in3(N__38262),
            .lcout(N_354_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // anda_plis_2
