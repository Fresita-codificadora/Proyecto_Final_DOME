// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Oct 3 2024 21:30:24

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "anda_plis" view "INTERFACE"

module anda_plis (
    uart_tx_o,
    uart_rx_i,
    reset,
    clk);

    output uart_tx_o;
    input uart_rx_i;
    input reset;
    input clk;

    wire N__24159;
    wire N__24158;
    wire N__24157;
    wire N__24150;
    wire N__24149;
    wire N__24148;
    wire N__24141;
    wire N__24140;
    wire N__24139;
    wire N__24132;
    wire N__24131;
    wire N__24130;
    wire N__24113;
    wire N__24110;
    wire N__24107;
    wire N__24104;
    wire N__24101;
    wire N__24098;
    wire N__24095;
    wire N__24094;
    wire N__24093;
    wire N__24092;
    wire N__24089;
    wire N__24086;
    wire N__24083;
    wire N__24082;
    wire N__24081;
    wire N__24078;
    wire N__24073;
    wire N__24070;
    wire N__24067;
    wire N__24064;
    wire N__24063;
    wire N__24060;
    wire N__24057;
    wire N__24054;
    wire N__24051;
    wire N__24048;
    wire N__24045;
    wire N__24042;
    wire N__24037;
    wire N__24032;
    wire N__24029;
    wire N__24020;
    wire N__24019;
    wire N__24018;
    wire N__24017;
    wire N__24016;
    wire N__24015;
    wire N__24014;
    wire N__24011;
    wire N__24006;
    wire N__24005;
    wire N__24004;
    wire N__24003;
    wire N__23998;
    wire N__23993;
    wire N__23992;
    wire N__23991;
    wire N__23990;
    wire N__23989;
    wire N__23988;
    wire N__23987;
    wire N__23986;
    wire N__23985;
    wire N__23984;
    wire N__23981;
    wire N__23978;
    wire N__23973;
    wire N__23970;
    wire N__23965;
    wire N__23960;
    wire N__23957;
    wire N__23950;
    wire N__23947;
    wire N__23942;
    wire N__23921;
    wire N__23920;
    wire N__23919;
    wire N__23918;
    wire N__23917;
    wire N__23916;
    wire N__23915;
    wire N__23914;
    wire N__23913;
    wire N__23912;
    wire N__23911;
    wire N__23910;
    wire N__23905;
    wire N__23904;
    wire N__23903;
    wire N__23902;
    wire N__23901;
    wire N__23900;
    wire N__23897;
    wire N__23894;
    wire N__23891;
    wire N__23886;
    wire N__23883;
    wire N__23878;
    wire N__23873;
    wire N__23870;
    wire N__23863;
    wire N__23858;
    wire N__23837;
    wire N__23836;
    wire N__23835;
    wire N__23834;
    wire N__23833;
    wire N__23832;
    wire N__23831;
    wire N__23830;
    wire N__23829;
    wire N__23824;
    wire N__23823;
    wire N__23822;
    wire N__23821;
    wire N__23820;
    wire N__23815;
    wire N__23810;
    wire N__23809;
    wire N__23804;
    wire N__23801;
    wire N__23798;
    wire N__23793;
    wire N__23790;
    wire N__23787;
    wire N__23782;
    wire N__23779;
    wire N__23762;
    wire N__23759;
    wire N__23756;
    wire N__23755;
    wire N__23754;
    wire N__23753;
    wire N__23750;
    wire N__23749;
    wire N__23748;
    wire N__23743;
    wire N__23742;
    wire N__23741;
    wire N__23740;
    wire N__23739;
    wire N__23738;
    wire N__23735;
    wire N__23730;
    wire N__23729;
    wire N__23728;
    wire N__23727;
    wire N__23724;
    wire N__23721;
    wire N__23718;
    wire N__23715;
    wire N__23712;
    wire N__23709;
    wire N__23708;
    wire N__23707;
    wire N__23706;
    wire N__23705;
    wire N__23704;
    wire N__23703;
    wire N__23700;
    wire N__23695;
    wire N__23690;
    wire N__23685;
    wire N__23682;
    wire N__23679;
    wire N__23672;
    wire N__23667;
    wire N__23664;
    wire N__23661;
    wire N__23656;
    wire N__23647;
    wire N__23630;
    wire N__23629;
    wire N__23626;
    wire N__23625;
    wire N__23624;
    wire N__23623;
    wire N__23622;
    wire N__23621;
    wire N__23620;
    wire N__23619;
    wire N__23618;
    wire N__23617;
    wire N__23614;
    wire N__23613;
    wire N__23612;
    wire N__23609;
    wire N__23608;
    wire N__23607;
    wire N__23604;
    wire N__23603;
    wire N__23600;
    wire N__23599;
    wire N__23598;
    wire N__23595;
    wire N__23594;
    wire N__23593;
    wire N__23592;
    wire N__23591;
    wire N__23590;
    wire N__23589;
    wire N__23588;
    wire N__23583;
    wire N__23574;
    wire N__23571;
    wire N__23566;
    wire N__23563;
    wire N__23558;
    wire N__23553;
    wire N__23550;
    wire N__23545;
    wire N__23540;
    wire N__23533;
    wire N__23526;
    wire N__23519;
    wire N__23498;
    wire N__23497;
    wire N__23496;
    wire N__23495;
    wire N__23494;
    wire N__23491;
    wire N__23490;
    wire N__23489;
    wire N__23488;
    wire N__23485;
    wire N__23484;
    wire N__23483;
    wire N__23482;
    wire N__23479;
    wire N__23476;
    wire N__23475;
    wire N__23474;
    wire N__23471;
    wire N__23468;
    wire N__23465;
    wire N__23462;
    wire N__23459;
    wire N__23456;
    wire N__23455;
    wire N__23452;
    wire N__23449;
    wire N__23446;
    wire N__23445;
    wire N__23442;
    wire N__23439;
    wire N__23436;
    wire N__23433;
    wire N__23430;
    wire N__23427;
    wire N__23420;
    wire N__23417;
    wire N__23412;
    wire N__23409;
    wire N__23406;
    wire N__23403;
    wire N__23398;
    wire N__23395;
    wire N__23392;
    wire N__23379;
    wire N__23366;
    wire N__23365;
    wire N__23362;
    wire N__23359;
    wire N__23354;
    wire N__23351;
    wire N__23348;
    wire N__23347;
    wire N__23346;
    wire N__23345;
    wire N__23344;
    wire N__23343;
    wire N__23342;
    wire N__23341;
    wire N__23336;
    wire N__23333;
    wire N__23330;
    wire N__23327;
    wire N__23324;
    wire N__23321;
    wire N__23320;
    wire N__23317;
    wire N__23316;
    wire N__23315;
    wire N__23314;
    wire N__23313;
    wire N__23310;
    wire N__23305;
    wire N__23302;
    wire N__23301;
    wire N__23296;
    wire N__23295;
    wire N__23294;
    wire N__23291;
    wire N__23286;
    wire N__23285;
    wire N__23282;
    wire N__23279;
    wire N__23276;
    wire N__23271;
    wire N__23268;
    wire N__23265;
    wire N__23262;
    wire N__23255;
    wire N__23252;
    wire N__23249;
    wire N__23238;
    wire N__23225;
    wire N__23222;
    wire N__23219;
    wire N__23218;
    wire N__23217;
    wire N__23216;
    wire N__23215;
    wire N__23212;
    wire N__23211;
    wire N__23210;
    wire N__23207;
    wire N__23206;
    wire N__23203;
    wire N__23202;
    wire N__23201;
    wire N__23200;
    wire N__23199;
    wire N__23196;
    wire N__23195;
    wire N__23192;
    wire N__23185;
    wire N__23182;
    wire N__23177;
    wire N__23176;
    wire N__23175;
    wire N__23174;
    wire N__23173;
    wire N__23168;
    wire N__23167;
    wire N__23166;
    wire N__23163;
    wire N__23158;
    wire N__23153;
    wire N__23152;
    wire N__23149;
    wire N__23144;
    wire N__23135;
    wire N__23134;
    wire N__23131;
    wire N__23126;
    wire N__23119;
    wire N__23116;
    wire N__23113;
    wire N__23110;
    wire N__23107;
    wire N__23104;
    wire N__23097;
    wire N__23084;
    wire N__23083;
    wire N__23082;
    wire N__23081;
    wire N__23078;
    wire N__23077;
    wire N__23076;
    wire N__23071;
    wire N__23068;
    wire N__23065;
    wire N__23064;
    wire N__23063;
    wire N__23060;
    wire N__23059;
    wire N__23058;
    wire N__23055;
    wire N__23054;
    wire N__23051;
    wire N__23048;
    wire N__23045;
    wire N__23038;
    wire N__23037;
    wire N__23036;
    wire N__23029;
    wire N__23028;
    wire N__23027;
    wire N__23024;
    wire N__23023;
    wire N__23022;
    wire N__23021;
    wire N__23012;
    wire N__23007;
    wire N__23004;
    wire N__22997;
    wire N__22996;
    wire N__22991;
    wire N__22988;
    wire N__22985;
    wire N__22982;
    wire N__22977;
    wire N__22974;
    wire N__22969;
    wire N__22966;
    wire N__22961;
    wire N__22952;
    wire N__22951;
    wire N__22950;
    wire N__22949;
    wire N__22948;
    wire N__22947;
    wire N__22946;
    wire N__22945;
    wire N__22928;
    wire N__22925;
    wire N__22922;
    wire N__22921;
    wire N__22920;
    wire N__22919;
    wire N__22918;
    wire N__22917;
    wire N__22916;
    wire N__22915;
    wire N__22914;
    wire N__22913;
    wire N__22912;
    wire N__22911;
    wire N__22910;
    wire N__22909;
    wire N__22908;
    wire N__22907;
    wire N__22906;
    wire N__22905;
    wire N__22904;
    wire N__22903;
    wire N__22902;
    wire N__22901;
    wire N__22900;
    wire N__22899;
    wire N__22898;
    wire N__22897;
    wire N__22896;
    wire N__22895;
    wire N__22894;
    wire N__22893;
    wire N__22892;
    wire N__22891;
    wire N__22890;
    wire N__22889;
    wire N__22888;
    wire N__22887;
    wire N__22886;
    wire N__22885;
    wire N__22884;
    wire N__22883;
    wire N__22882;
    wire N__22881;
    wire N__22880;
    wire N__22879;
    wire N__22878;
    wire N__22877;
    wire N__22876;
    wire N__22875;
    wire N__22778;
    wire N__22775;
    wire N__22772;
    wire N__22769;
    wire N__22766;
    wire N__22763;
    wire N__22760;
    wire N__22757;
    wire N__22754;
    wire N__22751;
    wire N__22750;
    wire N__22749;
    wire N__22748;
    wire N__22747;
    wire N__22746;
    wire N__22743;
    wire N__22740;
    wire N__22737;
    wire N__22734;
    wire N__22733;
    wire N__22730;
    wire N__22727;
    wire N__22724;
    wire N__22715;
    wire N__22710;
    wire N__22709;
    wire N__22708;
    wire N__22705;
    wire N__22700;
    wire N__22699;
    wire N__22698;
    wire N__22695;
    wire N__22694;
    wire N__22691;
    wire N__22690;
    wire N__22689;
    wire N__22686;
    wire N__22683;
    wire N__22680;
    wire N__22679;
    wire N__22676;
    wire N__22673;
    wire N__22670;
    wire N__22667;
    wire N__22664;
    wire N__22661;
    wire N__22658;
    wire N__22655;
    wire N__22650;
    wire N__22647;
    wire N__22642;
    wire N__22637;
    wire N__22634;
    wire N__22631;
    wire N__22624;
    wire N__22621;
    wire N__22618;
    wire N__22607;
    wire N__22606;
    wire N__22605;
    wire N__22602;
    wire N__22599;
    wire N__22598;
    wire N__22597;
    wire N__22596;
    wire N__22595;
    wire N__22594;
    wire N__22593;
    wire N__22590;
    wire N__22589;
    wire N__22588;
    wire N__22587;
    wire N__22582;
    wire N__22579;
    wire N__22578;
    wire N__22577;
    wire N__22574;
    wire N__22573;
    wire N__22572;
    wire N__22571;
    wire N__22570;
    wire N__22569;
    wire N__22566;
    wire N__22565;
    wire N__22564;
    wire N__22563;
    wire N__22562;
    wire N__22561;
    wire N__22558;
    wire N__22555;
    wire N__22554;
    wire N__22551;
    wire N__22550;
    wire N__22547;
    wire N__22544;
    wire N__22541;
    wire N__22538;
    wire N__22533;
    wire N__22530;
    wire N__22527;
    wire N__22524;
    wire N__22521;
    wire N__22518;
    wire N__22517;
    wire N__22516;
    wire N__22515;
    wire N__22514;
    wire N__22511;
    wire N__22510;
    wire N__22509;
    wire N__22506;
    wire N__22503;
    wire N__22502;
    wire N__22501;
    wire N__22500;
    wire N__22497;
    wire N__22496;
    wire N__22493;
    wire N__22490;
    wire N__22487;
    wire N__22484;
    wire N__22483;
    wire N__22482;
    wire N__22481;
    wire N__22480;
    wire N__22477;
    wire N__22472;
    wire N__22469;
    wire N__22468;
    wire N__22465;
    wire N__22462;
    wire N__22461;
    wire N__22456;
    wire N__22455;
    wire N__22454;
    wire N__22453;
    wire N__22448;
    wire N__22447;
    wire N__22444;
    wire N__22439;
    wire N__22432;
    wire N__22429;
    wire N__22426;
    wire N__22423;
    wire N__22420;
    wire N__22419;
    wire N__22416;
    wire N__22413;
    wire N__22412;
    wire N__22411;
    wire N__22410;
    wire N__22407;
    wire N__22406;
    wire N__22405;
    wire N__22402;
    wire N__22399;
    wire N__22396;
    wire N__22393;
    wire N__22392;
    wire N__22389;
    wire N__22388;
    wire N__22385;
    wire N__22382;
    wire N__22381;
    wire N__22380;
    wire N__22377;
    wire N__22374;
    wire N__22371;
    wire N__22368;
    wire N__22365;
    wire N__22362;
    wire N__22359;
    wire N__22356;
    wire N__22355;
    wire N__22354;
    wire N__22353;
    wire N__22352;
    wire N__22351;
    wire N__22348;
    wire N__22343;
    wire N__22340;
    wire N__22335;
    wire N__22332;
    wire N__22329;
    wire N__22326;
    wire N__22323;
    wire N__22320;
    wire N__22319;
    wire N__22318;
    wire N__22315;
    wire N__22312;
    wire N__22297;
    wire N__22294;
    wire N__22291;
    wire N__22288;
    wire N__22285;
    wire N__22282;
    wire N__22281;
    wire N__22280;
    wire N__22277;
    wire N__22274;
    wire N__22271;
    wire N__22268;
    wire N__22267;
    wire N__22264;
    wire N__22263;
    wire N__22256;
    wire N__22253;
    wire N__22252;
    wire N__22251;
    wire N__22248;
    wire N__22245;
    wire N__22244;
    wire N__22243;
    wire N__22242;
    wire N__22237;
    wire N__22234;
    wire N__22231;
    wire N__22230;
    wire N__22219;
    wire N__22216;
    wire N__22213;
    wire N__22210;
    wire N__22207;
    wire N__22204;
    wire N__22201;
    wire N__22198;
    wire N__22195;
    wire N__22188;
    wire N__22187;
    wire N__22182;
    wire N__22177;
    wire N__22174;
    wire N__22171;
    wire N__22168;
    wire N__22165;
    wire N__22162;
    wire N__22155;
    wire N__22150;
    wire N__22145;
    wire N__22142;
    wire N__22139;
    wire N__22136;
    wire N__22129;
    wire N__22126;
    wire N__22123;
    wire N__22120;
    wire N__22115;
    wire N__22114;
    wire N__22111;
    wire N__22108;
    wire N__22103;
    wire N__22102;
    wire N__22099;
    wire N__22096;
    wire N__22093;
    wire N__22090;
    wire N__22085;
    wire N__22084;
    wire N__22083;
    wire N__22082;
    wire N__22081;
    wire N__22078;
    wire N__22075;
    wire N__22072;
    wire N__22069;
    wire N__22064;
    wire N__22053;
    wire N__22050;
    wire N__22047;
    wire N__22044;
    wire N__22035;
    wire N__22030;
    wire N__22021;
    wire N__22014;
    wire N__22009;
    wire N__22006;
    wire N__22003;
    wire N__21998;
    wire N__21995;
    wire N__21992;
    wire N__21989;
    wire N__21986;
    wire N__21983;
    wire N__21978;
    wire N__21975;
    wire N__21972;
    wire N__21971;
    wire N__21968;
    wire N__21965;
    wire N__21964;
    wire N__21961;
    wire N__21948;
    wire N__21947;
    wire N__21946;
    wire N__21945;
    wire N__21940;
    wire N__21937;
    wire N__21932;
    wire N__21923;
    wire N__21916;
    wire N__21905;
    wire N__21902;
    wire N__21899;
    wire N__21894;
    wire N__21891;
    wire N__21890;
    wire N__21885;
    wire N__21884;
    wire N__21881;
    wire N__21878;
    wire N__21875;
    wire N__21874;
    wire N__21871;
    wire N__21866;
    wire N__21861;
    wire N__21850;
    wire N__21847;
    wire N__21844;
    wire N__21841;
    wire N__21838;
    wire N__21833;
    wire N__21830;
    wire N__21827;
    wire N__21824;
    wire N__21821;
    wire N__21818;
    wire N__21811;
    wire N__21804;
    wire N__21801;
    wire N__21798;
    wire N__21793;
    wire N__21788;
    wire N__21785;
    wire N__21782;
    wire N__21779;
    wire N__21776;
    wire N__21767;
    wire N__21766;
    wire N__21763;
    wire N__21760;
    wire N__21757;
    wire N__21752;
    wire N__21749;
    wire N__21748;
    wire N__21747;
    wire N__21742;
    wire N__21739;
    wire N__21734;
    wire N__21733;
    wire N__21732;
    wire N__21729;
    wire N__21726;
    wire N__21725;
    wire N__21724;
    wire N__21723;
    wire N__21720;
    wire N__21715;
    wire N__21712;
    wire N__21709;
    wire N__21706;
    wire N__21695;
    wire N__21694;
    wire N__21693;
    wire N__21692;
    wire N__21691;
    wire N__21690;
    wire N__21689;
    wire N__21686;
    wire N__21681;
    wire N__21678;
    wire N__21675;
    wire N__21670;
    wire N__21667;
    wire N__21666;
    wire N__21663;
    wire N__21662;
    wire N__21661;
    wire N__21660;
    wire N__21659;
    wire N__21658;
    wire N__21657;
    wire N__21656;
    wire N__21653;
    wire N__21650;
    wire N__21647;
    wire N__21644;
    wire N__21643;
    wire N__21640;
    wire N__21639;
    wire N__21636;
    wire N__21633;
    wire N__21626;
    wire N__21623;
    wire N__21620;
    wire N__21617;
    wire N__21612;
    wire N__21607;
    wire N__21600;
    wire N__21581;
    wire N__21578;
    wire N__21575;
    wire N__21572;
    wire N__21569;
    wire N__21566;
    wire N__21563;
    wire N__21562;
    wire N__21561;
    wire N__21560;
    wire N__21559;
    wire N__21556;
    wire N__21553;
    wire N__21552;
    wire N__21549;
    wire N__21544;
    wire N__21543;
    wire N__21542;
    wire N__21539;
    wire N__21534;
    wire N__21533;
    wire N__21532;
    wire N__21531;
    wire N__21530;
    wire N__21529;
    wire N__21528;
    wire N__21527;
    wire N__21522;
    wire N__21517;
    wire N__21512;
    wire N__21507;
    wire N__21500;
    wire N__21495;
    wire N__21482;
    wire N__21479;
    wire N__21478;
    wire N__21477;
    wire N__21476;
    wire N__21473;
    wire N__21468;
    wire N__21467;
    wire N__21464;
    wire N__21463;
    wire N__21462;
    wire N__21457;
    wire N__21456;
    wire N__21455;
    wire N__21454;
    wire N__21453;
    wire N__21450;
    wire N__21445;
    wire N__21444;
    wire N__21443;
    wire N__21440;
    wire N__21439;
    wire N__21436;
    wire N__21431;
    wire N__21426;
    wire N__21421;
    wire N__21416;
    wire N__21411;
    wire N__21404;
    wire N__21395;
    wire N__21392;
    wire N__21389;
    wire N__21386;
    wire N__21383;
    wire N__21380;
    wire N__21377;
    wire N__21374;
    wire N__21371;
    wire N__21368;
    wire N__21365;
    wire N__21362;
    wire N__21359;
    wire N__21356;
    wire N__21355;
    wire N__21354;
    wire N__21353;
    wire N__21352;
    wire N__21351;
    wire N__21348;
    wire N__21345;
    wire N__21342;
    wire N__21339;
    wire N__21336;
    wire N__21333;
    wire N__21330;
    wire N__21327;
    wire N__21324;
    wire N__21311;
    wire N__21310;
    wire N__21305;
    wire N__21302;
    wire N__21299;
    wire N__21296;
    wire N__21293;
    wire N__21290;
    wire N__21287;
    wire N__21284;
    wire N__21281;
    wire N__21278;
    wire N__21275;
    wire N__21272;
    wire N__21269;
    wire N__21266;
    wire N__21265;
    wire N__21262;
    wire N__21261;
    wire N__21258;
    wire N__21255;
    wire N__21252;
    wire N__21251;
    wire N__21248;
    wire N__21243;
    wire N__21240;
    wire N__21233;
    wire N__21232;
    wire N__21229;
    wire N__21226;
    wire N__21225;
    wire N__21224;
    wire N__21223;
    wire N__21222;
    wire N__21221;
    wire N__21220;
    wire N__21215;
    wire N__21210;
    wire N__21207;
    wire N__21206;
    wire N__21205;
    wire N__21204;
    wire N__21197;
    wire N__21190;
    wire N__21183;
    wire N__21176;
    wire N__21175;
    wire N__21174;
    wire N__21173;
    wire N__21172;
    wire N__21165;
    wire N__21162;
    wire N__21159;
    wire N__21158;
    wire N__21157;
    wire N__21156;
    wire N__21155;
    wire N__21152;
    wire N__21147;
    wire N__21146;
    wire N__21145;
    wire N__21142;
    wire N__21135;
    wire N__21134;
    wire N__21133;
    wire N__21128;
    wire N__21125;
    wire N__21122;
    wire N__21119;
    wire N__21116;
    wire N__21111;
    wire N__21106;
    wire N__21095;
    wire N__21094;
    wire N__21093;
    wire N__21092;
    wire N__21091;
    wire N__21090;
    wire N__21087;
    wire N__21086;
    wire N__21085;
    wire N__21084;
    wire N__21083;
    wire N__21080;
    wire N__21077;
    wire N__21072;
    wire N__21069;
    wire N__21066;
    wire N__21063;
    wire N__21060;
    wire N__21059;
    wire N__21058;
    wire N__21053;
    wire N__21046;
    wire N__21039;
    wire N__21038;
    wire N__21035;
    wire N__21032;
    wire N__21029;
    wire N__21024;
    wire N__21021;
    wire N__21018;
    wire N__21005;
    wire N__21004;
    wire N__21003;
    wire N__21002;
    wire N__20997;
    wire N__20994;
    wire N__20991;
    wire N__20990;
    wire N__20987;
    wire N__20984;
    wire N__20981;
    wire N__20978;
    wire N__20975;
    wire N__20972;
    wire N__20969;
    wire N__20966;
    wire N__20957;
    wire N__20954;
    wire N__20953;
    wire N__20950;
    wire N__20947;
    wire N__20944;
    wire N__20941;
    wire N__20936;
    wire N__20935;
    wire N__20934;
    wire N__20933;
    wire N__20932;
    wire N__20929;
    wire N__20928;
    wire N__20927;
    wire N__20924;
    wire N__20921;
    wire N__20918;
    wire N__20915;
    wire N__20914;
    wire N__20913;
    wire N__20912;
    wire N__20909;
    wire N__20906;
    wire N__20903;
    wire N__20900;
    wire N__20899;
    wire N__20898;
    wire N__20897;
    wire N__20890;
    wire N__20883;
    wire N__20878;
    wire N__20873;
    wire N__20872;
    wire N__20869;
    wire N__20868;
    wire N__20867;
    wire N__20862;
    wire N__20857;
    wire N__20852;
    wire N__20847;
    wire N__20842;
    wire N__20831;
    wire N__20828;
    wire N__20827;
    wire N__20826;
    wire N__20825;
    wire N__20824;
    wire N__20823;
    wire N__20822;
    wire N__20815;
    wire N__20812;
    wire N__20809;
    wire N__20804;
    wire N__20801;
    wire N__20798;
    wire N__20797;
    wire N__20792;
    wire N__20789;
    wire N__20786;
    wire N__20783;
    wire N__20780;
    wire N__20777;
    wire N__20768;
    wire N__20765;
    wire N__20764;
    wire N__20763;
    wire N__20760;
    wire N__20757;
    wire N__20756;
    wire N__20755;
    wire N__20754;
    wire N__20751;
    wire N__20748;
    wire N__20745;
    wire N__20742;
    wire N__20737;
    wire N__20734;
    wire N__20723;
    wire N__20722;
    wire N__20719;
    wire N__20716;
    wire N__20713;
    wire N__20712;
    wire N__20711;
    wire N__20710;
    wire N__20707;
    wire N__20704;
    wire N__20699;
    wire N__20696;
    wire N__20687;
    wire N__20686;
    wire N__20685;
    wire N__20682;
    wire N__20677;
    wire N__20674;
    wire N__20671;
    wire N__20666;
    wire N__20665;
    wire N__20664;
    wire N__20661;
    wire N__20658;
    wire N__20653;
    wire N__20650;
    wire N__20647;
    wire N__20642;
    wire N__20639;
    wire N__20638;
    wire N__20637;
    wire N__20636;
    wire N__20635;
    wire N__20634;
    wire N__20633;
    wire N__20632;
    wire N__20631;
    wire N__20630;
    wire N__20627;
    wire N__20624;
    wire N__20621;
    wire N__20618;
    wire N__20617;
    wire N__20614;
    wire N__20611;
    wire N__20610;
    wire N__20605;
    wire N__20604;
    wire N__20603;
    wire N__20600;
    wire N__20597;
    wire N__20588;
    wire N__20585;
    wire N__20580;
    wire N__20579;
    wire N__20578;
    wire N__20577;
    wire N__20576;
    wire N__20573;
    wire N__20570;
    wire N__20565;
    wire N__20562;
    wire N__20561;
    wire N__20558;
    wire N__20557;
    wire N__20550;
    wire N__20547;
    wire N__20540;
    wire N__20531;
    wire N__20528;
    wire N__20525;
    wire N__20522;
    wire N__20519;
    wire N__20504;
    wire N__20503;
    wire N__20502;
    wire N__20501;
    wire N__20500;
    wire N__20495;
    wire N__20494;
    wire N__20493;
    wire N__20492;
    wire N__20489;
    wire N__20486;
    wire N__20485;
    wire N__20484;
    wire N__20483;
    wire N__20482;
    wire N__20479;
    wire N__20478;
    wire N__20477;
    wire N__20476;
    wire N__20473;
    wire N__20468;
    wire N__20465;
    wire N__20462;
    wire N__20459;
    wire N__20454;
    wire N__20453;
    wire N__20448;
    wire N__20445;
    wire N__20442;
    wire N__20441;
    wire N__20436;
    wire N__20425;
    wire N__20422;
    wire N__20419;
    wire N__20416;
    wire N__20411;
    wire N__20408;
    wire N__20407;
    wire N__20406;
    wire N__20405;
    wire N__20404;
    wire N__20403;
    wire N__20402;
    wire N__20399;
    wire N__20394;
    wire N__20391;
    wire N__20384;
    wire N__20375;
    wire N__20370;
    wire N__20367;
    wire N__20354;
    wire N__20351;
    wire N__20348;
    wire N__20345;
    wire N__20342;
    wire N__20339;
    wire N__20336;
    wire N__20333;
    wire N__20332;
    wire N__20331;
    wire N__20330;
    wire N__20329;
    wire N__20328;
    wire N__20327;
    wire N__20326;
    wire N__20325;
    wire N__20324;
    wire N__20323;
    wire N__20320;
    wire N__20317;
    wire N__20312;
    wire N__20309;
    wire N__20304;
    wire N__20299;
    wire N__20298;
    wire N__20297;
    wire N__20296;
    wire N__20295;
    wire N__20294;
    wire N__20291;
    wire N__20286;
    wire N__20281;
    wire N__20278;
    wire N__20277;
    wire N__20276;
    wire N__20271;
    wire N__20266;
    wire N__20257;
    wire N__20254;
    wire N__20249;
    wire N__20246;
    wire N__20243;
    wire N__20242;
    wire N__20239;
    wire N__20234;
    wire N__20227;
    wire N__20222;
    wire N__20213;
    wire N__20210;
    wire N__20207;
    wire N__20204;
    wire N__20201;
    wire N__20198;
    wire N__20195;
    wire N__20192;
    wire N__20189;
    wire N__20186;
    wire N__20183;
    wire N__20180;
    wire N__20179;
    wire N__20176;
    wire N__20173;
    wire N__20168;
    wire N__20165;
    wire N__20162;
    wire N__20159;
    wire N__20156;
    wire N__20153;
    wire N__20150;
    wire N__20147;
    wire N__20146;
    wire N__20143;
    wire N__20142;
    wire N__20141;
    wire N__20140;
    wire N__20139;
    wire N__20136;
    wire N__20133;
    wire N__20128;
    wire N__20125;
    wire N__20124;
    wire N__20123;
    wire N__20118;
    wire N__20117;
    wire N__20116;
    wire N__20115;
    wire N__20114;
    wire N__20113;
    wire N__20110;
    wire N__20107;
    wire N__20106;
    wire N__20103;
    wire N__20098;
    wire N__20097;
    wire N__20096;
    wire N__20095;
    wire N__20094;
    wire N__20093;
    wire N__20090;
    wire N__20085;
    wire N__20082;
    wire N__20077;
    wire N__20072;
    wire N__20069;
    wire N__20064;
    wire N__20059;
    wire N__20054;
    wire N__20051;
    wire N__20048;
    wire N__20027;
    wire N__20024;
    wire N__20021;
    wire N__20020;
    wire N__20019;
    wire N__20016;
    wire N__20013;
    wire N__20010;
    wire N__20007;
    wire N__20000;
    wire N__19997;
    wire N__19994;
    wire N__19991;
    wire N__19988;
    wire N__19985;
    wire N__19982;
    wire N__19979;
    wire N__19976;
    wire N__19973;
    wire N__19970;
    wire N__19967;
    wire N__19964;
    wire N__19963;
    wire N__19962;
    wire N__19961;
    wire N__19952;
    wire N__19949;
    wire N__19946;
    wire N__19943;
    wire N__19940;
    wire N__19937;
    wire N__19934;
    wire N__19933;
    wire N__19930;
    wire N__19927;
    wire N__19926;
    wire N__19921;
    wire N__19920;
    wire N__19917;
    wire N__19914;
    wire N__19911;
    wire N__19908;
    wire N__19905;
    wire N__19900;
    wire N__19895;
    wire N__19894;
    wire N__19891;
    wire N__19890;
    wire N__19889;
    wire N__19886;
    wire N__19883;
    wire N__19880;
    wire N__19877;
    wire N__19876;
    wire N__19875;
    wire N__19874;
    wire N__19873;
    wire N__19870;
    wire N__19869;
    wire N__19866;
    wire N__19863;
    wire N__19862;
    wire N__19857;
    wire N__19852;
    wire N__19849;
    wire N__19846;
    wire N__19843;
    wire N__19838;
    wire N__19835;
    wire N__19830;
    wire N__19817;
    wire N__19816;
    wire N__19815;
    wire N__19812;
    wire N__19809;
    wire N__19808;
    wire N__19807;
    wire N__19806;
    wire N__19805;
    wire N__19804;
    wire N__19801;
    wire N__19798;
    wire N__19795;
    wire N__19792;
    wire N__19789;
    wire N__19786;
    wire N__19781;
    wire N__19778;
    wire N__19773;
    wire N__19760;
    wire N__19759;
    wire N__19758;
    wire N__19757;
    wire N__19756;
    wire N__19755;
    wire N__19754;
    wire N__19751;
    wire N__19744;
    wire N__19741;
    wire N__19740;
    wire N__19735;
    wire N__19728;
    wire N__19727;
    wire N__19726;
    wire N__19725;
    wire N__19724;
    wire N__19723;
    wire N__19722;
    wire N__19721;
    wire N__19718;
    wire N__19713;
    wire N__19708;
    wire N__19703;
    wire N__19696;
    wire N__19685;
    wire N__19682;
    wire N__19679;
    wire N__19676;
    wire N__19673;
    wire N__19672;
    wire N__19671;
    wire N__19668;
    wire N__19667;
    wire N__19666;
    wire N__19665;
    wire N__19660;
    wire N__19657;
    wire N__19656;
    wire N__19655;
    wire N__19652;
    wire N__19649;
    wire N__19646;
    wire N__19643;
    wire N__19640;
    wire N__19637;
    wire N__19634;
    wire N__19631;
    wire N__19616;
    wire N__19615;
    wire N__19614;
    wire N__19613;
    wire N__19610;
    wire N__19607;
    wire N__19604;
    wire N__19603;
    wire N__19598;
    wire N__19595;
    wire N__19592;
    wire N__19589;
    wire N__19588;
    wire N__19587;
    wire N__19584;
    wire N__19581;
    wire N__19576;
    wire N__19573;
    wire N__19570;
    wire N__19563;
    wire N__19556;
    wire N__19553;
    wire N__19550;
    wire N__19549;
    wire N__19548;
    wire N__19541;
    wire N__19538;
    wire N__19537;
    wire N__19536;
    wire N__19533;
    wire N__19530;
    wire N__19523;
    wire N__19520;
    wire N__19519;
    wire N__19518;
    wire N__19517;
    wire N__19516;
    wire N__19515;
    wire N__19514;
    wire N__19511;
    wire N__19508;
    wire N__19505;
    wire N__19504;
    wire N__19501;
    wire N__19498;
    wire N__19495;
    wire N__19492;
    wire N__19489;
    wire N__19486;
    wire N__19483;
    wire N__19478;
    wire N__19473;
    wire N__19472;
    wire N__19469;
    wire N__19468;
    wire N__19467;
    wire N__19466;
    wire N__19463;
    wire N__19460;
    wire N__19455;
    wire N__19452;
    wire N__19449;
    wire N__19446;
    wire N__19439;
    wire N__19432;
    wire N__19429;
    wire N__19418;
    wire N__19417;
    wire N__19416;
    wire N__19415;
    wire N__19412;
    wire N__19411;
    wire N__19408;
    wire N__19405;
    wire N__19402;
    wire N__19399;
    wire N__19396;
    wire N__19385;
    wire N__19382;
    wire N__19379;
    wire N__19376;
    wire N__19373;
    wire N__19372;
    wire N__19369;
    wire N__19366;
    wire N__19363;
    wire N__19362;
    wire N__19361;
    wire N__19358;
    wire N__19357;
    wire N__19354;
    wire N__19351;
    wire N__19348;
    wire N__19345;
    wire N__19342;
    wire N__19331;
    wire N__19328;
    wire N__19325;
    wire N__19322;
    wire N__19321;
    wire N__19320;
    wire N__19319;
    wire N__19316;
    wire N__19315;
    wire N__19312;
    wire N__19309;
    wire N__19306;
    wire N__19303;
    wire N__19302;
    wire N__19301;
    wire N__19296;
    wire N__19293;
    wire N__19290;
    wire N__19287;
    wire N__19282;
    wire N__19277;
    wire N__19274;
    wire N__19265;
    wire N__19264;
    wire N__19261;
    wire N__19260;
    wire N__19257;
    wire N__19256;
    wire N__19255;
    wire N__19252;
    wire N__19249;
    wire N__19246;
    wire N__19243;
    wire N__19240;
    wire N__19237;
    wire N__19234;
    wire N__19229;
    wire N__19220;
    wire N__19217;
    wire N__19214;
    wire N__19213;
    wire N__19212;
    wire N__19209;
    wire N__19206;
    wire N__19205;
    wire N__19202;
    wire N__19201;
    wire N__19200;
    wire N__19199;
    wire N__19198;
    wire N__19195;
    wire N__19192;
    wire N__19189;
    wire N__19186;
    wire N__19181;
    wire N__19176;
    wire N__19169;
    wire N__19160;
    wire N__19159;
    wire N__19156;
    wire N__19153;
    wire N__19150;
    wire N__19149;
    wire N__19146;
    wire N__19143;
    wire N__19140;
    wire N__19137;
    wire N__19130;
    wire N__19127;
    wire N__19126;
    wire N__19123;
    wire N__19120;
    wire N__19119;
    wire N__19116;
    wire N__19113;
    wire N__19112;
    wire N__19109;
    wire N__19106;
    wire N__19103;
    wire N__19098;
    wire N__19091;
    wire N__19088;
    wire N__19085;
    wire N__19082;
    wire N__19081;
    wire N__19080;
    wire N__19077;
    wire N__19076;
    wire N__19075;
    wire N__19072;
    wire N__19071;
    wire N__19070;
    wire N__19067;
    wire N__19066;
    wire N__19063;
    wire N__19062;
    wire N__19059;
    wire N__19056;
    wire N__19053;
    wire N__19052;
    wire N__19049;
    wire N__19048;
    wire N__19045;
    wire N__19042;
    wire N__19039;
    wire N__19036;
    wire N__19033;
    wire N__19026;
    wire N__19023;
    wire N__19020;
    wire N__19017;
    wire N__18998;
    wire N__18997;
    wire N__18994;
    wire N__18991;
    wire N__18990;
    wire N__18987;
    wire N__18986;
    wire N__18985;
    wire N__18984;
    wire N__18983;
    wire N__18982;
    wire N__18981;
    wire N__18978;
    wire N__18975;
    wire N__18972;
    wire N__18969;
    wire N__18962;
    wire N__18957;
    wire N__18952;
    wire N__18941;
    wire N__18940;
    wire N__18939;
    wire N__18938;
    wire N__18937;
    wire N__18934;
    wire N__18933;
    wire N__18932;
    wire N__18931;
    wire N__18928;
    wire N__18927;
    wire N__18924;
    wire N__18923;
    wire N__18922;
    wire N__18919;
    wire N__18918;
    wire N__18917;
    wire N__18916;
    wire N__18915;
    wire N__18914;
    wire N__18911;
    wire N__18908;
    wire N__18905;
    wire N__18900;
    wire N__18897;
    wire N__18892;
    wire N__18887;
    wire N__18884;
    wire N__18881;
    wire N__18876;
    wire N__18873;
    wire N__18870;
    wire N__18867;
    wire N__18864;
    wire N__18863;
    wire N__18860;
    wire N__18857;
    wire N__18854;
    wire N__18849;
    wire N__18842;
    wire N__18841;
    wire N__18836;
    wire N__18831;
    wire N__18828;
    wire N__18825;
    wire N__18822;
    wire N__18817;
    wire N__18814;
    wire N__18811;
    wire N__18808;
    wire N__18803;
    wire N__18800;
    wire N__18787;
    wire N__18782;
    wire N__18779;
    wire N__18776;
    wire N__18775;
    wire N__18774;
    wire N__18773;
    wire N__18772;
    wire N__18771;
    wire N__18770;
    wire N__18769;
    wire N__18768;
    wire N__18767;
    wire N__18766;
    wire N__18765;
    wire N__18764;
    wire N__18763;
    wire N__18762;
    wire N__18759;
    wire N__18756;
    wire N__18753;
    wire N__18750;
    wire N__18749;
    wire N__18746;
    wire N__18745;
    wire N__18742;
    wire N__18735;
    wire N__18730;
    wire N__18727;
    wire N__18724;
    wire N__18719;
    wire N__18716;
    wire N__18713;
    wire N__18710;
    wire N__18709;
    wire N__18708;
    wire N__18707;
    wire N__18704;
    wire N__18703;
    wire N__18700;
    wire N__18699;
    wire N__18696;
    wire N__18693;
    wire N__18686;
    wire N__18683;
    wire N__18678;
    wire N__18675;
    wire N__18670;
    wire N__18667;
    wire N__18662;
    wire N__18659;
    wire N__18656;
    wire N__18653;
    wire N__18650;
    wire N__18639;
    wire N__18620;
    wire N__18617;
    wire N__18614;
    wire N__18613;
    wire N__18610;
    wire N__18607;
    wire N__18606;
    wire N__18605;
    wire N__18604;
    wire N__18603;
    wire N__18602;
    wire N__18601;
    wire N__18596;
    wire N__18593;
    wire N__18590;
    wire N__18587;
    wire N__18584;
    wire N__18581;
    wire N__18578;
    wire N__18575;
    wire N__18568;
    wire N__18561;
    wire N__18558;
    wire N__18553;
    wire N__18552;
    wire N__18547;
    wire N__18544;
    wire N__18539;
    wire N__18536;
    wire N__18533;
    wire N__18530;
    wire N__18529;
    wire N__18528;
    wire N__18527;
    wire N__18520;
    wire N__18517;
    wire N__18512;
    wire N__18509;
    wire N__18506;
    wire N__18503;
    wire N__18500;
    wire N__18497;
    wire N__18494;
    wire N__18491;
    wire N__18488;
    wire N__18485;
    wire N__18482;
    wire N__18479;
    wire N__18476;
    wire N__18473;
    wire N__18470;
    wire N__18467;
    wire N__18464;
    wire N__18461;
    wire N__18458;
    wire N__18455;
    wire N__18452;
    wire N__18449;
    wire N__18448;
    wire N__18445;
    wire N__18442;
    wire N__18437;
    wire N__18434;
    wire N__18431;
    wire N__18428;
    wire N__18425;
    wire N__18422;
    wire N__18419;
    wire N__18416;
    wire N__18413;
    wire N__18410;
    wire N__18407;
    wire N__18404;
    wire N__18401;
    wire N__18398;
    wire N__18395;
    wire N__18394;
    wire N__18393;
    wire N__18392;
    wire N__18391;
    wire N__18390;
    wire N__18389;
    wire N__18386;
    wire N__18383;
    wire N__18382;
    wire N__18381;
    wire N__18378;
    wire N__18375;
    wire N__18372;
    wire N__18367;
    wire N__18364;
    wire N__18361;
    wire N__18356;
    wire N__18353;
    wire N__18338;
    wire N__18337;
    wire N__18336;
    wire N__18333;
    wire N__18332;
    wire N__18331;
    wire N__18330;
    wire N__18327;
    wire N__18324;
    wire N__18321;
    wire N__18316;
    wire N__18313;
    wire N__18302;
    wire N__18299;
    wire N__18296;
    wire N__18293;
    wire N__18290;
    wire N__18287;
    wire N__18284;
    wire N__18281;
    wire N__18278;
    wire N__18275;
    wire N__18272;
    wire N__18269;
    wire N__18266;
    wire N__18263;
    wire N__18260;
    wire N__18259;
    wire N__18256;
    wire N__18255;
    wire N__18252;
    wire N__18251;
    wire N__18248;
    wire N__18245;
    wire N__18240;
    wire N__18239;
    wire N__18236;
    wire N__18231;
    wire N__18228;
    wire N__18227;
    wire N__18226;
    wire N__18225;
    wire N__18224;
    wire N__18221;
    wire N__18218;
    wire N__18215;
    wire N__18210;
    wire N__18205;
    wire N__18194;
    wire N__18193;
    wire N__18192;
    wire N__18191;
    wire N__18188;
    wire N__18187;
    wire N__18186;
    wire N__18185;
    wire N__18184;
    wire N__18179;
    wire N__18176;
    wire N__18169;
    wire N__18166;
    wire N__18165;
    wire N__18164;
    wire N__18163;
    wire N__18160;
    wire N__18153;
    wire N__18150;
    wire N__18147;
    wire N__18142;
    wire N__18139;
    wire N__18136;
    wire N__18125;
    wire N__18124;
    wire N__18123;
    wire N__18120;
    wire N__18119;
    wire N__18114;
    wire N__18111;
    wire N__18108;
    wire N__18105;
    wire N__18104;
    wire N__18103;
    wire N__18102;
    wire N__18099;
    wire N__18094;
    wire N__18091;
    wire N__18090;
    wire N__18089;
    wire N__18088;
    wire N__18083;
    wire N__18080;
    wire N__18075;
    wire N__18070;
    wire N__18067;
    wire N__18056;
    wire N__18053;
    wire N__18050;
    wire N__18047;
    wire N__18044;
    wire N__18041;
    wire N__18038;
    wire N__18035;
    wire N__18032;
    wire N__18029;
    wire N__18028;
    wire N__18027;
    wire N__18026;
    wire N__18023;
    wire N__18020;
    wire N__18019;
    wire N__18018;
    wire N__18013;
    wire N__18008;
    wire N__18007;
    wire N__18006;
    wire N__18005;
    wire N__18004;
    wire N__18003;
    wire N__18002;
    wire N__17999;
    wire N__17996;
    wire N__17991;
    wire N__17984;
    wire N__17975;
    wire N__17974;
    wire N__17973;
    wire N__17970;
    wire N__17963;
    wire N__17962;
    wire N__17959;
    wire N__17958;
    wire N__17955;
    wire N__17952;
    wire N__17949;
    wire N__17946;
    wire N__17939;
    wire N__17930;
    wire N__17927;
    wire N__17924;
    wire N__17921;
    wire N__17918;
    wire N__17915;
    wire N__17912;
    wire N__17909;
    wire N__17906;
    wire N__17903;
    wire N__17900;
    wire N__17897;
    wire N__17894;
    wire N__17891;
    wire N__17888;
    wire N__17885;
    wire N__17882;
    wire N__17879;
    wire N__17876;
    wire N__17875;
    wire N__17874;
    wire N__17873;
    wire N__17872;
    wire N__17871;
    wire N__17870;
    wire N__17869;
    wire N__17868;
    wire N__17865;
    wire N__17858;
    wire N__17853;
    wire N__17848;
    wire N__17845;
    wire N__17834;
    wire N__17831;
    wire N__17828;
    wire N__17825;
    wire N__17824;
    wire N__17823;
    wire N__17820;
    wire N__17815;
    wire N__17810;
    wire N__17807;
    wire N__17804;
    wire N__17801;
    wire N__17798;
    wire N__17795;
    wire N__17794;
    wire N__17793;
    wire N__17792;
    wire N__17791;
    wire N__17790;
    wire N__17787;
    wire N__17786;
    wire N__17783;
    wire N__17782;
    wire N__17781;
    wire N__17780;
    wire N__17777;
    wire N__17774;
    wire N__17773;
    wire N__17770;
    wire N__17769;
    wire N__17768;
    wire N__17765;
    wire N__17764;
    wire N__17761;
    wire N__17756;
    wire N__17753;
    wire N__17742;
    wire N__17737;
    wire N__17730;
    wire N__17717;
    wire N__17716;
    wire N__17715;
    wire N__17714;
    wire N__17707;
    wire N__17704;
    wire N__17703;
    wire N__17702;
    wire N__17701;
    wire N__17700;
    wire N__17699;
    wire N__17698;
    wire N__17693;
    wire N__17692;
    wire N__17687;
    wire N__17684;
    wire N__17683;
    wire N__17680;
    wire N__17679;
    wire N__17676;
    wire N__17673;
    wire N__17670;
    wire N__17669;
    wire N__17668;
    wire N__17667;
    wire N__17666;
    wire N__17663;
    wire N__17660;
    wire N__17657;
    wire N__17654;
    wire N__17651;
    wire N__17648;
    wire N__17645;
    wire N__17640;
    wire N__17639;
    wire N__17636;
    wire N__17633;
    wire N__17628;
    wire N__17625;
    wire N__17622;
    wire N__17613;
    wire N__17608;
    wire N__17605;
    wire N__17588;
    wire N__17585;
    wire N__17582;
    wire N__17579;
    wire N__17576;
    wire N__17573;
    wire N__17572;
    wire N__17569;
    wire N__17566;
    wire N__17563;
    wire N__17560;
    wire N__17557;
    wire N__17552;
    wire N__17549;
    wire N__17546;
    wire N__17543;
    wire N__17540;
    wire N__17537;
    wire N__17536;
    wire N__17535;
    wire N__17534;
    wire N__17527;
    wire N__17526;
    wire N__17525;
    wire N__17522;
    wire N__17519;
    wire N__17514;
    wire N__17507;
    wire N__17506;
    wire N__17503;
    wire N__17500;
    wire N__17495;
    wire N__17492;
    wire N__17489;
    wire N__17486;
    wire N__17483;
    wire N__17482;
    wire N__17479;
    wire N__17476;
    wire N__17471;
    wire N__17468;
    wire N__17467;
    wire N__17464;
    wire N__17461;
    wire N__17458;
    wire N__17455;
    wire N__17452;
    wire N__17449;
    wire N__17444;
    wire N__17441;
    wire N__17438;
    wire N__17435;
    wire N__17432;
    wire N__17429;
    wire N__17426;
    wire N__17423;
    wire N__17420;
    wire N__17417;
    wire N__17414;
    wire N__17411;
    wire N__17410;
    wire N__17409;
    wire N__17404;
    wire N__17401;
    wire N__17400;
    wire N__17399;
    wire N__17398;
    wire N__17395;
    wire N__17392;
    wire N__17391;
    wire N__17390;
    wire N__17387;
    wire N__17384;
    wire N__17381;
    wire N__17380;
    wire N__17377;
    wire N__17374;
    wire N__17371;
    wire N__17368;
    wire N__17363;
    wire N__17360;
    wire N__17357;
    wire N__17342;
    wire N__17341;
    wire N__17338;
    wire N__17335;
    wire N__17332;
    wire N__17327;
    wire N__17324;
    wire N__17321;
    wire N__17318;
    wire N__17315;
    wire N__17312;
    wire N__17309;
    wire N__17306;
    wire N__17303;
    wire N__17300;
    wire N__17297;
    wire N__17294;
    wire N__17291;
    wire N__17288;
    wire N__17285;
    wire N__17282;
    wire N__17279;
    wire N__17276;
    wire N__17273;
    wire N__17270;
    wire N__17267;
    wire N__17264;
    wire N__17261;
    wire N__17258;
    wire N__17255;
    wire N__17252;
    wire N__17249;
    wire N__17246;
    wire N__17243;
    wire N__17240;
    wire N__17237;
    wire N__17234;
    wire N__17231;
    wire N__17228;
    wire N__17225;
    wire N__17222;
    wire N__17219;
    wire N__17216;
    wire N__17213;
    wire N__17210;
    wire N__17207;
    wire N__17204;
    wire N__17201;
    wire N__17198;
    wire N__17195;
    wire N__17192;
    wire N__17189;
    wire N__17186;
    wire N__17183;
    wire N__17180;
    wire N__17177;
    wire N__17176;
    wire N__17175;
    wire N__17174;
    wire N__17173;
    wire N__17172;
    wire N__17171;
    wire N__17170;
    wire N__17167;
    wire N__17154;
    wire N__17151;
    wire N__17148;
    wire N__17145;
    wire N__17142;
    wire N__17139;
    wire N__17136;
    wire N__17133;
    wire N__17126;
    wire N__17123;
    wire N__17120;
    wire N__17117;
    wire N__17116;
    wire N__17115;
    wire N__17114;
    wire N__17113;
    wire N__17112;
    wire N__17109;
    wire N__17108;
    wire N__17105;
    wire N__17102;
    wire N__17099;
    wire N__17094;
    wire N__17089;
    wire N__17088;
    wire N__17087;
    wire N__17084;
    wire N__17081;
    wire N__17074;
    wire N__17069;
    wire N__17060;
    wire N__17057;
    wire N__17054;
    wire N__17051;
    wire N__17048;
    wire N__17045;
    wire N__17042;
    wire N__17039;
    wire N__17036;
    wire N__17033;
    wire N__17032;
    wire N__17031;
    wire N__17030;
    wire N__17021;
    wire N__17020;
    wire N__17019;
    wire N__17018;
    wire N__17017;
    wire N__17014;
    wire N__17013;
    wire N__17012;
    wire N__17011;
    wire N__17004;
    wire N__17001;
    wire N__17000;
    wire N__16997;
    wire N__16994;
    wire N__16991;
    wire N__16988;
    wire N__16985;
    wire N__16982;
    wire N__16979;
    wire N__16976;
    wire N__16969;
    wire N__16958;
    wire N__16957;
    wire N__16954;
    wire N__16953;
    wire N__16952;
    wire N__16951;
    wire N__16950;
    wire N__16947;
    wire N__16946;
    wire N__16943;
    wire N__16940;
    wire N__16937;
    wire N__16936;
    wire N__16935;
    wire N__16930;
    wire N__16927;
    wire N__16924;
    wire N__16921;
    wire N__16916;
    wire N__16911;
    wire N__16906;
    wire N__16895;
    wire N__16892;
    wire N__16889;
    wire N__16886;
    wire N__16883;
    wire N__16880;
    wire N__16877;
    wire N__16874;
    wire N__16871;
    wire N__16868;
    wire N__16865;
    wire N__16862;
    wire N__16859;
    wire N__16856;
    wire N__16855;
    wire N__16852;
    wire N__16849;
    wire N__16844;
    wire N__16841;
    wire N__16838;
    wire N__16835;
    wire N__16832;
    wire N__16829;
    wire N__16826;
    wire N__16823;
    wire N__16820;
    wire N__16817;
    wire N__16814;
    wire N__16811;
    wire N__16808;
    wire N__16805;
    wire N__16804;
    wire N__16803;
    wire N__16800;
    wire N__16797;
    wire N__16794;
    wire N__16787;
    wire N__16784;
    wire N__16781;
    wire N__16778;
    wire N__16775;
    wire N__16772;
    wire N__16769;
    wire N__16766;
    wire N__16763;
    wire N__16760;
    wire N__16757;
    wire N__16754;
    wire N__16751;
    wire N__16748;
    wire N__16745;
    wire N__16742;
    wire N__16739;
    wire N__16736;
    wire N__16733;
    wire N__16732;
    wire N__16729;
    wire N__16726;
    wire N__16725;
    wire N__16724;
    wire N__16723;
    wire N__16722;
    wire N__16719;
    wire N__16716;
    wire N__16713;
    wire N__16706;
    wire N__16697;
    wire N__16694;
    wire N__16691;
    wire N__16688;
    wire N__16685;
    wire N__16682;
    wire N__16679;
    wire N__16678;
    wire N__16677;
    wire N__16674;
    wire N__16673;
    wire N__16670;
    wire N__16667;
    wire N__16664;
    wire N__16661;
    wire N__16656;
    wire N__16651;
    wire N__16648;
    wire N__16645;
    wire N__16642;
    wire N__16639;
    wire N__16634;
    wire N__16633;
    wire N__16628;
    wire N__16625;
    wire N__16622;
    wire N__16619;
    wire N__16616;
    wire N__16613;
    wire N__16610;
    wire N__16607;
    wire N__16604;
    wire N__16601;
    wire N__16598;
    wire N__16595;
    wire N__16592;
    wire N__16589;
    wire N__16586;
    wire N__16583;
    wire N__16580;
    wire N__16577;
    wire N__16574;
    wire N__16571;
    wire N__16568;
    wire N__16565;
    wire N__16562;
    wire N__16559;
    wire N__16556;
    wire N__16553;
    wire N__16550;
    wire N__16547;
    wire N__16544;
    wire N__16541;
    wire N__16538;
    wire N__16535;
    wire N__16532;
    wire N__16529;
    wire N__16526;
    wire N__16523;
    wire N__16520;
    wire N__16517;
    wire N__16514;
    wire N__16511;
    wire N__16508;
    wire N__16505;
    wire N__16502;
    wire N__16499;
    wire N__16496;
    wire N__16493;
    wire N__16490;
    wire N__16487;
    wire N__16484;
    wire N__16481;
    wire N__16480;
    wire N__16479;
    wire N__16478;
    wire N__16475;
    wire N__16474;
    wire N__16473;
    wire N__16470;
    wire N__16467;
    wire N__16466;
    wire N__16465;
    wire N__16462;
    wire N__16459;
    wire N__16458;
    wire N__16455;
    wire N__16452;
    wire N__16445;
    wire N__16442;
    wire N__16437;
    wire N__16434;
    wire N__16431;
    wire N__16418;
    wire N__16415;
    wire N__16412;
    wire N__16409;
    wire N__16406;
    wire N__16405;
    wire N__16402;
    wire N__16401;
    wire N__16400;
    wire N__16397;
    wire N__16396;
    wire N__16395;
    wire N__16394;
    wire N__16391;
    wire N__16388;
    wire N__16381;
    wire N__16378;
    wire N__16375;
    wire N__16374;
    wire N__16371;
    wire N__16368;
    wire N__16361;
    wire N__16358;
    wire N__16349;
    wire N__16346;
    wire N__16343;
    wire N__16340;
    wire N__16337;
    wire N__16334;
    wire N__16331;
    wire N__16330;
    wire N__16327;
    wire N__16324;
    wire N__16321;
    wire N__16318;
    wire N__16315;
    wire N__16312;
    wire N__16309;
    wire N__16304;
    wire N__16301;
    wire N__16298;
    wire N__16295;
    wire N__16292;
    wire N__16289;
    wire N__16286;
    wire N__16283;
    wire N__16280;
    wire N__16277;
    wire N__16274;
    wire N__16271;
    wire N__16270;
    wire N__16267;
    wire N__16264;
    wire N__16259;
    wire N__16256;
    wire N__16253;
    wire N__16250;
    wire N__16247;
    wire N__16244;
    wire N__16241;
    wire N__16238;
    wire N__16235;
    wire N__16232;
    wire N__16229;
    wire N__16228;
    wire N__16225;
    wire N__16224;
    wire N__16223;
    wire N__16222;
    wire N__16221;
    wire N__16218;
    wire N__16217;
    wire N__16214;
    wire N__16211;
    wire N__16206;
    wire N__16203;
    wire N__16202;
    wire N__16199;
    wire N__16196;
    wire N__16187;
    wire N__16184;
    wire N__16175;
    wire N__16174;
    wire N__16173;
    wire N__16172;
    wire N__16171;
    wire N__16170;
    wire N__16169;
    wire N__16168;
    wire N__16165;
    wire N__16162;
    wire N__16159;
    wire N__16152;
    wire N__16151;
    wire N__16150;
    wire N__16147;
    wire N__16144;
    wire N__16141;
    wire N__16138;
    wire N__16133;
    wire N__16128;
    wire N__16115;
    wire N__16114;
    wire N__16113;
    wire N__16112;
    wire N__16111;
    wire N__16108;
    wire N__16105;
    wire N__16102;
    wire N__16101;
    wire N__16100;
    wire N__16097;
    wire N__16094;
    wire N__16091;
    wire N__16088;
    wire N__16085;
    wire N__16078;
    wire N__16077;
    wire N__16076;
    wire N__16069;
    wire N__16064;
    wire N__16059;
    wire N__16056;
    wire N__16051;
    wire N__16046;
    wire N__16045;
    wire N__16044;
    wire N__16041;
    wire N__16038;
    wire N__16037;
    wire N__16034;
    wire N__16031;
    wire N__16028;
    wire N__16025;
    wire N__16024;
    wire N__16023;
    wire N__16020;
    wire N__16017;
    wire N__16014;
    wire N__16011;
    wire N__16008;
    wire N__16005;
    wire N__15992;
    wire N__15989;
    wire N__15986;
    wire N__15983;
    wire N__15980;
    wire N__15977;
    wire N__15974;
    wire N__15971;
    wire N__15968;
    wire N__15965;
    wire N__15962;
    wire N__15959;
    wire N__15956;
    wire N__15953;
    wire N__15950;
    wire N__15947;
    wire N__15946;
    wire N__15945;
    wire N__15942;
    wire N__15937;
    wire N__15934;
    wire N__15931;
    wire N__15926;
    wire N__15923;
    wire N__15920;
    wire N__15917;
    wire N__15914;
    wire N__15911;
    wire N__15910;
    wire N__15907;
    wire N__15904;
    wire N__15903;
    wire N__15902;
    wire N__15901;
    wire N__15896;
    wire N__15893;
    wire N__15890;
    wire N__15887;
    wire N__15884;
    wire N__15879;
    wire N__15872;
    wire N__15871;
    wire N__15868;
    wire N__15867;
    wire N__15866;
    wire N__15865;
    wire N__15862;
    wire N__15859;
    wire N__15854;
    wire N__15851;
    wire N__15848;
    wire N__15847;
    wire N__15846;
    wire N__15845;
    wire N__15844;
    wire N__15841;
    wire N__15838;
    wire N__15835;
    wire N__15832;
    wire N__15829;
    wire N__15822;
    wire N__15809;
    wire N__15806;
    wire N__15803;
    wire N__15800;
    wire N__15797;
    wire N__15794;
    wire N__15791;
    wire N__15788;
    wire N__15787;
    wire N__15782;
    wire N__15779;
    wire N__15776;
    wire N__15775;
    wire N__15770;
    wire N__15767;
    wire N__15764;
    wire N__15761;
    wire N__15758;
    wire N__15755;
    wire N__15752;
    wire N__15749;
    wire N__15746;
    wire N__15743;
    wire N__15742;
    wire N__15739;
    wire N__15736;
    wire N__15731;
    wire N__15728;
    wire N__15725;
    wire N__15722;
    wire N__15721;
    wire N__15720;
    wire N__15719;
    wire N__15716;
    wire N__15711;
    wire N__15708;
    wire N__15705;
    wire N__15702;
    wire N__15699;
    wire N__15696;
    wire N__15693;
    wire N__15686;
    wire N__15685;
    wire N__15684;
    wire N__15683;
    wire N__15682;
    wire N__15681;
    wire N__15680;
    wire N__15679;
    wire N__15678;
    wire N__15677;
    wire N__15674;
    wire N__15671;
    wire N__15668;
    wire N__15665;
    wire N__15660;
    wire N__15655;
    wire N__15652;
    wire N__15645;
    wire N__15642;
    wire N__15639;
    wire N__15634;
    wire N__15633;
    wire N__15632;
    wire N__15629;
    wire N__15626;
    wire N__15621;
    wire N__15618;
    wire N__15613;
    wire N__15608;
    wire N__15599;
    wire N__15598;
    wire N__15597;
    wire N__15596;
    wire N__15595;
    wire N__15594;
    wire N__15581;
    wire N__15578;
    wire N__15577;
    wire N__15576;
    wire N__15575;
    wire N__15572;
    wire N__15567;
    wire N__15566;
    wire N__15565;
    wire N__15564;
    wire N__15563;
    wire N__15560;
    wire N__15559;
    wire N__15554;
    wire N__15541;
    wire N__15536;
    wire N__15535;
    wire N__15534;
    wire N__15531;
    wire N__15526;
    wire N__15521;
    wire N__15518;
    wire N__15515;
    wire N__15512;
    wire N__15509;
    wire N__15506;
    wire N__15503;
    wire N__15500;
    wire N__15497;
    wire N__15494;
    wire N__15491;
    wire N__15490;
    wire N__15487;
    wire N__15484;
    wire N__15481;
    wire N__15478;
    wire N__15477;
    wire N__15474;
    wire N__15471;
    wire N__15470;
    wire N__15469;
    wire N__15466;
    wire N__15463;
    wire N__15460;
    wire N__15457;
    wire N__15454;
    wire N__15451;
    wire N__15440;
    wire N__15439;
    wire N__15434;
    wire N__15431;
    wire N__15428;
    wire N__15425;
    wire N__15422;
    wire N__15419;
    wire N__15416;
    wire N__15413;
    wire N__15412;
    wire N__15409;
    wire N__15406;
    wire N__15403;
    wire N__15400;
    wire N__15395;
    wire N__15392;
    wire N__15389;
    wire N__15386;
    wire N__15383;
    wire N__15380;
    wire N__15377;
    wire N__15376;
    wire N__15375;
    wire N__15374;
    wire N__15373;
    wire N__15372;
    wire N__15371;
    wire N__15370;
    wire N__15369;
    wire N__15366;
    wire N__15363;
    wire N__15360;
    wire N__15357;
    wire N__15350;
    wire N__15345;
    wire N__15332;
    wire N__15329;
    wire N__15326;
    wire N__15325;
    wire N__15324;
    wire N__15321;
    wire N__15318;
    wire N__15317;
    wire N__15316;
    wire N__15315;
    wire N__15312;
    wire N__15301;
    wire N__15296;
    wire N__15293;
    wire N__15290;
    wire N__15287;
    wire N__15284;
    wire N__15281;
    wire N__15278;
    wire N__15275;
    wire N__15274;
    wire N__15271;
    wire N__15268;
    wire N__15263;
    wire N__15260;
    wire N__15257;
    wire N__15254;
    wire N__15251;
    wire N__15248;
    wire N__15245;
    wire N__15242;
    wire N__15239;
    wire N__15236;
    wire N__15235;
    wire N__15234;
    wire N__15231;
    wire N__15228;
    wire N__15225;
    wire N__15224;
    wire N__15219;
    wire N__15216;
    wire N__15215;
    wire N__15214;
    wire N__15213;
    wire N__15210;
    wire N__15207;
    wire N__15204;
    wire N__15197;
    wire N__15194;
    wire N__15185;
    wire N__15184;
    wire N__15183;
    wire N__15182;
    wire N__15181;
    wire N__15180;
    wire N__15177;
    wire N__15174;
    wire N__15165;
    wire N__15162;
    wire N__15157;
    wire N__15154;
    wire N__15151;
    wire N__15146;
    wire N__15145;
    wire N__15140;
    wire N__15139;
    wire N__15138;
    wire N__15135;
    wire N__15132;
    wire N__15129;
    wire N__15126;
    wire N__15119;
    wire N__15116;
    wire N__15113;
    wire N__15110;
    wire N__15107;
    wire N__15104;
    wire N__15103;
    wire N__15100;
    wire N__15097;
    wire N__15094;
    wire N__15091;
    wire N__15086;
    wire N__15083;
    wire N__15080;
    wire N__15077;
    wire N__15074;
    wire N__15073;
    wire N__15070;
    wire N__15067;
    wire N__15062;
    wire N__15061;
    wire N__15060;
    wire N__15059;
    wire N__15058;
    wire N__15055;
    wire N__15054;
    wire N__15053;
    wire N__15046;
    wire N__15043;
    wire N__15036;
    wire N__15029;
    wire N__15028;
    wire N__15027;
    wire N__15026;
    wire N__15023;
    wire N__15022;
    wire N__15021;
    wire N__15020;
    wire N__15017;
    wire N__15008;
    wire N__15003;
    wire N__14998;
    wire N__14993;
    wire N__14990;
    wire N__14989;
    wire N__14988;
    wire N__14987;
    wire N__14986;
    wire N__14985;
    wire N__14984;
    wire N__14981;
    wire N__14978;
    wire N__14975;
    wire N__14966;
    wire N__14957;
    wire N__14956;
    wire N__14955;
    wire N__14954;
    wire N__14953;
    wire N__14952;
    wire N__14949;
    wire N__14942;
    wire N__14939;
    wire N__14936;
    wire N__14927;
    wire N__14926;
    wire N__14925;
    wire N__14924;
    wire N__14919;
    wire N__14916;
    wire N__14913;
    wire N__14906;
    wire N__14905;
    wire N__14902;
    wire N__14899;
    wire N__14898;
    wire N__14897;
    wire N__14892;
    wire N__14889;
    wire N__14886;
    wire N__14883;
    wire N__14880;
    wire N__14873;
    wire N__14872;
    wire N__14869;
    wire N__14866;
    wire N__14863;
    wire N__14860;
    wire N__14859;
    wire N__14858;
    wire N__14857;
    wire N__14856;
    wire N__14853;
    wire N__14850;
    wire N__14847;
    wire N__14844;
    wire N__14839;
    wire N__14834;
    wire N__14825;
    wire N__14824;
    wire N__14821;
    wire N__14820;
    wire N__14817;
    wire N__14814;
    wire N__14811;
    wire N__14808;
    wire N__14801;
    wire N__14798;
    wire N__14797;
    wire N__14796;
    wire N__14795;
    wire N__14794;
    wire N__14793;
    wire N__14792;
    wire N__14791;
    wire N__14788;
    wire N__14787;
    wire N__14786;
    wire N__14785;
    wire N__14782;
    wire N__14781;
    wire N__14778;
    wire N__14769;
    wire N__14766;
    wire N__14763;
    wire N__14756;
    wire N__14753;
    wire N__14750;
    wire N__14747;
    wire N__14744;
    wire N__14741;
    wire N__14736;
    wire N__14731;
    wire N__14728;
    wire N__14725;
    wire N__14718;
    wire N__14713;
    wire N__14710;
    wire N__14705;
    wire N__14704;
    wire N__14701;
    wire N__14698;
    wire N__14695;
    wire N__14694;
    wire N__14693;
    wire N__14690;
    wire N__14687;
    wire N__14684;
    wire N__14681;
    wire N__14678;
    wire N__14675;
    wire N__14670;
    wire N__14663;
    wire N__14660;
    wire N__14659;
    wire N__14658;
    wire N__14655;
    wire N__14652;
    wire N__14649;
    wire N__14648;
    wire N__14643;
    wire N__14640;
    wire N__14637;
    wire N__14634;
    wire N__14631;
    wire N__14624;
    wire N__14621;
    wire N__14618;
    wire N__14615;
    wire N__14612;
    wire N__14609;
    wire N__14606;
    wire N__14605;
    wire N__14602;
    wire N__14599;
    wire N__14594;
    wire N__14591;
    wire N__14588;
    wire N__14585;
    wire N__14584;
    wire N__14583;
    wire N__14576;
    wire N__14573;
    wire N__14570;
    wire N__14567;
    wire N__14564;
    wire N__14561;
    wire N__14558;
    wire N__14555;
    wire N__14552;
    wire N__14549;
    wire N__14546;
    wire N__14545;
    wire N__14542;
    wire N__14539;
    wire N__14536;
    wire N__14533;
    wire N__14530;
    wire N__14525;
    wire N__14522;
    wire N__14519;
    wire N__14516;
    wire N__14513;
    wire N__14510;
    wire N__14509;
    wire N__14506;
    wire N__14503;
    wire N__14498;
    wire N__14495;
    wire N__14492;
    wire N__14489;
    wire N__14486;
    wire N__14485;
    wire N__14482;
    wire N__14479;
    wire N__14476;
    wire N__14473;
    wire N__14470;
    wire N__14465;
    wire N__14462;
    wire N__14459;
    wire N__14456;
    wire N__14455;
    wire N__14452;
    wire N__14449;
    wire N__14446;
    wire N__14443;
    wire N__14440;
    wire N__14437;
    wire N__14434;
    wire N__14429;
    wire N__14426;
    wire N__14423;
    wire N__14420;
    wire N__14419;
    wire N__14418;
    wire N__14417;
    wire N__14416;
    wire N__14415;
    wire N__14414;
    wire N__14413;
    wire N__14410;
    wire N__14405;
    wire N__14394;
    wire N__14389;
    wire N__14386;
    wire N__14383;
    wire N__14380;
    wire N__14375;
    wire N__14372;
    wire N__14371;
    wire N__14368;
    wire N__14365;
    wire N__14362;
    wire N__14359;
    wire N__14356;
    wire N__14353;
    wire N__14348;
    wire N__14347;
    wire N__14346;
    wire N__14345;
    wire N__14344;
    wire N__14343;
    wire N__14342;
    wire N__14341;
    wire N__14340;
    wire N__14339;
    wire N__14328;
    wire N__14323;
    wire N__14322;
    wire N__14321;
    wire N__14314;
    wire N__14311;
    wire N__14308;
    wire N__14303;
    wire N__14300;
    wire N__14299;
    wire N__14298;
    wire N__14295;
    wire N__14292;
    wire N__14287;
    wire N__14282;
    wire N__14279;
    wire N__14270;
    wire N__14269;
    wire N__14266;
    wire N__14261;
    wire N__14258;
    wire N__14255;
    wire N__14254;
    wire N__14251;
    wire N__14248;
    wire N__14243;
    wire N__14242;
    wire N__14241;
    wire N__14238;
    wire N__14235;
    wire N__14232;
    wire N__14231;
    wire N__14228;
    wire N__14225;
    wire N__14222;
    wire N__14219;
    wire N__14216;
    wire N__14209;
    wire N__14204;
    wire N__14201;
    wire N__14200;
    wire N__14199;
    wire N__14198;
    wire N__14195;
    wire N__14192;
    wire N__14189;
    wire N__14186;
    wire N__14181;
    wire N__14178;
    wire N__14171;
    wire N__14168;
    wire N__14165;
    wire N__14162;
    wire N__14159;
    wire N__14156;
    wire N__14153;
    wire N__14150;
    wire N__14147;
    wire N__14144;
    wire N__14141;
    wire N__14138;
    wire N__14135;
    wire N__14132;
    wire N__14129;
    wire N__14126;
    wire N__14123;
    wire N__14120;
    wire N__14117;
    wire N__14114;
    wire N__14111;
    wire N__14108;
    wire N__14105;
    wire N__14102;
    wire N__14099;
    wire N__14096;
    wire N__14095;
    wire N__14094;
    wire N__14089;
    wire N__14086;
    wire N__14083;
    wire N__14078;
    wire N__14075;
    wire N__14072;
    wire N__14069;
    wire N__14066;
    wire N__14063;
    wire N__14060;
    wire N__14059;
    wire N__14056;
    wire N__14053;
    wire N__14050;
    wire N__14047;
    wire N__14044;
    wire N__14041;
    wire N__14038;
    wire N__14033;
    wire N__14030;
    wire N__14027;
    wire N__14026;
    wire N__14023;
    wire N__14020;
    wire N__14017;
    wire N__14014;
    wire N__14011;
    wire N__14006;
    wire N__14003;
    wire N__14000;
    wire N__13999;
    wire N__13996;
    wire N__13993;
    wire N__13990;
    wire N__13987;
    wire N__13984;
    wire N__13981;
    wire N__13978;
    wire N__13973;
    wire N__13970;
    wire N__13967;
    wire N__13964;
    wire N__13963;
    wire N__13962;
    wire N__13959;
    wire N__13954;
    wire N__13949;
    wire N__13946;
    wire N__13943;
    wire N__13940;
    wire N__13937;
    wire N__13936;
    wire N__13933;
    wire N__13930;
    wire N__13927;
    wire N__13924;
    wire N__13919;
    wire N__13916;
    wire N__13913;
    wire N__13912;
    wire N__13909;
    wire N__13906;
    wire N__13903;
    wire N__13900;
    wire N__13895;
    wire N__13894;
    wire N__13893;
    wire N__13892;
    wire N__13889;
    wire N__13886;
    wire N__13881;
    wire N__13874;
    wire N__13871;
    wire N__13868;
    wire N__13867;
    wire N__13864;
    wire N__13861;
    wire N__13858;
    wire N__13853;
    wire N__13852;
    wire N__13851;
    wire N__13848;
    wire N__13845;
    wire N__13842;
    wire N__13835;
    wire N__13832;
    wire N__13829;
    wire N__13828;
    wire N__13823;
    wire N__13820;
    wire N__13817;
    wire N__13816;
    wire N__13811;
    wire N__13808;
    wire N__13805;
    wire N__13804;
    wire N__13803;
    wire N__13802;
    wire N__13801;
    wire N__13800;
    wire N__13797;
    wire N__13796;
    wire N__13793;
    wire N__13790;
    wire N__13787;
    wire N__13778;
    wire N__13769;
    wire N__13766;
    wire N__13763;
    wire N__13760;
    wire N__13759;
    wire N__13758;
    wire N__13757;
    wire N__13754;
    wire N__13751;
    wire N__13746;
    wire N__13745;
    wire N__13744;
    wire N__13743;
    wire N__13742;
    wire N__13741;
    wire N__13734;
    wire N__13723;
    wire N__13718;
    wire N__13715;
    wire N__13712;
    wire N__13709;
    wire N__13706;
    wire N__13703;
    wire N__13700;
    wire N__13697;
    wire N__13694;
    wire N__13691;
    wire N__13688;
    wire N__13687;
    wire N__13686;
    wire N__13683;
    wire N__13680;
    wire N__13675;
    wire N__13670;
    wire N__13669;
    wire N__13668;
    wire N__13667;
    wire N__13666;
    wire N__13665;
    wire N__13662;
    wire N__13659;
    wire N__13650;
    wire N__13643;
    wire N__13642;
    wire N__13639;
    wire N__13638;
    wire N__13635;
    wire N__13632;
    wire N__13629;
    wire N__13626;
    wire N__13623;
    wire N__13620;
    wire N__13619;
    wire N__13612;
    wire N__13609;
    wire N__13604;
    wire N__13603;
    wire N__13602;
    wire N__13601;
    wire N__13598;
    wire N__13595;
    wire N__13592;
    wire N__13589;
    wire N__13586;
    wire N__13583;
    wire N__13578;
    wire N__13575;
    wire N__13568;
    wire N__13565;
    wire N__13562;
    wire N__13559;
    wire N__13556;
    wire N__13553;
    wire N__13552;
    wire N__13549;
    wire N__13546;
    wire N__13545;
    wire N__13542;
    wire N__13539;
    wire N__13536;
    wire N__13535;
    wire N__13532;
    wire N__13529;
    wire N__13526;
    wire N__13523;
    wire N__13514;
    wire N__13513;
    wire N__13510;
    wire N__13509;
    wire N__13508;
    wire N__13505;
    wire N__13502;
    wire N__13499;
    wire N__13496;
    wire N__13493;
    wire N__13488;
    wire N__13481;
    wire N__13480;
    wire N__13477;
    wire N__13474;
    wire N__13471;
    wire N__13468;
    wire N__13463;
    wire N__13460;
    wire N__13459;
    wire N__13456;
    wire N__13453;
    wire N__13450;
    wire N__13447;
    wire N__13444;
    wire N__13441;
    wire N__13436;
    wire N__13433;
    wire N__13430;
    wire N__13427;
    wire N__13424;
    wire N__13421;
    wire N__13418;
    wire N__13415;
    wire N__13412;
    wire N__13411;
    wire N__13408;
    wire N__13405;
    wire N__13402;
    wire N__13399;
    wire N__13394;
    wire N__13391;
    wire N__13388;
    wire N__13385;
    wire N__13382;
    wire N__13381;
    wire N__13380;
    wire N__13379;
    wire N__13376;
    wire N__13373;
    wire N__13370;
    wire N__13365;
    wire N__13358;
    wire N__13357;
    wire N__13356;
    wire N__13355;
    wire N__13352;
    wire N__13351;
    wire N__13350;
    wire N__13349;
    wire N__13348;
    wire N__13347;
    wire N__13344;
    wire N__13339;
    wire N__13336;
    wire N__13333;
    wire N__13330;
    wire N__13325;
    wire N__13322;
    wire N__13317;
    wire N__13304;
    wire N__13303;
    wire N__13302;
    wire N__13301;
    wire N__13300;
    wire N__13297;
    wire N__13294;
    wire N__13287;
    wire N__13280;
    wire N__13277;
    wire N__13274;
    wire N__13271;
    wire N__13268;
    wire N__13267;
    wire N__13266;
    wire N__13263;
    wire N__13260;
    wire N__13257;
    wire N__13254;
    wire N__13251;
    wire N__13248;
    wire N__13241;
    wire N__13238;
    wire N__13237;
    wire N__13234;
    wire N__13233;
    wire N__13232;
    wire N__13231;
    wire N__13230;
    wire N__13229;
    wire N__13228;
    wire N__13227;
    wire N__13224;
    wire N__13223;
    wire N__13220;
    wire N__13219;
    wire N__13218;
    wire N__13215;
    wire N__13210;
    wire N__13207;
    wire N__13204;
    wire N__13199;
    wire N__13196;
    wire N__13193;
    wire N__13190;
    wire N__13185;
    wire N__13180;
    wire N__13173;
    wire N__13170;
    wire N__13163;
    wire N__13158;
    wire N__13151;
    wire N__13148;
    wire N__13145;
    wire N__13142;
    wire N__13141;
    wire N__13138;
    wire N__13135;
    wire N__13130;
    wire N__13127;
    wire N__13124;
    wire N__13121;
    wire N__13118;
    wire N__13115;
    wire N__13112;
    wire N__13109;
    wire N__13106;
    wire N__13103;
    wire N__13102;
    wire N__13099;
    wire N__13096;
    wire N__13095;
    wire N__13092;
    wire N__13089;
    wire N__13086;
    wire N__13085;
    wire N__13080;
    wire N__13077;
    wire N__13074;
    wire N__13067;
    wire N__13064;
    wire N__13061;
    wire N__13060;
    wire N__13059;
    wire N__13058;
    wire N__13055;
    wire N__13052;
    wire N__13049;
    wire N__13046;
    wire N__13041;
    wire N__13038;
    wire N__13031;
    wire N__13028;
    wire N__13027;
    wire N__13024;
    wire N__13021;
    wire N__13020;
    wire N__13017;
    wire N__13014;
    wire N__13011;
    wire N__13010;
    wire N__13005;
    wire N__13002;
    wire N__12999;
    wire N__12992;
    wire N__12991;
    wire N__12988;
    wire N__12987;
    wire N__12986;
    wire N__12983;
    wire N__12980;
    wire N__12977;
    wire N__12974;
    wire N__12971;
    wire N__12966;
    wire N__12959;
    wire N__12958;
    wire N__12955;
    wire N__12952;
    wire N__12951;
    wire N__12948;
    wire N__12945;
    wire N__12942;
    wire N__12941;
    wire N__12936;
    wire N__12933;
    wire N__12930;
    wire N__12923;
    wire N__12920;
    wire N__12919;
    wire N__12916;
    wire N__12915;
    wire N__12914;
    wire N__12911;
    wire N__12908;
    wire N__12905;
    wire N__12902;
    wire N__12899;
    wire N__12894;
    wire N__12887;
    wire N__12886;
    wire N__12883;
    wire N__12880;
    wire N__12879;
    wire N__12876;
    wire N__12873;
    wire N__12870;
    wire N__12869;
    wire N__12864;
    wire N__12861;
    wire N__12858;
    wire N__12851;
    wire N__12848;
    wire N__12847;
    wire N__12846;
    wire N__12845;
    wire N__12842;
    wire N__12839;
    wire N__12836;
    wire N__12833;
    wire N__12830;
    wire N__12827;
    wire N__12824;
    wire N__12821;
    wire N__12812;
    wire N__12809;
    wire N__12808;
    wire N__12807;
    wire N__12804;
    wire N__12801;
    wire N__12798;
    wire N__12791;
    wire N__12788;
    wire N__12785;
    wire N__12784;
    wire N__12783;
    wire N__12780;
    wire N__12777;
    wire N__12774;
    wire N__12767;
    wire N__12764;
    wire N__12763;
    wire N__12762;
    wire N__12759;
    wire N__12756;
    wire N__12753;
    wire N__12750;
    wire N__12747;
    wire N__12744;
    wire N__12737;
    wire N__12736;
    wire N__12735;
    wire N__12732;
    wire N__12729;
    wire N__12726;
    wire N__12723;
    wire N__12720;
    wire N__12717;
    wire N__12714;
    wire N__12707;
    wire N__12704;
    wire N__12703;
    wire N__12702;
    wire N__12699;
    wire N__12696;
    wire N__12693;
    wire N__12690;
    wire N__12687;
    wire N__12684;
    wire N__12677;
    wire N__12676;
    wire N__12675;
    wire N__12672;
    wire N__12669;
    wire N__12666;
    wire N__12663;
    wire N__12660;
    wire N__12657;
    wire N__12654;
    wire N__12647;
    wire N__12644;
    wire N__12643;
    wire N__12642;
    wire N__12639;
    wire N__12636;
    wire N__12633;
    wire N__12630;
    wire N__12627;
    wire N__12624;
    wire N__12617;
    wire N__12614;
    wire N__12613;
    wire N__12612;
    wire N__12609;
    wire N__12606;
    wire N__12603;
    wire N__12600;
    wire N__12597;
    wire N__12594;
    wire N__12587;
    wire N__12584;
    wire N__12583;
    wire N__12582;
    wire N__12579;
    wire N__12576;
    wire N__12573;
    wire N__12570;
    wire N__12567;
    wire N__12564;
    wire N__12557;
    wire N__12556;
    wire N__12553;
    wire N__12550;
    wire N__12545;
    wire N__12542;
    wire N__12541;
    wire N__12538;
    wire N__12535;
    wire N__12532;
    wire N__12529;
    wire N__12526;
    wire N__12523;
    wire N__12520;
    wire N__12515;
    wire N__12512;
    wire N__12509;
    wire N__12506;
    wire N__12503;
    wire N__12500;
    wire N__12499;
    wire N__12498;
    wire N__12497;
    wire N__12496;
    wire N__12495;
    wire N__12494;
    wire N__12493;
    wire N__12492;
    wire N__12487;
    wire N__12474;
    wire N__12473;
    wire N__12470;
    wire N__12467;
    wire N__12464;
    wire N__12461;
    wire N__12452;
    wire N__12449;
    wire N__12448;
    wire N__12443;
    wire N__12440;
    wire N__12439;
    wire N__12438;
    wire N__12437;
    wire N__12434;
    wire N__12431;
    wire N__12428;
    wire N__12427;
    wire N__12426;
    wire N__12423;
    wire N__12422;
    wire N__12421;
    wire N__12418;
    wire N__12405;
    wire N__12402;
    wire N__12395;
    wire N__12392;
    wire N__12389;
    wire N__12386;
    wire N__12383;
    wire N__12380;
    wire N__12377;
    wire N__12374;
    wire N__12371;
    wire N__12368;
    wire N__12365;
    wire N__12362;
    wire N__12359;
    wire N__12356;
    wire N__12353;
    wire N__12350;
    wire N__12349;
    wire N__12346;
    wire N__12343;
    wire N__12338;
    wire N__12337;
    wire N__12334;
    wire N__12331;
    wire N__12326;
    wire N__12325;
    wire N__12322;
    wire N__12319;
    wire N__12314;
    wire N__12313;
    wire N__12310;
    wire N__12307;
    wire N__12302;
    wire N__12301;
    wire N__12298;
    wire N__12295;
    wire N__12292;
    wire N__12287;
    wire N__12284;
    wire N__12281;
    wire N__12278;
    wire N__12277;
    wire N__12276;
    wire N__12273;
    wire N__12266;
    wire N__12265;
    wire N__12264;
    wire N__12261;
    wire N__12258;
    wire N__12255;
    wire N__12252;
    wire N__12245;
    wire N__12242;
    wire N__12241;
    wire N__12238;
    wire N__12237;
    wire N__12236;
    wire N__12235;
    wire N__12234;
    wire N__12233;
    wire N__12232;
    wire N__12229;
    wire N__12226;
    wire N__12221;
    wire N__12216;
    wire N__12211;
    wire N__12200;
    wire N__12199;
    wire N__12198;
    wire N__12195;
    wire N__12194;
    wire N__12193;
    wire N__12188;
    wire N__12181;
    wire N__12176;
    wire N__12173;
    wire N__12172;
    wire N__12167;
    wire N__12166;
    wire N__12165;
    wire N__12162;
    wire N__12161;
    wire N__12160;
    wire N__12159;
    wire N__12158;
    wire N__12157;
    wire N__12154;
    wire N__12153;
    wire N__12150;
    wire N__12147;
    wire N__12142;
    wire N__12135;
    wire N__12130;
    wire N__12119;
    wire N__12118;
    wire N__12117;
    wire N__12116;
    wire N__12115;
    wire N__12114;
    wire N__12109;
    wire N__12100;
    wire N__12095;
    wire N__12092;
    wire N__12089;
    wire N__12088;
    wire N__12085;
    wire N__12082;
    wire N__12081;
    wire N__12080;
    wire N__12079;
    wire N__12076;
    wire N__12071;
    wire N__12066;
    wire N__12059;
    wire N__12058;
    wire N__12057;
    wire N__12056;
    wire N__12053;
    wire N__12050;
    wire N__12045;
    wire N__12038;
    wire N__12035;
    wire N__12034;
    wire N__12033;
    wire N__12030;
    wire N__12025;
    wire N__12020;
    wire N__12017;
    wire N__12014;
    wire N__12013;
    wire N__12012;
    wire N__12011;
    wire N__12010;
    wire N__12009;
    wire N__12008;
    wire N__12007;
    wire N__12004;
    wire N__11989;
    wire N__11984;
    wire N__11981;
    wire N__11978;
    wire N__11977;
    wire N__11976;
    wire N__11975;
    wire N__11974;
    wire N__11973;
    wire N__11972;
    wire N__11971;
    wire N__11968;
    wire N__11953;
    wire N__11948;
    wire N__11947;
    wire N__11946;
    wire N__11945;
    wire N__11944;
    wire N__11941;
    wire N__11938;
    wire N__11935;
    wire N__11932;
    wire N__11929;
    wire N__11926;
    wire N__11925;
    wire N__11924;
    wire N__11923;
    wire N__11914;
    wire N__11911;
    wire N__11908;
    wire N__11905;
    wire N__11902;
    wire N__11897;
    wire N__11890;
    wire N__11887;
    wire N__11882;
    wire N__11879;
    wire N__11876;
    wire N__11873;
    wire N__11870;
    wire N__11869;
    wire N__11868;
    wire N__11867;
    wire N__11864;
    wire N__11857;
    wire N__11852;
    wire N__11849;
    wire N__11846;
    wire N__11845;
    wire N__11844;
    wire N__11841;
    wire N__11838;
    wire N__11835;
    wire N__11834;
    wire N__11833;
    wire N__11832;
    wire N__11829;
    wire N__11826;
    wire N__11823;
    wire N__11816;
    wire N__11813;
    wire N__11810;
    wire N__11801;
    wire N__11798;
    wire N__11795;
    wire N__11794;
    wire N__11791;
    wire N__11788;
    wire N__11787;
    wire N__11784;
    wire N__11779;
    wire N__11776;
    wire N__11773;
    wire N__11768;
    wire N__11765;
    wire N__11764;
    wire N__11761;
    wire N__11760;
    wire N__11759;
    wire N__11756;
    wire N__11755;
    wire N__11752;
    wire N__11747;
    wire N__11742;
    wire N__11735;
    wire N__11732;
    wire N__11729;
    wire N__11726;
    wire N__11723;
    wire N__11720;
    wire N__11717;
    wire N__11714;
    wire N__11713;
    wire N__11710;
    wire N__11707;
    wire N__11706;
    wire N__11701;
    wire N__11698;
    wire N__11695;
    wire N__11690;
    wire N__11689;
    wire N__11688;
    wire N__11683;
    wire N__11680;
    wire N__11675;
    wire N__11672;
    wire N__11671;
    wire N__11670;
    wire N__11669;
    wire N__11662;
    wire N__11659;
    wire N__11654;
    wire N__11653;
    wire N__11650;
    wire N__11647;
    wire N__11644;
    wire N__11639;
    wire N__11636;
    wire N__11635;
    wire N__11632;
    wire N__11629;
    wire N__11626;
    wire N__11623;
    wire N__11620;
    wire N__11617;
    wire N__11614;
    wire N__11609;
    wire N__11606;
    wire N__11603;
    wire N__11600;
    wire N__11597;
    wire N__11594;
    wire N__11591;
    wire N__11590;
    wire N__11589;
    wire N__11588;
    wire N__11583;
    wire N__11578;
    wire N__11573;
    wire N__11572;
    wire N__11571;
    wire N__11570;
    wire N__11565;
    wire N__11560;
    wire N__11555;
    wire N__11552;
    wire N__11551;
    wire N__11550;
    wire N__11547;
    wire N__11540;
    wire N__11537;
    wire N__11536;
    wire N__11533;
    wire N__11530;
    wire N__11525;
    wire N__11522;
    wire N__11519;
    wire N__11516;
    wire N__11513;
    wire N__11512;
    wire N__11511;
    wire N__11510;
    wire N__11507;
    wire N__11506;
    wire N__11503;
    wire N__11500;
    wire N__11497;
    wire N__11494;
    wire N__11491;
    wire N__11488;
    wire N__11485;
    wire N__11474;
    wire N__11473;
    wire N__11472;
    wire N__11471;
    wire N__11468;
    wire N__11465;
    wire N__11462;
    wire N__11459;
    wire N__11458;
    wire N__11455;
    wire N__11452;
    wire N__11449;
    wire N__11446;
    wire N__11443;
    wire N__11438;
    wire N__11429;
    wire N__11428;
    wire N__11427;
    wire N__11426;
    wire N__11423;
    wire N__11420;
    wire N__11419;
    wire N__11416;
    wire N__11413;
    wire N__11410;
    wire N__11407;
    wire N__11404;
    wire N__11401;
    wire N__11390;
    wire N__11389;
    wire N__11388;
    wire N__11387;
    wire N__11386;
    wire N__11383;
    wire N__11380;
    wire N__11377;
    wire N__11374;
    wire N__11371;
    wire N__11368;
    wire N__11365;
    wire N__11362;
    wire N__11359;
    wire N__11356;
    wire N__11345;
    wire N__11344;
    wire N__11341;
    wire N__11338;
    wire N__11337;
    wire N__11334;
    wire N__11331;
    wire N__11328;
    wire N__11327;
    wire N__11326;
    wire N__11319;
    wire N__11314;
    wire N__11309;
    wire N__11308;
    wire N__11305;
    wire N__11304;
    wire N__11303;
    wire N__11300;
    wire N__11297;
    wire N__11294;
    wire N__11293;
    wire N__11290;
    wire N__11287;
    wire N__11284;
    wire N__11281;
    wire N__11278;
    wire N__11267;
    wire N__11264;
    wire N__11263;
    wire N__11262;
    wire N__11259;
    wire N__11256;
    wire N__11253;
    wire N__11250;
    wire N__11247;
    wire N__11244;
    wire N__11243;
    wire N__11242;
    wire N__11235;
    wire N__11232;
    wire N__11229;
    wire N__11222;
    wire N__11221;
    wire N__11218;
    wire N__11217;
    wire N__11214;
    wire N__11213;
    wire N__11210;
    wire N__11207;
    wire N__11204;
    wire N__11203;
    wire N__11200;
    wire N__11197;
    wire N__11194;
    wire N__11191;
    wire N__11188;
    wire N__11185;
    wire N__11178;
    wire N__11175;
    wire N__11168;
    wire N__11167;
    wire N__11164;
    wire N__11163;
    wire N__11160;
    wire N__11157;
    wire N__11156;
    wire N__11155;
    wire N__11152;
    wire N__11149;
    wire N__11146;
    wire N__11143;
    wire N__11140;
    wire N__11129;
    wire N__11126;
    wire N__11125;
    wire N__11122;
    wire N__11121;
    wire N__11118;
    wire N__11115;
    wire N__11112;
    wire N__11109;
    wire N__11102;
    wire N__11099;
    wire N__11098;
    wire N__11095;
    wire N__11094;
    wire N__11091;
    wire N__11088;
    wire N__11085;
    wire N__11082;
    wire N__11075;
    wire N__11074;
    wire N__11071;
    wire N__11070;
    wire N__11067;
    wire N__11064;
    wire N__11061;
    wire N__11060;
    wire N__11057;
    wire N__11056;
    wire N__11051;
    wire N__11048;
    wire N__11045;
    wire N__11042;
    wire N__11033;
    wire N__11032;
    wire N__11029;
    wire N__11026;
    wire N__11023;
    wire N__11022;
    wire N__11021;
    wire N__11018;
    wire N__11015;
    wire N__11012;
    wire N__11011;
    wire N__11008;
    wire N__11003;
    wire N__11000;
    wire N__10997;
    wire N__10988;
    wire N__10985;
    wire N__10984;
    wire N__10981;
    wire N__10980;
    wire N__10977;
    wire N__10974;
    wire N__10971;
    wire N__10968;
    wire N__10963;
    wire N__10958;
    wire N__10955;
    wire N__10954;
    wire N__10951;
    wire N__10950;
    wire N__10947;
    wire N__10946;
    wire N__10943;
    wire N__10942;
    wire N__10939;
    wire N__10936;
    wire N__10933;
    wire N__10930;
    wire N__10927;
    wire N__10916;
    wire N__10913;
    wire N__10910;
    wire N__10909;
    wire N__10906;
    wire N__10905;
    wire N__10902;
    wire N__10899;
    wire N__10896;
    wire N__10893;
    wire N__10886;
    wire N__10885;
    wire N__10884;
    wire N__10881;
    wire N__10878;
    wire N__10875;
    wire N__10872;
    wire N__10871;
    wire N__10870;
    wire N__10865;
    wire N__10862;
    wire N__10859;
    wire N__10856;
    wire N__10847;
    wire N__10846;
    wire N__10845;
    wire N__10842;
    wire N__10839;
    wire N__10836;
    wire N__10833;
    wire N__10830;
    wire N__10829;
    wire N__10828;
    wire N__10825;
    wire N__10822;
    wire N__10819;
    wire N__10816;
    wire N__10813;
    wire N__10802;
    wire N__10801;
    wire N__10798;
    wire N__10795;
    wire N__10794;
    wire N__10793;
    wire N__10790;
    wire N__10787;
    wire N__10784;
    wire N__10783;
    wire N__10780;
    wire N__10777;
    wire N__10774;
    wire N__10771;
    wire N__10768;
    wire N__10757;
    wire N__10756;
    wire N__10753;
    wire N__10752;
    wire N__10749;
    wire N__10746;
    wire N__10743;
    wire N__10740;
    wire N__10735;
    wire N__10730;
    wire N__10727;
    wire N__10724;
    wire N__10721;
    wire N__10718;
    wire N__10715;
    wire N__10712;
    wire N__10709;
    wire N__10706;
    wire N__10705;
    wire N__10702;
    wire N__10701;
    wire N__10700;
    wire N__10697;
    wire N__10696;
    wire N__10695;
    wire N__10692;
    wire N__10689;
    wire N__10688;
    wire N__10685;
    wire N__10682;
    wire N__10681;
    wire N__10680;
    wire N__10679;
    wire N__10678;
    wire N__10673;
    wire N__10668;
    wire N__10665;
    wire N__10662;
    wire N__10659;
    wire N__10654;
    wire N__10649;
    wire N__10646;
    wire N__10641;
    wire N__10628;
    wire N__10625;
    wire N__10622;
    wire N__10619;
    wire N__10616;
    wire N__10613;
    wire N__10612;
    wire N__10611;
    wire N__10610;
    wire N__10607;
    wire N__10604;
    wire N__10601;
    wire N__10598;
    wire N__10589;
    wire N__10586;
    wire N__10583;
    wire N__10580;
    wire N__10577;
    wire N__10574;
    wire N__10571;
    wire N__10570;
    wire N__10569;
    wire N__10568;
    wire N__10567;
    wire N__10564;
    wire N__10563;
    wire N__10562;
    wire N__10559;
    wire N__10558;
    wire N__10557;
    wire N__10554;
    wire N__10553;
    wire N__10548;
    wire N__10547;
    wire N__10546;
    wire N__10545;
    wire N__10544;
    wire N__10543;
    wire N__10542;
    wire N__10541;
    wire N__10540;
    wire N__10537;
    wire N__10534;
    wire N__10531;
    wire N__10528;
    wire N__10519;
    wire N__10518;
    wire N__10517;
    wire N__10516;
    wire N__10515;
    wire N__10514;
    wire N__10513;
    wire N__10512;
    wire N__10511;
    wire N__10510;
    wire N__10507;
    wire N__10494;
    wire N__10489;
    wire N__10482;
    wire N__10477;
    wire N__10472;
    wire N__10467;
    wire N__10456;
    wire N__10451;
    wire N__10444;
    wire N__10433;
    wire N__10432;
    wire N__10431;
    wire N__10430;
    wire N__10429;
    wire N__10428;
    wire N__10427;
    wire N__10426;
    wire N__10425;
    wire N__10420;
    wire N__10419;
    wire N__10414;
    wire N__10411;
    wire N__10406;
    wire N__10401;
    wire N__10398;
    wire N__10395;
    wire N__10392;
    wire N__10383;
    wire N__10376;
    wire N__10373;
    wire N__10370;
    wire N__10367;
    wire N__10364;
    wire N__10361;
    wire N__10358;
    wire N__10355;
    wire N__10352;
    wire N__10351;
    wire N__10350;
    wire N__10349;
    wire N__10346;
    wire N__10343;
    wire N__10340;
    wire N__10337;
    wire N__10334;
    wire N__10333;
    wire N__10330;
    wire N__10327;
    wire N__10324;
    wire N__10321;
    wire N__10318;
    wire N__10315;
    wire N__10312;
    wire N__10307;
    wire N__10302;
    wire N__10295;
    wire N__10294;
    wire N__10291;
    wire N__10288;
    wire N__10287;
    wire N__10286;
    wire N__10283;
    wire N__10282;
    wire N__10279;
    wire N__10276;
    wire N__10273;
    wire N__10270;
    wire N__10267;
    wire N__10264;
    wire N__10259;
    wire N__10250;
    wire N__10247;
    wire N__10246;
    wire N__10243;
    wire N__10242;
    wire N__10239;
    wire N__10236;
    wire N__10233;
    wire N__10230;
    wire N__10223;
    wire N__10220;
    wire N__10217;
    wire N__10214;
    wire N__10211;
    wire N__10210;
    wire N__10209;
    wire N__10208;
    wire N__10207;
    wire N__10206;
    wire N__10203;
    wire N__10198;
    wire N__10191;
    wire N__10184;
    wire N__10183;
    wire N__10182;
    wire N__10175;
    wire N__10172;
    wire N__10171;
    wire N__10168;
    wire N__10165;
    wire N__10164;
    wire N__10161;
    wire N__10158;
    wire N__10157;
    wire N__10154;
    wire N__10151;
    wire N__10148;
    wire N__10145;
    wire N__10144;
    wire N__10143;
    wire N__10140;
    wire N__10137;
    wire N__10134;
    wire N__10131;
    wire N__10126;
    wire N__10123;
    wire N__10120;
    wire N__10117;
    wire N__10106;
    wire N__10103;
    wire N__10100;
    wire N__10097;
    wire N__10094;
    wire N__10091;
    wire N__10088;
    wire N__10085;
    wire N__10082;
    wire N__10079;
    wire N__10076;
    wire N__10073;
    wire N__10070;
    wire N__10067;
    wire N__10064;
    wire N__10061;
    wire N__10058;
    wire N__10055;
    wire N__10052;
    wire N__10049;
    wire N__10046;
    wire N__10043;
    wire N__10040;
    wire N__10037;
    wire N__10034;
    wire N__10031;
    wire N__10028;
    wire N__10027;
    wire N__10024;
    wire N__10023;
    wire N__10020;
    wire N__10017;
    wire N__10014;
    wire N__10011;
    wire N__10008;
    wire N__10005;
    wire N__10002;
    wire N__9995;
    wire N__9992;
    wire N__9989;
    wire N__9986;
    wire N__9983;
    wire N__9980;
    wire N__9977;
    wire N__9974;
    wire N__9971;
    wire N__9970;
    wire N__9967;
    wire N__9964;
    wire N__9959;
    wire N__9956;
    wire N__9953;
    wire N__9950;
    wire N__9947;
    wire N__9946;
    wire N__9943;
    wire N__9940;
    wire N__9935;
    wire N__9932;
    wire N__9929;
    wire N__9926;
    wire N__9923;
    wire N__9920;
    wire N__9917;
    wire N__9914;
    wire N__9911;
    wire N__9908;
    wire N__9905;
    wire N__9902;
    wire N__9899;
    wire N__9896;
    wire N__9893;
    wire N__9890;
    wire N__9887;
    wire N__9884;
    wire N__9881;
    wire N__9878;
    wire N__9875;
    wire N__9872;
    wire N__9871;
    wire N__9868;
    wire N__9865;
    wire N__9862;
    wire N__9859;
    wire N__9854;
    wire N__9853;
    wire N__9850;
    wire N__9847;
    wire N__9844;
    wire N__9841;
    wire N__9836;
    wire N__9835;
    wire N__9832;
    wire N__9829;
    wire N__9826;
    wire N__9823;
    wire N__9818;
    wire N__9817;
    wire N__9814;
    wire N__9811;
    wire N__9808;
    wire N__9805;
    wire N__9802;
    wire N__9797;
    wire N__9796;
    wire N__9793;
    wire N__9790;
    wire N__9787;
    wire N__9784;
    wire N__9781;
    wire N__9776;
    wire N__9775;
    wire N__9772;
    wire N__9769;
    wire N__9766;
    wire N__9763;
    wire N__9760;
    wire N__9757;
    wire N__9752;
    wire N__9751;
    wire N__9748;
    wire N__9745;
    wire N__9742;
    wire N__9739;
    wire N__9736;
    wire N__9731;
    wire N__9728;
    wire N__9727;
    wire N__9724;
    wire N__9721;
    wire N__9716;
    wire N__9713;
    wire N__9710;
    wire N__9707;
    wire N__9704;
    wire N__9701;
    wire N__9698;
    wire N__9695;
    wire N__9692;
    wire N__9689;
    wire N__9686;
    wire N__9683;
    wire N__9680;
    wire N__9677;
    wire N__9674;
    wire N__9671;
    wire N__9670;
    wire N__9669;
    wire N__9668;
    wire N__9663;
    wire N__9660;
    wire N__9657;
    wire N__9650;
    wire N__9647;
    wire N__9644;
    wire N__9641;
    wire N__9638;
    wire N__9635;
    wire N__9632;
    wire N__9629;
    wire N__9628;
    wire N__9625;
    wire N__9622;
    wire N__9619;
    wire N__9616;
    wire N__9611;
    wire N__9608;
    wire N__9605;
    wire N__9604;
    wire N__9601;
    wire N__9598;
    wire N__9593;
    wire N__9590;
    wire N__9589;
    wire N__9586;
    wire N__9583;
    wire N__9580;
    wire N__9575;
    wire N__9572;
    wire N__9569;
    wire N__9566;
    wire N__9563;
    wire N__9560;
    wire N__9557;
    wire N__9554;
    wire N__9551;
    wire N__9548;
    wire N__9545;
    wire N__9542;
    wire N__9539;
    wire N__9536;
    wire N__9533;
    wire N__9530;
    wire N__9527;
    wire N__9526;
    wire N__9523;
    wire N__9520;
    wire N__9517;
    wire N__9512;
    wire N__9511;
    wire N__9510;
    wire N__9509;
    wire N__9506;
    wire N__9499;
    wire N__9494;
    wire N__9491;
    wire N__9488;
    wire N__9485;
    wire N__9484;
    wire N__9483;
    wire N__9482;
    wire N__9479;
    wire N__9472;
    wire N__9467;
    wire N__9464;
    wire N__9461;
    wire N__9458;
    wire N__9455;
    wire N__9454;
    wire N__9453;
    wire N__9452;
    wire N__9447;
    wire N__9444;
    wire N__9441;
    wire N__9436;
    wire N__9431;
    wire N__9428;
    wire N__9427;
    wire N__9426;
    wire N__9425;
    wire N__9422;
    wire N__9419;
    wire N__9414;
    wire N__9407;
    wire N__9404;
    wire N__9401;
    wire N__9398;
    wire N__9397;
    wire N__9396;
    wire N__9393;
    wire N__9392;
    wire N__9389;
    wire N__9386;
    wire N__9383;
    wire N__9380;
    wire N__9371;
    wire N__9368;
    wire N__9365;
    wire N__9362;
    wire N__9359;
    wire N__9356;
    wire N__9353;
    wire N__9350;
    wire N__9347;
    wire N__9344;
    wire N__9341;
    wire N__9340;
    wire N__9339;
    wire N__9338;
    wire N__9337;
    wire N__9336;
    wire N__9323;
    wire N__9320;
    wire N__9317;
    wire N__9314;
    wire N__9311;
    wire N__9310;
    wire N__9309;
    wire N__9308;
    wire N__9305;
    wire N__9302;
    wire N__9297;
    wire N__9290;
    wire N__9287;
    wire N__9284;
    wire N__9283;
    wire N__9282;
    wire N__9281;
    wire N__9278;
    wire N__9271;
    wire N__9266;
    wire N__9263;
    wire N__9262;
    wire N__9259;
    wire N__9258;
    wire N__9257;
    wire N__9252;
    wire N__9249;
    wire N__9246;
    wire N__9239;
    wire N__9236;
    wire N__9235;
    wire N__9234;
    wire N__9233;
    wire N__9230;
    wire N__9223;
    wire N__9218;
    wire N__9215;
    wire N__9212;
    wire N__9209;
    wire N__9208;
    wire N__9207;
    wire N__9206;
    wire N__9203;
    wire N__9196;
    wire N__9191;
    wire N__9188;
    wire N__9187;
    wire N__9186;
    wire N__9185;
    wire N__9182;
    wire N__9179;
    wire N__9174;
    wire N__9167;
    wire N__9164;
    wire N__9161;
    wire N__9158;
    wire N__9157;
    wire N__9156;
    wire N__9155;
    wire N__9152;
    wire N__9149;
    wire N__9144;
    wire N__9137;
    wire N__9134;
    wire N__9131;
    wire N__9128;
    wire N__9125;
    wire N__9124;
    wire N__9119;
    wire N__9116;
    wire N__9113;
    wire N__9110;
    wire N__9107;
    wire N__9104;
    wire N__9101;
    wire N__9098;
    wire N__9095;
    wire N__9092;
    wire N__9089;
    wire N__9086;
    wire N__9083;
    wire N__9080;
    wire N__9077;
    wire N__9074;
    wire N__9071;
    wire N__9068;
    wire N__9065;
    wire N__9062;
    wire N__9059;
    wire N__9056;
    wire N__9053;
    wire N__9050;
    wire N__9047;
    wire N__9044;
    wire N__9041;
    wire N__9038;
    wire N__9035;
    wire N__9032;
    wire N__9029;
    wire N__9026;
    wire N__9023;
    wire N__9020;
    wire N__9017;
    wire N__9014;
    wire N__9011;
    wire N__9008;
    wire N__9005;
    wire N__9002;
    wire N__8999;
    wire N__8996;
    wire N__8993;
    wire N__8990;
    wire N__8987;
    wire N__8984;
    wire N__8981;
    wire N__8978;
    wire N__8975;
    wire N__8972;
    wire N__8969;
    wire N__8966;
    wire N__8963;
    wire N__8960;
    wire N__8959;
    wire N__8956;
    wire N__8953;
    wire N__8948;
    wire N__8945;
    wire N__8942;
    wire N__8939;
    wire N__8936;
    wire N__8933;
    wire N__8930;
    wire N__8927;
    wire N__8924;
    wire N__8921;
    wire N__8918;
    wire N__8915;
    wire N__8912;
    wire N__8909;
    wire N__8906;
    wire N__8903;
    wire N__8900;
    wire N__8897;
    wire N__8894;
    wire N__8891;
    wire N__8888;
    wire N__8885;
    wire N__8884;
    wire N__8883;
    wire N__8882;
    wire N__8881;
    wire N__8880;
    wire N__8879;
    wire N__8878;
    wire N__8873;
    wire N__8860;
    wire N__8855;
    wire N__8852;
    wire N__8849;
    wire N__8846;
    wire N__8843;
    wire N__8840;
    wire N__8837;
    wire N__8834;
    wire N__8831;
    wire N__8828;
    wire N__8825;
    wire N__8822;
    wire N__8819;
    wire N__8816;
    wire N__8813;
    wire N__8810;
    wire N__8807;
    wire N__8804;
    wire N__8801;
    wire N__8798;
    wire N__8795;
    wire N__8792;
    wire N__8789;
    wire N__8786;
    wire N__8783;
    wire N__8780;
    wire N__8777;
    wire N__8774;
    wire N__8771;
    wire N__8768;
    wire N__8765;
    wire N__8762;
    wire N__8759;
    wire N__8756;
    wire N__8753;
    wire N__8750;
    wire N__8747;
    wire N__8744;
    wire N__8741;
    wire N__8738;
    wire N__8735;
    wire N__8732;
    wire N__8729;
    wire N__8726;
    wire N__8723;
    wire N__8720;
    wire N__8717;
    wire N__8714;
    wire N__8711;
    wire N__8708;
    wire N__8705;
    wire N__8702;
    wire N__8699;
    wire N__8696;
    wire N__8693;
    wire N__8690;
    wire N__8687;
    wire N__8684;
    wire N__8681;
    wire N__8678;
    wire N__8675;
    wire N__8672;
    wire N__8669;
    wire N__8666;
    wire N__8663;
    wire N__8662;
    wire N__8659;
    wire N__8656;
    wire N__8653;
    wire N__8648;
    wire N__8647;
    wire N__8644;
    wire N__8641;
    wire N__8636;
    wire N__8635;
    wire N__8632;
    wire N__8629;
    wire N__8624;
    wire N__8623;
    wire N__8620;
    wire N__8617;
    wire N__8612;
    wire N__8609;
    wire N__8606;
    wire N__8603;
    wire N__8600;
    wire N__8597;
    wire N__8594;
    wire N__8591;
    wire N__8588;
    wire N__8585;
    wire N__8582;
    wire N__8579;
    wire N__8576;
    wire N__8573;
    wire N__8570;
    wire N__8567;
    wire N__8564;
    wire N__8561;
    wire N__8558;
    wire N__8555;
    wire N__8552;
    wire N__8549;
    wire N__8546;
    wire N__8543;
    wire N__8542;
    wire N__8539;
    wire N__8536;
    wire N__8535;
    wire N__8534;
    wire N__8533;
    wire N__8526;
    wire N__8521;
    wire N__8516;
    wire N__8513;
    wire N__8512;
    wire N__8511;
    wire N__8510;
    wire N__8509;
    wire N__8508;
    wire N__8505;
    wire N__8496;
    wire N__8493;
    wire N__8486;
    wire N__8483;
    wire N__8480;
    wire N__8477;
    wire N__8474;
    wire N__8471;
    wire N__8468;
    wire N__8465;
    wire N__8462;
    wire N__8461;
    wire N__8460;
    wire N__8457;
    wire N__8452;
    wire N__8447;
    wire N__8446;
    wire N__8445;
    wire N__8444;
    wire N__8441;
    wire N__8436;
    wire N__8433;
    wire N__8426;
    wire N__8425;
    wire N__8424;
    wire N__8423;
    wire N__8420;
    wire N__8415;
    wire N__8414;
    wire N__8413;
    wire N__8412;
    wire N__8411;
    wire N__8408;
    wire N__8403;
    wire N__8394;
    wire N__8387;
    wire N__8386;
    wire N__8383;
    wire N__8380;
    wire N__8379;
    wire N__8378;
    wire N__8373;
    wire N__8368;
    wire N__8363;
    wire N__8362;
    wire N__8359;
    wire N__8356;
    wire N__8355;
    wire N__8354;
    wire N__8353;
    wire N__8352;
    wire N__8351;
    wire N__8350;
    wire N__8341;
    wire N__8338;
    wire N__8331;
    wire N__8328;
    wire N__8321;
    wire N__8318;
    wire N__8315;
    wire N__8312;
    wire N__8309;
    wire N__8306;
    wire N__8303;
    wire N__8300;
    wire N__8297;
    wire N__8294;
    wire N__8291;
    wire N__8288;
    wire N__8285;
    wire N__8282;
    wire GNDG0;
    wire VCCG0;
    wire \b2v_inst.cuenta_pixel_RNO_0Z0Z_1 ;
    wire \b2v_inst.g0_10_a3_0_4 ;
    wire \b2v_inst.g0_10_a3_0_7_cascade_ ;
    wire \b2v_inst.g0_10_a3_0_5 ;
    wire \b2v_inst.g0_10_a3_5_cascade_ ;
    wire \b2v_inst.g0_10_a3_4 ;
    wire \b2v_inst.un1_cuenta_pixel_c6 ;
    wire \b2v_inst.un1_cuenta_pixel_c6_cascade_ ;
    wire \b2v_inst.cuenta_pixelZ0Z_7 ;
    wire \b2v_inst.cuenta_pixelZ0Z_2 ;
    wire \b2v_inst.N_6_i ;
    wire \b2v_inst.g0_6_1_cascade_ ;
    wire \b2v_inst.N_4 ;
    wire \b2v_inst.un11_cuenta_pixel_6_cascade_ ;
    wire \b2v_inst.un11_cuenta_pixel_6 ;
    wire \b2v_inst.cuenta_pixel_RNI3FD32_0Z0Z_5 ;
    wire \b2v_inst.cuenta_pixelZ0Z_3 ;
    wire \b2v_inst.un1_cuenta_pixel_c3 ;
    wire \b2v_inst.cuenta_pixelZ0Z_4 ;
    wire bfn_1_15_0_;
    wire \b2v_inst.eventos_cry_0 ;
    wire \b2v_inst.eventos_cry_1 ;
    wire \b2v_inst.eventos_cry_2 ;
    wire \b2v_inst.eventos_cry_3 ;
    wire \b2v_inst.eventos_cry_4 ;
    wire \b2v_inst.eventos_cry_5 ;
    wire \b2v_inst.eventos_cry_6 ;
    wire \b2v_inst.eventosZ0Z_3 ;
    wire \b2v_inst.eventosZ0Z_4 ;
    wire \b2v_inst.eventosZ0Z_0 ;
    wire \b2v_inst.eventosZ0Z_5 ;
    wire \b2v_inst.N_47_i ;
    wire \b2v_inst.reg_ancho_1_i_0 ;
    wire bfn_1_17_0_;
    wire \b2v_inst.reg_ancho_1_i_1 ;
    wire \b2v_inst.un3_valor_max1_cry_0 ;
    wire \b2v_inst.reg_ancho_1_i_2 ;
    wire \b2v_inst.un3_valor_max1_cry_1 ;
    wire \b2v_inst.reg_ancho_1_i_3 ;
    wire \b2v_inst.un3_valor_max1_cry_2 ;
    wire \b2v_inst.reg_ancho_1_i_4 ;
    wire \b2v_inst.un3_valor_max1_cry_3 ;
    wire \b2v_inst.reg_ancho_1_i_5 ;
    wire \b2v_inst.un3_valor_max1_cry_4 ;
    wire \b2v_inst.reg_ancho_1_i_6 ;
    wire \b2v_inst.un3_valor_max1_cry_5 ;
    wire \b2v_inst.reg_ancho_1_i_7 ;
    wire \b2v_inst.un3_valor_max1_cry_6 ;
    wire \b2v_inst.un3_valor_max1 ;
    wire bfn_1_18_0_;
    wire bfn_1_19_0_;
    wire \b2v_inst.valor_max_final5_3_cry_0 ;
    wire \b2v_inst.valor_max_final5_3_cry_1 ;
    wire \b2v_inst.valor_max_final5_3_cry_2 ;
    wire \b2v_inst.valor_max_final5_3_cry_3 ;
    wire \b2v_inst.valor_max_final5_3_cry_4 ;
    wire \b2v_inst.valor_max_final5_3_cry_5 ;
    wire \b2v_inst.valor_max_final5_3_cry_6 ;
    wire \b2v_inst.valor_max_final53 ;
    wire bfn_1_20_0_;
    wire \b2v_inst.g0_10_1 ;
    wire \b2v_inst.g0_10_a3_7 ;
    wire bfn_2_11_0_;
    wire \b2v_inst.un1_pix_count_anterior_0_data_tmp_0 ;
    wire \b2v_inst.un1_pix_count_anterior_0_data_tmp_1 ;
    wire \b2v_inst.un1_pix_count_anterior_0_data_tmp_2 ;
    wire \b2v_inst.un1_pix_count_anterior_0_data_tmp_3 ;
    wire \b2v_inst.un1_pix_count_anterior_0_data_tmp_4 ;
    wire \b2v_inst.un1_pix_count_anterior_0_data_tmp_5 ;
    wire \b2v_inst.un1_pix_count_anterior_0_N_2 ;
    wire \b2v_inst.un1_pix_count_anterior_0_I_15_c_RNOZ0 ;
    wire \b2v_inst.pix_count_anteriorZ0Z_4 ;
    wire \b2v_inst.pix_count_anteriorZ0Z_5 ;
    wire \b2v_inst.pix_count_anteriorZ0Z_1 ;
    wire \b2v_inst.un1_pix_count_anterior_0_I_1_c_RNOZ0 ;
    wire \b2v_inst.pix_count_anteriorZ0Z_0 ;
    wire \b2v_inst.pix_count_anteriorZ0Z_12 ;
    wire \b2v_inst.un1_pix_count_anterior_0_I_39_c_RNOZ0 ;
    wire \b2v_inst.un1_pix_count_anterior_0_I_21_c_RNOZ0 ;
    wire \b2v_inst.pix_count_anteriorZ0Z_6 ;
    wire \b2v_inst4.un1_pix_count_int_0_sqmuxa_8_cascade_ ;
    wire \b2v_inst.pix_count_anteriorZ0Z_7 ;
    wire \b2v_inst.pix_count_anteriorZ0Z_8 ;
    wire \b2v_inst.un1_pix_count_anterior_0_I_51_c_RNOZ0 ;
    wire \b2v_inst.pix_count_anteriorZ0Z_9 ;
    wire \b2v_inst.un1_state_17_0 ;
    wire \b2v_inst.ignorar_anchoZ0Z_1 ;
    wire \b2v_inst.data_a_escribir_RNO_3Z0Z_4_cascade_ ;
    wire \b2v_inst.data_a_escribir_RNO_3Z0Z_0_cascade_ ;
    wire \b2v_inst.un1_reg_anterior_iv_0_0_0_0 ;
    wire \b2v_inst.un1_m3_2_0 ;
    wire \b2v_inst.data_a_escribir_RNO_1Z0Z_0_cascade_ ;
    wire \b2v_inst.un1_reg_anterior_iv_0_0_1_1_3 ;
    wire \b2v_inst.N_315_cascade_ ;
    wire \b2v_inst.un1_reg_anterior_iv_0_0_1_3 ;
    wire \b2v_inst.un1_reg_anterior_iv_0_0_a2_6_0_1_cascade_ ;
    wire \b2v_inst.N_317 ;
    wire \b2v_inst.un1_reg_anterior_iv_0_0_a2_4_tz_1_2 ;
    wire \b2v_inst.eventosZ0Z_2 ;
    wire \b2v_inst.N_320_tz_cascade_ ;
    wire \b2v_inst.un1_m3_0_m3_ns_1_cascade_ ;
    wire \b2v_inst.N_318 ;
    wire \b2v_inst.data_a_escribir_RNO_0Z0Z_4 ;
    wire \b2v_inst.un1_reg_anterior_iv_0_0_0_4 ;
    wire N_211_i;
    wire N_219_i;
    wire N_217_i;
    wire N_215_i;
    wire \b2v_inst.state_ns_i_i_a2_4Z0Z_6 ;
    wire \b2v_inst.state_ns_i_i_a2_4Z0Z_6_cascade_ ;
    wire \b2v_inst.N_497_cascade_ ;
    wire \b2v_inst.N_361 ;
    wire \b2v_inst.state_ns_i_i_a2_5Z0Z_6 ;
    wire \b2v_inst.N_254_i ;
    wire \b2v_inst.pix_count_anteriorZ0Z_2 ;
    wire \b2v_inst.un1_pix_count_anterior_0_I_27_c_RNOZ0 ;
    wire \b2v_inst.pix_count_anteriorZ0Z_3 ;
    wire \b2v_inst.pix_count_anteriorZ0Z_10 ;
    wire \b2v_inst.un1_pix_count_anterior_0_I_9_c_RNOZ0 ;
    wire \b2v_inst.pix_count_anteriorZ0Z_11 ;
    wire \b2v_inst.N_254_i_g ;
    wire SYNTHESIZED_WIRE_2_0;
    wire \b2v_inst4.pix_count_int_RNO_0Z0Z_0 ;
    wire bfn_3_13_0_;
    wire SYNTHESIZED_WIRE_2_1;
    wire \b2v_inst4.un1_pix_count_int_cry_0 ;
    wire SYNTHESIZED_WIRE_2_2;
    wire \b2v_inst4.un1_pix_count_int_cry_1 ;
    wire SYNTHESIZED_WIRE_2_3;
    wire \b2v_inst4.pix_count_int_RNO_0Z0Z_3 ;
    wire \b2v_inst4.un1_pix_count_int_cry_2 ;
    wire SYNTHESIZED_WIRE_2_4;
    wire \b2v_inst4.un1_pix_count_int_cry_3 ;
    wire SYNTHESIZED_WIRE_2_5;
    wire \b2v_inst4.pix_count_int_RNO_0Z0Z_5 ;
    wire \b2v_inst4.un1_pix_count_int_cry_4 ;
    wire SYNTHESIZED_WIRE_2_6;
    wire \b2v_inst4.un1_pix_count_int_cry_5 ;
    wire SYNTHESIZED_WIRE_2_7;
    wire \b2v_inst4.pix_count_int_RNO_0Z0Z_7 ;
    wire \b2v_inst4.un1_pix_count_int_cry_6 ;
    wire \b2v_inst4.un1_pix_count_int_cry_7 ;
    wire SYNTHESIZED_WIRE_2_8;
    wire \b2v_inst4.pix_count_int_RNO_0Z0Z_8 ;
    wire bfn_3_14_0_;
    wire \b2v_inst4.un1_pix_count_int_cry_8 ;
    wire SYNTHESIZED_WIRE_2_10;
    wire \b2v_inst4.un1_pix_count_int_cry_9 ;
    wire SYNTHESIZED_WIRE_2_11;
    wire \b2v_inst4.pix_count_int_RNO_0Z0Z_11 ;
    wire \b2v_inst4.un1_pix_count_int_cry_10 ;
    wire SYNTHESIZED_WIRE_2_12;
    wire \b2v_inst4.un1_pix_count_int_cry_11 ;
    wire \b2v_inst4.pix_count_int_RNO_0Z0Z_12 ;
    wire \b2v_inst.data_a_escribir9_0_and ;
    wire bfn_3_15_0_;
    wire \b2v_inst.data_a_escribir9_1_and ;
    wire \b2v_inst.data_a_escribir9_0 ;
    wire \b2v_inst.data_a_escribir9_2_and ;
    wire \b2v_inst.data_a_escribir9_1 ;
    wire \b2v_inst.data_a_escribir9_3_and ;
    wire \b2v_inst.data_a_escribir9_2 ;
    wire \b2v_inst.data_a_escribir9_3 ;
    wire \b2v_inst.data_a_escribir9_4 ;
    wire \b2v_inst.data_a_escribir9_5 ;
    wire \b2v_inst.data_a_escribir9_6 ;
    wire \b2v_inst.data_a_escribir10 ;
    wire bfn_3_16_0_;
    wire \b2v_inst.eventosZ0Z_7 ;
    wire \b2v_inst.eventosZ0Z_1 ;
    wire \b2v_inst.eventosZ0Z_6 ;
    wire \b2v_inst.un1_reg_anterior_iv_0_0_2_1_1_cascade_ ;
    wire \b2v_inst.data_a_escribir_RNO_4Z0Z_1_cascade_ ;
    wire \b2v_inst.un1_reg_anterior_iv_0_0_0_1 ;
    wire \b2v_inst.data_a_escribir_RNO_0Z0Z_1 ;
    wire \b2v_inst.data_a_escribir_RNO_1Z0Z_1_cascade_ ;
    wire \b2v_inst.N_497 ;
    wire \b2v_inst.un1_reg_anterior_iv_0_0_2_tz_2 ;
    wire \b2v_inst.data_a_escribir_RNO_1Z0Z_2_cascade_ ;
    wire \b2v_inst.un1_reg_anterior_iv_0_0_1_2 ;
    wire \b2v_inst.data_a_escribir_RNO_4Z0Z_5_cascade_ ;
    wire \b2v_inst.un1_reg_anterior_iv_0_0_2_1_5_cascade_ ;
    wire \b2v_inst.un1_reg_anterior_iv_0_0_a2_4_0_1 ;
    wire \b2v_inst.un1_reg_anterior_iv_0_0_0_5 ;
    wire \b2v_inst.data_a_escribir_RNO_0Z0Z_5_cascade_ ;
    wire \b2v_inst.data_a_escribir_RNO_1Z0Z_5 ;
    wire \b2v_inst.reg_anterior_i_0 ;
    wire bfn_3_19_0_;
    wire \b2v_inst.reg_anterior_i_1 ;
    wire \b2v_inst.valor_max_final5_1_cry_0 ;
    wire \b2v_inst.reg_anterior_i_2 ;
    wire \b2v_inst.valor_max_final5_1_cry_1 ;
    wire \b2v_inst.reg_anterior_i_3 ;
    wire \b2v_inst.valor_max_final5_1_cry_2 ;
    wire \b2v_inst.reg_anterior_i_4 ;
    wire \b2v_inst.valor_max_final5_1_cry_3 ;
    wire \b2v_inst.reg_anterior_i_5 ;
    wire \b2v_inst.valor_max_final5_1_cry_4 ;
    wire \b2v_inst.reg_anterior_i_6 ;
    wire \b2v_inst.valor_max_final5_1_cry_5 ;
    wire \b2v_inst.reg_anterior_i_7 ;
    wire \b2v_inst.valor_max_final5_1_cry_6 ;
    wire \b2v_inst.valor_max_final51 ;
    wire \b2v_inst.valor_max_final53_THRU_CO ;
    wire \b2v_inst.un1_m3_0_m3_ns_1 ;
    wire bfn_3_20_0_;
    wire \b2v_inst.un1_reg_anterior_iv_0_0_2_tz_4 ;
    wire \b2v_inst3.fsm_state_ns_0_0_0_1_cascade_ ;
    wire N_230_cascade_;
    wire \b2v_inst3.N_434 ;
    wire \b2v_inst3.N_490 ;
    wire \b2v_inst3.fsm_state_ns_i_i_1_0_cascade_ ;
    wire \b2v_inst3.un1_m2_0_a2_2_cascade_ ;
    wire \b2v_inst3.un1_cycle_counter_5_c5 ;
    wire \b2v_inst3.un1_cycle_counter_5_c5_cascade_ ;
    wire SYNTHESIZED_WIRE_10_0;
    wire SYNTHESIZED_WIRE_3_0;
    wire SYNTHESIZED_WIRE_3_1;
    wire SYNTHESIZED_WIRE_3_2;
    wire SYNTHESIZED_WIRE_3_3;
    wire SYNTHESIZED_WIRE_3_4;
    wire SYNTHESIZED_WIRE_3_5;
    wire SYNTHESIZED_WIRE_3_6;
    wire SYNTHESIZED_WIRE_3_7;
    wire \b2v_inst4.pix_count_int_0_sqmuxa ;
    wire \b2v_inst.we_0_a2_0_a2_4_cascade_ ;
    wire SYNTHESIZED_WIRE_4;
    wire \b2v_inst.we_0_a2_0_a2_3 ;
    wire N_458_cascade_;
    wire \b2v_inst.N_429_cascade_ ;
    wire \b2v_inst.un1_pix_count_anterior_0_N_2_THRU_CO ;
    wire \b2v_inst.stateZ0Z_3 ;
    wire \b2v_inst.stateZ0Z_2 ;
    wire \b2v_inst.data_a_escribir9_4_and ;
    wire \b2v_inst.data_a_escribir9_5_and ;
    wire \b2v_inst.un3_valor_max1_THRU_CO ;
    wire \b2v_inst.data_a_escribir_RNO_3Z0Z_6 ;
    wire \b2v_inst.un1_reg_anterior_iv_0_0_a2_6_0_1 ;
    wire \b2v_inst.un1_m3_0_0 ;
    wire \b2v_inst.un1_reg_anterior_iv_0_0_0_6 ;
    wire \b2v_inst.data_a_escribir_RNO_1Z0Z_6_cascade_ ;
    wire \b2v_inst.data_a_escribir10_THRU_CO ;
    wire \b2v_inst.N_264 ;
    wire \b2v_inst.un1_reg_anterior_iv_0_0_0_7 ;
    wire \b2v_inst.un1_reg_anterior_iv_0_0_3_0_7_cascade_ ;
    wire \b2v_inst.un1_reg_anterior_iv_0_0_2_0_tz_7 ;
    wire \b2v_inst.un1_reset_inv_2_0 ;
    wire \b2v_inst.reg_ancho_1Z0Z_0 ;
    wire \b2v_inst.reg_ancho_3Z0Z_0 ;
    wire bfn_5_17_0_;
    wire \b2v_inst.reg_ancho_1Z0Z_1 ;
    wire \b2v_inst.reg_ancho_3Z0Z_1 ;
    wire \b2v_inst.valor_max_final5_0_cry_0 ;
    wire \b2v_inst.reg_ancho_3Z0Z_2 ;
    wire \b2v_inst.reg_ancho_1Z0Z_2 ;
    wire \b2v_inst.valor_max_final5_0_cry_1 ;
    wire \b2v_inst.reg_ancho_1Z0Z_3 ;
    wire \b2v_inst.reg_ancho_3Z0Z_3 ;
    wire \b2v_inst.valor_max_final5_0_cry_2 ;
    wire \b2v_inst.reg_ancho_1Z0Z_4 ;
    wire \b2v_inst.reg_ancho_3Z0Z_4 ;
    wire \b2v_inst.valor_max_final5_0_cry_3 ;
    wire \b2v_inst.reg_ancho_1Z0Z_5 ;
    wire \b2v_inst.valor_max_final5_0_cry_4 ;
    wire \b2v_inst.reg_ancho_1Z0Z_6 ;
    wire \b2v_inst.valor_max_final5_0_cry_5 ;
    wire \b2v_inst.reg_ancho_1Z0Z_7 ;
    wire \b2v_inst.reg_ancho_3Z0Z_7 ;
    wire \b2v_inst.valor_max_final5_0_cry_6 ;
    wire \b2v_inst.valor_max_final50 ;
    wire bfn_5_18_0_;
    wire \b2v_inst.valor_max_final50_THRU_CO ;
    wire \b2v_inst.data_a_escribir9_6_and ;
    wire \b2v_inst.reg_ancho_2Z0Z_0 ;
    wire bfn_5_19_0_;
    wire \b2v_inst.reg_ancho_2Z0Z_1 ;
    wire \b2v_inst.valor_max_final5_2_cry_0 ;
    wire \b2v_inst.reg_ancho_2Z0Z_2 ;
    wire \b2v_inst.valor_max_final5_2_cry_1 ;
    wire \b2v_inst.reg_ancho_2Z0Z_3 ;
    wire \b2v_inst.valor_max_final5_2_cry_2 ;
    wire \b2v_inst.reg_ancho_2Z0Z_4 ;
    wire \b2v_inst.valor_max_final5_2_cry_3 ;
    wire \b2v_inst.reg_ancho_2Z0Z_5 ;
    wire \b2v_inst.valor_max_final5_2_cry_4 ;
    wire \b2v_inst.reg_ancho_2Z0Z_6 ;
    wire \b2v_inst.valor_max_final5_2_cry_5 ;
    wire \b2v_inst.reg_ancho_2Z0Z_7 ;
    wire \b2v_inst.valor_max_final5_2_cry_6 ;
    wire \b2v_inst.valor_max_final52 ;
    wire bfn_5_20_0_;
    wire \b2v_inst.valor_max_final52_THRU_CO ;
    wire \b2v_inst3.un1_bit_counter_3_c2 ;
    wire \b2v_inst3.un1_bit_counter_3_c2_cascade_ ;
    wire \b2v_inst3.N_258 ;
    wire \b2v_inst3.N_258_cascade_ ;
    wire \b2v_inst3.bit_counterZ0Z_2 ;
    wire \b2v_inst3.bit_counterZ1Z_1 ;
    wire \b2v_inst3.N_102_2_cascade_ ;
    wire \b2v_inst3.bit_counterZ0Z_3 ;
    wire \b2v_inst3.N_436 ;
    wire uart_tx_o;
    wire \b2v_inst4.stateZ0Z_0 ;
    wire \b2v_inst3.cycle_counterZ0Z_6 ;
    wire \b2v_inst3.cycle_counterZ0Z_5 ;
    wire \b2v_inst3.cycle_counterZ0Z_7 ;
    wire \b2v_inst3.next_bit_0_a3_4_cascade_ ;
    wire \b2v_inst3.next_bit_0_a3_3 ;
    wire SYNTHESIZED_WIRE_7;
    wire \b2v_inst3.N_105_7_cascade_ ;
    wire \b2v_inst3.fsm_stateZ0Z_0 ;
    wire \b2v_inst3.cycle_counterZ0Z_1 ;
    wire \b2v_inst3.fsm_stateZ0Z_1 ;
    wire \b2v_inst3.cycle_counterZ0Z_0 ;
    wire \b2v_inst3.un1_cycle_counter_5_c2 ;
    wire \b2v_inst3.cycle_counterZ0Z_2 ;
    wire \b2v_inst3.cycle_counterZ0Z_3 ;
    wire \b2v_inst3.un1_cycle_counter_5_c2_cascade_ ;
    wire \b2v_inst3.cycle_counterZ0Z_4 ;
    wire \b2v_inst4.un1_pix_count_int_0_sqmuxa_9 ;
    wire \b2v_inst4.un1_pix_count_int_0_sqmuxa_11 ;
    wire \b2v_inst4.un1_pix_count_int_0_sqmuxa_10 ;
    wire \b2v_inst4.pix_count_int_RNO_0Z0Z_9 ;
    wire SYNTHESIZED_WIRE_2_9;
    wire \b2v_inst.cuenta_pixelZ0Z_6 ;
    wire \b2v_inst.un11_cuenta_pixel_i_0_o2_0 ;
    wire \b2v_inst.cuenta_pixelZ0Z_5 ;
    wire \b2v_inst.cuenta_pixelZ0Z_0 ;
    wire \b2v_inst.cuenta_pixelZ0Z_1 ;
    wire \b2v_inst.cuenta_pixel_4_i_a2_0_6 ;
    wire N_213_i;
    wire N_209_i;
    wire N_207_i;
    wire SYNTHESIZED_WIRE_10_2;
    wire SYNTHESIZED_WIRE_10_3;
    wire SYNTHESIZED_WIRE_10_4;
    wire SYNTHESIZED_WIRE_10_5;
    wire SYNTHESIZED_WIRE_10_6;
    wire SYNTHESIZED_WIRE_10_7;
    wire \b2v_inst.addr_ram_1_iv_i_2_5_cascade_ ;
    wire N_54;
    wire \b2v_inst.addr_ram_1_iv_i_1_5 ;
    wire \b2v_inst.N_341 ;
    wire \b2v_inst.N_404_cascade_ ;
    wire \b2v_inst.reg_ancho_3Z0Z_6 ;
    wire \b2v_inst.reg_ancho_3Z0Z_5 ;
    wire \b2v_inst.reg_ancho_3_i_0 ;
    wire bfn_6_17_0_;
    wire \b2v_inst.reg_ancho_3_i_1 ;
    wire \b2v_inst.un3_valor_max2_cry_0 ;
    wire \b2v_inst.reg_ancho_3_i_2 ;
    wire \b2v_inst.un3_valor_max2_cry_1 ;
    wire \b2v_inst.reg_ancho_3_i_3 ;
    wire \b2v_inst.un3_valor_max2_cry_2 ;
    wire \b2v_inst.reg_ancho_3_i_4 ;
    wire \b2v_inst.un3_valor_max2_cry_3 ;
    wire \b2v_inst.reg_ancho_3_i_5 ;
    wire \b2v_inst.un3_valor_max2_cry_4 ;
    wire \b2v_inst.reg_ancho_3_i_6 ;
    wire \b2v_inst.un3_valor_max2_cry_5 ;
    wire \b2v_inst.reg_ancho_3_i_7 ;
    wire \b2v_inst.un3_valor_max2_cry_6 ;
    wire \b2v_inst.un3_valor_max2 ;
    wire bfn_6_18_0_;
    wire \b2v_inst.un3_valor_max2_THRU_CO ;
    wire reset_i;
    wire \b2v_inst3.un2_n_fsm_state_0_sqmuxa_2_0_i ;
    wire \b2v_inst1.r_RX_Bytece_0_6 ;
    wire SYNTHESIZED_WIRE_1_0;
    wire \b2v_inst.reg_anteriorZ0Z_0 ;
    wire SYNTHESIZED_WIRE_1_1;
    wire \b2v_inst.reg_anteriorZ0Z_1 ;
    wire SYNTHESIZED_WIRE_1_2;
    wire \b2v_inst.reg_anteriorZ0Z_2 ;
    wire SYNTHESIZED_WIRE_1_3;
    wire \b2v_inst.reg_anteriorZ0Z_3 ;
    wire SYNTHESIZED_WIRE_1_7;
    wire \b2v_inst.reg_anteriorZ0Z_7 ;
    wire \b2v_inst.data_a_escribir9_7_and ;
    wire SYNTHESIZED_WIRE_1_4;
    wire \b2v_inst.reg_anteriorZ0Z_4 ;
    wire b2v_inst_data_a_escribir_1;
    wire b2v_inst_data_a_escribir_0;
    wire \b2v_inst3.data_to_sendZ0Z_1 ;
    wire \b2v_inst3.data_to_sendZ0Z_0 ;
    wire b2v_inst_data_a_escribir_2;
    wire \b2v_inst3.data_to_sendZ0Z_2 ;
    wire \b2v_inst3.fsm_state_RNIEPSN1Z0Z_0 ;
    wire \b2v_inst3.N_105_7 ;
    wire \b2v_inst3.bit_counterZ0Z_0 ;
    wire \b2v_inst.state_ns_a2_0_a2_0_1_2 ;
    wire \b2v_inst.cuenta_5_i_a2_2_0_1_cascade_ ;
    wire \b2v_inst.un4_cuenta_c4_cascade_ ;
    wire \b2v_inst.cuentaZ0Z_3 ;
    wire \b2v_inst.cuentaZ0Z_2 ;
    wire \b2v_inst.un2_cuentalto7_3_cascade_ ;
    wire \b2v_inst.N_351_0_cascade_ ;
    wire \b2v_inst.cuenta_fastZ0Z_4 ;
    wire \b2v_inst.cuenta_RNIQ56K_0Z0Z_3 ;
    wire \b2v_inst.N_376_1 ;
    wire \b2v_inst.cuenta_RNIQI4FZ0Z_2 ;
    wire \b2v_inst.cuenta_RNIR03AZ0Z_1 ;
    wire \b2v_inst.N_376_1_cascade_ ;
    wire \b2v_inst.cuentaZ0Z_1 ;
    wire \b2v_inst.cuenta_5_i_a2_0_3 ;
    wire \b2v_inst.cuentaZ0Z_0 ;
    wire \b2v_inst.N_377 ;
    wire \b2v_inst.N_491_cascade_ ;
    wire \b2v_inst.state_RNIFQKOZ0Z_17 ;
    wire \b2v_inst.state_RNIFQKOZ0Z_17_cascade_ ;
    wire \b2v_inst.N_236_cascade_ ;
    wire \b2v_inst.stateZ0Z_9 ;
    wire \b2v_inst.N_399_cascade_ ;
    wire \b2v_inst.addr_ram_1_iv_i_1_6 ;
    wire \b2v_inst.addr_ram_1_iv_i_2_6_cascade_ ;
    wire N_165;
    wire \b2v_inst.stateZ0Z_12 ;
    wire \b2v_inst.N_235_cascade_ ;
    wire \b2v_inst.stateZ0Z_11 ;
    wire \b2v_inst.N_237_cascade_ ;
    wire \b2v_inst.addr_ram_1_iv_i_2_0 ;
    wire \b2v_inst.addr_ram_1_iv_i_1_0_cascade_ ;
    wire N_167;
    wire \b2v_inst.addr_ram_1_0_iv_i_0_1 ;
    wire N_60;
    wire \b2v_inst.addr_ram_1_0_iv_i_0_2_cascade_ ;
    wire N_56;
    wire \b2v_inst.dir_mem_315_0_cascade_ ;
    wire \b2v_inst.dir_mem_3Z0Z_1 ;
    wire \b2v_inst.addr_ram_1_0_iv_i_1_1 ;
    wire \b2v_inst.dir_mem_3Z0Z_0 ;
    wire \b2v_inst.dir_mem_3Z0Z_5 ;
    wire \b2v_inst.dir_mem_3Z0Z_6 ;
    wire N_205_i;
    wire \b2v_inst.dir_mem_2Z0Z_6 ;
    wire \b2v_inst1.r_RX_Bytece_0_3 ;
    wire \b2v_inst1.r_RX_Bytece_0_0_4 ;
    wire b2v_inst_data_a_escribir_3;
    wire \b2v_inst3.data_to_sendZ0Z_3 ;
    wire b2v_inst_data_a_escribir_4;
    wire \b2v_inst3.data_to_sendZ0Z_4 ;
    wire b2v_inst_data_a_escribir_5;
    wire \b2v_inst3.data_to_sendZ0Z_5 ;
    wire b2v_inst_data_a_escribir_6;
    wire \b2v_inst3.data_to_sendZ0Z_6 ;
    wire N_458;
    wire b2v_inst_data_a_escribir_7;
    wire N_230;
    wire \b2v_inst3.data_to_sendZ0Z_7 ;
    wire \b2v_inst3.un2_n_fsm_state_0_sqmuxa_2_0_i_0 ;
    wire SYNTHESIZED_WIRE_1_6;
    wire \b2v_inst.reg_anteriorZ0Z_6 ;
    wire SYNTHESIZED_WIRE_1_5;
    wire \b2v_inst.reg_anteriorZ0Z_5 ;
    wire \b2v_inst.un4_cuenta_ac0_11_0_cascade_ ;
    wire \b2v_inst.N_491 ;
    wire \b2v_inst.cuenta_5_i_o2_0_0_1_cascade_ ;
    wire \b2v_inst.state_ns_a2_0_o2_1_0_2_cascade_ ;
    wire \b2v_inst.cuenta_5_i_o2_0_0_1 ;
    wire \b2v_inst.state_17_rep1_RNICDKZ0Z34_cascade_ ;
    wire \b2v_inst.cuenta_RNIO2VO3Z0Z_4 ;
    wire \b2v_inst.N_374 ;
    wire \b2v_inst.cuentaZ0Z_5 ;
    wire \b2v_inst.cuentaZ0Z_4 ;
    wire \b2v_inst.un4_cuenta_ac0_9_0_cascade_ ;
    wire \b2v_inst.un4_cuenta_c4 ;
    wire \b2v_inst.cuentaZ0Z_6 ;
    wire \b2v_inst.cuentaZ0Z_7 ;
    wire \b2v_inst.N_399_i ;
    wire \b2v_inst.N_227 ;
    wire \b2v_inst.N_232 ;
    wire \b2v_inst.N_232_cascade_ ;
    wire \b2v_inst.stateZ0Z_7 ;
    wire \b2v_inst.stateZ0Z_14 ;
    wire \b2v_inst.stateZ0Z_6 ;
    wire \b2v_inst.state_RNITETBZ0Z_0 ;
    wire \b2v_inst.N_351_cascade_ ;
    wire \b2v_inst.addr_ram_1_iv_i_1_3 ;
    wire \b2v_inst.addr_ram_1_iv_i_2_3_cascade_ ;
    wire N_58;
    wire \b2v_inst.stateZ0Z_0 ;
    wire \b2v_inst.stateZ0Z_10 ;
    wire \b2v_inst.stateZ0Z_1 ;
    wire \b2v_inst.dir_mem_3Z0Z_4 ;
    wire \b2v_inst.addr_ram_1_0_iv_i_1_4_cascade_ ;
    wire N_163;
    wire \b2v_inst.g0_11_1_cascade_ ;
    wire \b2v_inst.dir_mem_1Z0Z_4 ;
    wire \b2v_inst.N_235 ;
    wire \b2v_inst.addr_ram_1_0_iv_i_0_4 ;
    wire \b2v_inst.dir_mem_315_0 ;
    wire \b2v_inst.dir_mem_3Z0Z_3 ;
    wire \b2v_inst.dir_mem_3Z0Z_7 ;
    wire \b2v_inst.N_138_i ;
    wire \b2v_inst1.r_RX_Bytece_0_5 ;
    wire \b2v_inst.dir_mem_3_RNO_0Z0Z_3 ;
    wire \b2v_inst1.r_RX_Bytece_0_0_1_cascade_ ;
    wire SYNTHESIZED_WIRE_10_1;
    wire \b2v_inst.dir_mem_2_RNO_0Z0Z_6 ;
    wire SYNTHESIZED_WIRE_9;
    wire \b2v_inst.stateZ0Z_16 ;
    wire \b2v_inst.ignorar_anteriorZ0 ;
    wire \b2v_inst.un1_state_19_0 ;
    wire \b2v_inst.N_5 ;
    wire \b2v_inst.N_7_1_cascade_ ;
    wire \b2v_inst.g2_2_cascade_ ;
    wire \b2v_inst.g1 ;
    wire \b2v_inst.un2_indice_21_s0_0_6 ;
    wire \b2v_inst.N_253_cascade_ ;
    wire \b2v_inst.state_fastZ0Z_17 ;
    wire \b2v_inst.state_fastZ0Z_15 ;
    wire \b2v_inst.N_253_i_cascade_ ;
    wire \b2v_inst.un2_indice_3_0_iv_0_a2_5_sx_2 ;
    wire \b2v_inst.N_452_cascade_ ;
    wire \b2v_inst.stateZ0Z_13 ;
    wire \b2v_inst.g2_3 ;
    wire \b2v_inst.borradoZ0 ;
    wire \b2v_inst.stateZ0Z_5 ;
    wire \b2v_inst.g4_0_cascade_ ;
    wire \b2v_inst.g0_0 ;
    wire \b2v_inst.state_ns_a2_0_o2_1_0_2 ;
    wire \b2v_inst.cuenta_RNI4SC81Z0Z_7 ;
    wire \b2v_inst.state_ns_a2_0_o2_0_2 ;
    wire \b2v_inst.stateZ0Z_8 ;
    wire \b2v_inst.dir_mem_2_RNO_0Z0Z_3_cascade_ ;
    wire \b2v_inst.dir_mem_2Z0Z_3 ;
    wire \b2v_inst.un1_dir_mem_3_ns_1_4 ;
    wire \b2v_inst.dir_mem_2_RNO_0Z0Z_7 ;
    wire \b2v_inst.N_237 ;
    wire \b2v_inst.dir_mem_2Z0Z_7 ;
    wire \b2v_inst.N_239 ;
    wire \b2v_inst.addr_ram_1_0_iv_i_1_7_cascade_ ;
    wire \b2v_inst.addr_ram_1_0_iv_i_0_7 ;
    wire N_50;
    wire \b2v_inst.g0_2_6_cascade_ ;
    wire \b2v_inst.g0_2_8 ;
    wire \b2v_inst.i4_mux_cascade_ ;
    wire \b2v_inst.dir_mem_1Z0Z_6 ;
    wire \b2v_inst.un2_dir_mem_3_c5 ;
    wire \b2v_inst.un2_dir_mem_3_ac0_3 ;
    wire \b2v_inst.un2_dir_mem_3_ac0_3_cascade_ ;
    wire \b2v_inst.un1_dir_mem_3_ns_1_5 ;
    wire \b2v_inst.m7_1 ;
    wire \b2v_inst.un8_dir_mem_3_c4_cascade_ ;
    wire \b2v_inst.un8_dir_mem_3_c6 ;
    wire \b2v_inst.un2_indice_1_1_4_cascade_ ;
    wire \b2v_inst.dir_mem_2Z0Z_4 ;
    wire \b2v_inst.dir_mem_2Z0Z_1 ;
    wire \b2v_inst.dir_mem_2Z0Z_2 ;
    wire \b2v_inst.dir_mem_215_0_cascade_ ;
    wire \b2v_inst.dir_mem_2Z0Z_0 ;
    wire \b2v_inst.dir_mem_215_0 ;
    wire \b2v_inst.dir_mem_2Z0Z_5 ;
    wire \b2v_inst.N_136_i ;
    wire \b2v_inst1.N_14 ;
    wire \b2v_inst.dir_mem_RNIGVEE1Z0Z_0 ;
    wire bfn_10_10_0_;
    wire \b2v_inst.dir_mem_RNII5PO1Z0Z_1 ;
    wire \b2v_inst.un2_indice_cry_0 ;
    wire \b2v_inst.dir_mem_RNIL33H1Z0Z_2 ;
    wire \b2v_inst.un2_indice_cry_1 ;
    wire \b2v_inst.dir_mem_RNIN53H1Z0Z_3 ;
    wire \b2v_inst.un2_indice_cry_2 ;
    wire \b2v_inst.un2_indice_cry_3 ;
    wire \b2v_inst.un2_indice_cry_4 ;
    wire \b2v_inst.dir_mem_RNITB3H1Z0Z_6 ;
    wire \b2v_inst.un2_indice_20_6 ;
    wire \b2v_inst.un2_indice_cry_5 ;
    wire \b2v_inst.un2_indice_cry_6 ;
    wire \b2v_inst.un2_indice_21_s0_1_cascade_ ;
    wire \b2v_inst.un2_indice_21_s0_1 ;
    wire \b2v_inst.un2_indice_20_1 ;
    wire \b2v_inst.dir_mem_RNO_2Z0Z_1 ;
    wire \b2v_inst.dir_mem_RNO_3Z0Z_1_cascade_ ;
    wire \b2v_inst.dir_mem_RNIP73H1Z0Z_4 ;
    wire \b2v_inst.dir_mem_RNIR93H1Z0Z_5 ;
    wire \b2v_inst.g1_0_3 ;
    wire \b2v_inst.g0_2_7 ;
    wire \b2v_inst.N_467 ;
    wire \b2v_inst.N_411_cascade_ ;
    wire \b2v_inst.un2_indice_20_5 ;
    wire \b2v_inst.un2_indice_3_iv_0_a2_2_sx_5 ;
    wire \b2v_inst.un2_indice_0_d0_c4_d ;
    wire \b2v_inst.un2_m1_e_0_cascade_ ;
    wire \b2v_inst.dir_mem_RNO_4Z0Z_4_cascade_ ;
    wire \b2v_inst.indice_RNIA33NZ0Z_1 ;
    wire \b2v_inst.N_238 ;
    wire \b2v_inst.N_236 ;
    wire \b2v_inst.dir_mem_3Z0Z_2 ;
    wire \b2v_inst.addr_ram_1_0_iv_i_1_2 ;
    wire \b2v_inst.un10_indice_cascade_ ;
    wire \b2v_inst1.r_RX_Bytece_0_2 ;
    wire \b2v_inst1.r_RX_Byte_1_sqmuxa ;
    wire \b2v_inst1.r_RX_Bytece_0_0_0 ;
    wire \b2v_inst.indice_3_repZ0Z1 ;
    wire \b2v_inst.un2_dir_mem_2_c4_d ;
    wire \b2v_inst1.N_7_cascade_ ;
    wire \b2v_inst1.g0_0_i_a6_1_2 ;
    wire \b2v_inst1.N_9_cascade_ ;
    wire \b2v_inst1.g0_0_i_a6_3_5 ;
    wire \b2v_inst1.N_19_cascade_ ;
    wire \b2v_inst1.N_6 ;
    wire \b2v_inst1.r_SM_Main_1_sqmuxa_1_0 ;
    wire \b2v_inst1.g0_3_4 ;
    wire \b2v_inst1.g0_0_i_a6_2_2_cascade_ ;
    wire \b2v_inst1.g0_0_i_a6_2_1 ;
    wire \b2v_inst1.N_18 ;
    wire \b2v_inst.dir_mem_RNO_2Z0Z_4 ;
    wire \b2v_inst.un2_indice_3_0_i_1_4_cascade_ ;
    wire \b2v_inst.un2_indice_20_4 ;
    wire \b2v_inst.dir_mem_RNO_2Z0Z_7 ;
    wire \b2v_inst.un2_indice_20_7 ;
    wire \b2v_inst.un2_indice_3_0_iv_0_0_7_cascade_ ;
    wire \b2v_inst.un2_indice_21_s0_2 ;
    wire \b2v_inst.un2_indice_20_2 ;
    wire \b2v_inst.un2_indice_21_s1_2 ;
    wire \b2v_inst.un2_indice_3_0_iv_0_1_2_cascade_ ;
    wire \b2v_inst.dir_mem_RNO_3Z0Z_4 ;
    wire \b2v_inst.un2_indice_0_d1_c2 ;
    wire \b2v_inst.N_451 ;
    wire \b2v_inst.un2_indice_21_s0_3 ;
    wire \b2v_inst.un2_indice_20_3 ;
    wire \b2v_inst.un2_indice_21_s1_3 ;
    wire \b2v_inst.un2_indice_3_0_iv_0_0_3_cascade_ ;
    wire \b2v_inst.dir_mem_RNO_5Z0Z_4 ;
    wire \b2v_inst.un2_indice_3_iv_0_1_0_5 ;
    wire \b2v_inst.N_410 ;
    wire \b2v_inst.un2_indice_3_iv_0_0_1 ;
    wire \b2v_inst.N_253_i ;
    wire \b2v_inst.stateZ0Z_17 ;
    wire \b2v_inst.un2_indice_20_0_cascade_ ;
    wire \b2v_inst.N_4_0 ;
    wire \b2v_inst.un2_cuentalto7_3 ;
    wire \b2v_inst.N_228_cascade_ ;
    wire \b2v_inst.cuenta_RNI925FZ0Z_7 ;
    wire \b2v_inst.N_234 ;
    wire \b2v_inst.un2_indice_3_0_iv_0_a2_0_8_2_2 ;
    wire \b2v_inst.N_228 ;
    wire \b2v_inst.N_383_8_cascade_ ;
    wire \b2v_inst.un2_indice_3_0_iv_0_a2_0_8_3_2 ;
    wire \b2v_inst.un10_indice_2_cascade_ ;
    wire \b2v_inst.indice_fast_RNIDAJGZ0Z_2 ;
    wire \b2v_inst.dir_mem_115lto6_1_cascade_ ;
    wire \b2v_inst.un1_dir_mem_1_mb_1_7_cascade_ ;
    wire \b2v_inst.dir_mem_1Z0Z_7 ;
    wire \b2v_inst.indiceZ0Z_4 ;
    wire \b2v_inst.un2_dir_mem_2_c5 ;
    wire \b2v_inst.N_4_0_0_cascade_ ;
    wire \b2v_inst.N_8_0 ;
    wire \b2v_inst.dir_mem_315lto8_a0_1_cascade_ ;
    wire \b2v_inst.indice_fast_RNIRFV61Z0Z_3 ;
    wire \b2v_inst.indice_0_repZ0Z1 ;
    wire \b2v_inst.indice_0_rep1_RNIFJJGZ0 ;
    wire \b2v_inst.indice_1_repZ0Z1 ;
    wire \b2v_inst.indice_fastZ0Z_2 ;
    wire \b2v_inst.dir_mem_215lt6_0_cascade_ ;
    wire \b2v_inst.dir_mem_215lt8 ;
    wire \b2v_inst1.g0_0_i_a6_3_4 ;
    wire \b2v_inst1.r_rx_byteZ0Z_7 ;
    wire \b2v_inst1.r_rx_byteZ0Z_7_cascade_ ;
    wire \b2v_inst1.r_Bit_IndexZ0Z_2 ;
    wire \b2v_inst1.r_Bit_IndexZ0Z_0 ;
    wire \b2v_inst1.r_Bit_IndexZ0Z_1 ;
    wire \b2v_inst1.N_11_0_0 ;
    wire \b2v_inst1.N_9 ;
    wire \b2v_inst1.un1_r_Clk_Count_ac0_1_out_cascade_ ;
    wire \b2v_inst1.m22_ns_1 ;
    wire \b2v_inst1.N_29_mux_cascade_ ;
    wire \b2v_inst1.N_11_cascade_ ;
    wire \b2v_inst1.g0_0_i_1 ;
    wire \b2v_inst1.N_14_0 ;
    wire \b2v_inst1.g0_0_i_0 ;
    wire \b2v_inst1.m6_2_cascade_ ;
    wire \b2v_inst1.N_10_0 ;
    wire \b2v_inst1.g0_7_1 ;
    wire \b2v_inst1.g0_i_1_cascade_ ;
    wire \b2v_inst1.N_11_0 ;
    wire \b2v_inst1.N_32_mux ;
    wire \b2v_inst1.N_10_cascade_ ;
    wire \b2v_inst1.g2_1_cascade_ ;
    wire \b2v_inst1.g2_0 ;
    wire \b2v_inst1.m6_2 ;
    wire \b2v_inst.un2_indice_0_d1_c5 ;
    wire \b2v_inst.dir_memZ0Z_4 ;
    wire \b2v_inst.un2_indice_0_d1_ac0_7_s_0_0 ;
    wire \b2v_inst.dir_memZ0Z_3 ;
    wire \b2v_inst.dir_memZ0Z_5 ;
    wire \b2v_inst.un2_indice_0_d1_ac0_7_s_0_0_cascade_ ;
    wire \b2v_inst.dir_memZ0Z_2 ;
    wire \b2v_inst.dir_memZ0Z_7 ;
    wire \b2v_inst.un2_indice_0_d1_ac0_9_0_cascade_ ;
    wire \b2v_inst.dir_memZ0Z_6 ;
    wire \b2v_inst.un2_indice_21_s1_7 ;
    wire \b2v_inst.state_17_repZ0Z1 ;
    wire \b2v_inst.stateZ0Z_15 ;
    wire reset;
    wire \b2v_inst.N_351_0 ;
    wire CONSTANT_ONE_NET;
    wire \b2v_inst.N_384_cascade_ ;
    wire \b2v_inst.state_17_rep1_RNIN75CZ0Z3 ;
    wire \b2v_inst.un2_indice_3_0_iv_0_0_2 ;
    wire \b2v_inst.dir_memZ0Z_0 ;
    wire \b2v_inst.dir_memZ0Z_1 ;
    wire \b2v_inst.N_253 ;
    wire \b2v_inst.un2_indice_21_s1_1 ;
    wire \b2v_inst.un10_indice_2 ;
    wire \b2v_inst.CO1 ;
    wire \b2v_inst.CO1_cascade_ ;
    wire \b2v_inst.un2_dir_mem_2_c2_cascade_ ;
    wire \b2v_inst.indice_fastZ0Z_0 ;
    wire \b2v_inst.indice_fastZ0Z_1 ;
    wire \b2v_inst.indice_2_repZ0Z1 ;
    wire \b2v_inst.indiceZ0Z_3 ;
    wire \b2v_inst.dir_mem_1_RNO_0Z0Z_3_cascade_ ;
    wire \b2v_inst.dir_mem_1Z0Z_3 ;
    wire \b2v_inst.indice_fast_RNIF91EZ0Z_0 ;
    wire \b2v_inst.dir_mem_115lto8_1 ;
    wire \b2v_inst.dir_mem_115lto6_1 ;
    wire \b2v_inst.un8_dir_mem_1_c7 ;
    wire \b2v_inst.dir_mem_115lto8_1_cascade_ ;
    wire \b2v_inst.dir_mem_115_0_cascade_ ;
    wire \b2v_inst.dir_mem_1Z0Z_0 ;
    wire \b2v_inst.indiceZ0Z_2 ;
    wire \b2v_inst.un2_dir_mem_2_c2 ;
    wire \b2v_inst.dir_mem_1Z0Z_2 ;
    wire \b2v_inst.dir_mem_1_RNO_0Z0Z_5 ;
    wire \b2v_inst.dir_mem_1Z0Z_5 ;
    wire \b2v_inst.dir_mem_115_0 ;
    wire \b2v_inst.dir_mem_1Z0Z_1 ;
    wire \b2v_inst.N_134_i ;
    wire \b2v_inst.un8_dir_mem_3_ac0_9_0_cascade_ ;
    wire \b2v_inst.un10_indice ;
    wire \b2v_inst.indice_4_repZ0Z1 ;
    wire \b2v_inst.indice_1_repZ0Z2 ;
    wire \b2v_inst.indice_0_repZ0Z2 ;
    wire \b2v_inst.un10_indice_2_0 ;
    wire \b2v_inst.un8_dir_mem_3_ac0_9_0 ;
    wire \b2v_inst.indiceZ0Z_7 ;
    wire \b2v_inst.un8_dir_mem_3_c4 ;
    wire \b2v_inst.indice_fastZ0Z_4 ;
    wire \b2v_inst.indice_fastZ0Z_3 ;
    wire \b2v_inst.un8_dir_mem_1_ac0_7_out ;
    wire \b2v_inst.un8_dir_mem_2_c4 ;
    wire \b2v_inst.indiceZ0Z_6 ;
    wire \b2v_inst.indiceZ0Z_5 ;
    wire \b2v_inst.dir_mem_2_RNO_1Z0Z_6 ;
    wire \b2v_inst1.g0_i_o5_0_2 ;
    wire \b2v_inst1.g0_1_4_cascade_ ;
    wire \b2v_inst1.N_28_mux ;
    wire \b2v_inst1.un1_r_SM_Main_3_0 ;
    wire \b2v_inst1.g0_1_cascade_ ;
    wire \b2v_inst1.N_29_mux_1 ;
    wire \b2v_inst1.N_14_0_1_cascade_ ;
    wire \b2v_inst1.g0_0_i_a6_1_5_cascade_ ;
    wire \b2v_inst1.g0_0_i_a6_1_1 ;
    wire \b2v_inst1.un1_r_Clk_Count_ac0_3_out ;
    wire \b2v_inst1.N_29_mux ;
    wire \b2v_inst1.r_SM_Main_1_sqmuxa_1_cascade_ ;
    wire \b2v_inst1.un1_r_SM_Main_1_sqmuxa_0 ;
    wire \b2v_inst1.un1_r_Clk_Count_ac0_1_out ;
    wire \b2v_inst1.r_Clk_CountZ0Z_3 ;
    wire \b2v_inst1.g0_3_1_cascade_ ;
    wire \b2v_inst1.N_14_0_0 ;
    wire \b2v_inst1.N_14_0_0_cascade_ ;
    wire \b2v_inst1.N_29_mux_0 ;
    wire \b2v_inst1.r_Clk_CountZ0Z_0 ;
    wire \b2v_inst1.g3_1_cascade_ ;
    wire \b2v_inst1.r_Clk_CountZ0Z_1 ;
    wire \b2v_inst1.g3 ;
    wire \b2v_inst1.N_9_0 ;
    wire \b2v_inst1.N_13_cascade_ ;
    wire \b2v_inst1.g0_0_i_a6_3_0 ;
    wire \b2v_inst1.g0_0_i_a6_1_6 ;
    wire \b2v_inst1.g0_0_i_1_0_cascade_ ;
    wire \b2v_inst1.N_7_0 ;
    wire \b2v_inst1.r_SM_Main_d_4 ;
    wire \b2v_inst1.r_Clk_CountZ0Z_6 ;
    wire \b2v_inst1.r_Clk_CountZ0Z_5 ;
    wire \b2v_inst1.r_Clk_CountZ0Z_2 ;
    wire \b2v_inst1.g2_1_4 ;
    wire \b2v_inst1.r_SM_MainZ0Z_0 ;
    wire \b2v_inst1.r_SM_MainZ0Z_1 ;
    wire \b2v_inst1.r_SM_MainZ0Z_2 ;
    wire \b2v_inst1.N_11_1 ;
    wire \b2v_inst1.g0_0_i_a6_2_0_cascade_ ;
    wire \b2v_inst1.r_Clk_CountZ0Z_4 ;
    wire \b2v_inst1.g0_0_i_0_0 ;
    wire \b2v_inst.indiceZ0Z_0 ;
    wire \b2v_inst.indiceZ0Z_1 ;
    wire \b2v_inst.state_g_2 ;
    wire reset_i_g;
    wire uart_rx_i;
    wire \b2v_inst1.r_RX_Data_RZ0 ;
    wire \b2v_inst1.r_RX_DataZ0 ;
    wire clk;
    wire _gnd_net_;

    defparam \b2v_inst2.mem_0_mem_0_0_0_physical .WRITE_MODE=0;
    defparam \b2v_inst2.mem_0_mem_0_0_0_physical .READ_MODE=0;
    SB_RAM40_4K \b2v_inst2.mem_0_mem_0_0_0_physical  (
            .RDATA({dangling_wire_0,dangling_wire_1,dangling_wire_2,dangling_wire_3,dangling_wire_4,dangling_wire_5,dangling_wire_6,dangling_wire_7,SYNTHESIZED_WIRE_1_7,SYNTHESIZED_WIRE_1_6,SYNTHESIZED_WIRE_1_5,SYNTHESIZED_WIRE_1_4,SYNTHESIZED_WIRE_1_3,SYNTHESIZED_WIRE_1_2,SYNTHESIZED_WIRE_1_1,SYNTHESIZED_WIRE_1_0}),
            .RADDR({dangling_wire_8,dangling_wire_9,dangling_wire_10,N__16330,N__13937,N__12541,N__15416,N__15107,N__13999,N__14026,N__14059}),
            .WADDR({dangling_wire_11,dangling_wire_12,dangling_wire_13,N__16334,N__13936,N__12542,N__15412,N__15103,N__14000,N__14027,N__14060}),
            .MASK({dangling_wire_14,dangling_wire_15,dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29}),
            .WDATA({dangling_wire_30,dangling_wire_31,dangling_wire_32,dangling_wire_33,dangling_wire_34,dangling_wire_35,dangling_wire_36,dangling_wire_37,N__14126,N__12362,N__12374,N__9047,N__12386,N__9008,N__9020,N__9035}),
            .RCLKE(),
            .RCLK(N__22577),
            .RE(N__18613),
            .WCLKE(N__9992),
            .WCLK(N__22483),
            .WE(N__18620));
    IO_PAD ipInertedIOPad_uart_tx_o_iopad (
            .OE(N__24159),
            .DIN(N__24158),
            .DOUT(N__24157),
            .PACKAGEPIN(uart_tx_o));
    defparam ipInertedIOPad_uart_tx_o_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_uart_tx_o_preio (
            .PADOEN(N__24159),
            .PADOUT(N__24158),
            .PADIN(N__24157),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__11735),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_uart_rx_i_iopad (
            .OE(N__24150),
            .DIN(N__24149),
            .DOUT(N__24148),
            .PACKAGEPIN(uart_rx_i));
    defparam ipInertedIOPad_uart_rx_i_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_uart_rx_i_preio (
            .PADOEN(N__24150),
            .PADOUT(N__24149),
            .PADIN(N__24148),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(uart_rx_i),
            .DIN1());
    IO_PAD ipInertedIOPad_reset_iopad (
            .OE(N__24141),
            .DIN(N__24140),
            .DOUT(N__24139),
            .PACKAGEPIN(reset));
    defparam ipInertedIOPad_reset_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_reset_preio (
            .PADOEN(N__24141),
            .PADOUT(N__24140),
            .PADIN(N__24139),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(reset),
            .DIN1());
    IO_PAD ipInertedIOPad_clk_iopad (
            .OE(N__24132),
            .DIN(N__24131),
            .DOUT(N__24130),
            .PACKAGEPIN(clk));
    defparam ipInertedIOPad_clk_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_clk_preio (
            .PADOEN(N__24132),
            .PADOUT(N__24131),
            .PADIN(N__24130),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(clk),
            .DIN1());
    InMux I__5972 (
            .O(N__24113),
            .I(N__24110));
    LocalMux I__5971 (
            .O(N__24110),
            .I(N__24107));
    Odrv4 I__5970 (
            .O(N__24107),
            .I(\b2v_inst1.g0_0_i_a6_1_6 ));
    CascadeMux I__5969 (
            .O(N__24104),
            .I(\b2v_inst1.g0_0_i_1_0_cascade_ ));
    InMux I__5968 (
            .O(N__24101),
            .I(N__24098));
    LocalMux I__5967 (
            .O(N__24098),
            .I(\b2v_inst1.N_7_0 ));
    SRMux I__5966 (
            .O(N__24095),
            .I(N__24089));
    SRMux I__5965 (
            .O(N__24094),
            .I(N__24086));
    SRMux I__5964 (
            .O(N__24093),
            .I(N__24083));
    SRMux I__5963 (
            .O(N__24092),
            .I(N__24078));
    LocalMux I__5962 (
            .O(N__24089),
            .I(N__24073));
    LocalMux I__5961 (
            .O(N__24086),
            .I(N__24073));
    LocalMux I__5960 (
            .O(N__24083),
            .I(N__24070));
    SRMux I__5959 (
            .O(N__24082),
            .I(N__24067));
    SRMux I__5958 (
            .O(N__24081),
            .I(N__24064));
    LocalMux I__5957 (
            .O(N__24078),
            .I(N__24060));
    Span4Mux_v I__5956 (
            .O(N__24073),
            .I(N__24057));
    Span4Mux_v I__5955 (
            .O(N__24070),
            .I(N__24054));
    LocalMux I__5954 (
            .O(N__24067),
            .I(N__24051));
    LocalMux I__5953 (
            .O(N__24064),
            .I(N__24048));
    SRMux I__5952 (
            .O(N__24063),
            .I(N__24045));
    Span12Mux_s10_v I__5951 (
            .O(N__24060),
            .I(N__24042));
    Sp12to4 I__5950 (
            .O(N__24057),
            .I(N__24037));
    Sp12to4 I__5949 (
            .O(N__24054),
            .I(N__24037));
    Span4Mux_v I__5948 (
            .O(N__24051),
            .I(N__24032));
    Span4Mux_h I__5947 (
            .O(N__24048),
            .I(N__24032));
    LocalMux I__5946 (
            .O(N__24045),
            .I(N__24029));
    Odrv12 I__5945 (
            .O(N__24042),
            .I(\b2v_inst1.r_SM_Main_d_4 ));
    Odrv12 I__5944 (
            .O(N__24037),
            .I(\b2v_inst1.r_SM_Main_d_4 ));
    Odrv4 I__5943 (
            .O(N__24032),
            .I(\b2v_inst1.r_SM_Main_d_4 ));
    Odrv12 I__5942 (
            .O(N__24029),
            .I(\b2v_inst1.r_SM_Main_d_4 ));
    InMux I__5941 (
            .O(N__24020),
            .I(N__24011));
    InMux I__5940 (
            .O(N__24019),
            .I(N__24006));
    InMux I__5939 (
            .O(N__24018),
            .I(N__24006));
    InMux I__5938 (
            .O(N__24017),
            .I(N__23998));
    InMux I__5937 (
            .O(N__24016),
            .I(N__23998));
    InMux I__5936 (
            .O(N__24015),
            .I(N__23993));
    InMux I__5935 (
            .O(N__24014),
            .I(N__23993));
    LocalMux I__5934 (
            .O(N__24011),
            .I(N__23981));
    LocalMux I__5933 (
            .O(N__24006),
            .I(N__23978));
    InMux I__5932 (
            .O(N__24005),
            .I(N__23973));
    InMux I__5931 (
            .O(N__24004),
            .I(N__23973));
    InMux I__5930 (
            .O(N__24003),
            .I(N__23970));
    LocalMux I__5929 (
            .O(N__23998),
            .I(N__23965));
    LocalMux I__5928 (
            .O(N__23993),
            .I(N__23965));
    InMux I__5927 (
            .O(N__23992),
            .I(N__23960));
    InMux I__5926 (
            .O(N__23991),
            .I(N__23960));
    InMux I__5925 (
            .O(N__23990),
            .I(N__23957));
    InMux I__5924 (
            .O(N__23989),
            .I(N__23950));
    InMux I__5923 (
            .O(N__23988),
            .I(N__23950));
    InMux I__5922 (
            .O(N__23987),
            .I(N__23950));
    InMux I__5921 (
            .O(N__23986),
            .I(N__23947));
    InMux I__5920 (
            .O(N__23985),
            .I(N__23942));
    InMux I__5919 (
            .O(N__23984),
            .I(N__23942));
    Odrv4 I__5918 (
            .O(N__23981),
            .I(\b2v_inst1.r_Clk_CountZ0Z_6 ));
    Odrv4 I__5917 (
            .O(N__23978),
            .I(\b2v_inst1.r_Clk_CountZ0Z_6 ));
    LocalMux I__5916 (
            .O(N__23973),
            .I(\b2v_inst1.r_Clk_CountZ0Z_6 ));
    LocalMux I__5915 (
            .O(N__23970),
            .I(\b2v_inst1.r_Clk_CountZ0Z_6 ));
    Odrv4 I__5914 (
            .O(N__23965),
            .I(\b2v_inst1.r_Clk_CountZ0Z_6 ));
    LocalMux I__5913 (
            .O(N__23960),
            .I(\b2v_inst1.r_Clk_CountZ0Z_6 ));
    LocalMux I__5912 (
            .O(N__23957),
            .I(\b2v_inst1.r_Clk_CountZ0Z_6 ));
    LocalMux I__5911 (
            .O(N__23950),
            .I(\b2v_inst1.r_Clk_CountZ0Z_6 ));
    LocalMux I__5910 (
            .O(N__23947),
            .I(\b2v_inst1.r_Clk_CountZ0Z_6 ));
    LocalMux I__5909 (
            .O(N__23942),
            .I(\b2v_inst1.r_Clk_CountZ0Z_6 ));
    InMux I__5908 (
            .O(N__23921),
            .I(N__23905));
    InMux I__5907 (
            .O(N__23920),
            .I(N__23905));
    InMux I__5906 (
            .O(N__23919),
            .I(N__23897));
    InMux I__5905 (
            .O(N__23918),
            .I(N__23894));
    InMux I__5904 (
            .O(N__23917),
            .I(N__23891));
    InMux I__5903 (
            .O(N__23916),
            .I(N__23886));
    InMux I__5902 (
            .O(N__23915),
            .I(N__23886));
    InMux I__5901 (
            .O(N__23914),
            .I(N__23883));
    InMux I__5900 (
            .O(N__23913),
            .I(N__23878));
    InMux I__5899 (
            .O(N__23912),
            .I(N__23878));
    InMux I__5898 (
            .O(N__23911),
            .I(N__23873));
    InMux I__5897 (
            .O(N__23910),
            .I(N__23873));
    LocalMux I__5896 (
            .O(N__23905),
            .I(N__23870));
    InMux I__5895 (
            .O(N__23904),
            .I(N__23863));
    InMux I__5894 (
            .O(N__23903),
            .I(N__23863));
    InMux I__5893 (
            .O(N__23902),
            .I(N__23863));
    InMux I__5892 (
            .O(N__23901),
            .I(N__23858));
    InMux I__5891 (
            .O(N__23900),
            .I(N__23858));
    LocalMux I__5890 (
            .O(N__23897),
            .I(\b2v_inst1.r_Clk_CountZ0Z_5 ));
    LocalMux I__5889 (
            .O(N__23894),
            .I(\b2v_inst1.r_Clk_CountZ0Z_5 ));
    LocalMux I__5888 (
            .O(N__23891),
            .I(\b2v_inst1.r_Clk_CountZ0Z_5 ));
    LocalMux I__5887 (
            .O(N__23886),
            .I(\b2v_inst1.r_Clk_CountZ0Z_5 ));
    LocalMux I__5886 (
            .O(N__23883),
            .I(\b2v_inst1.r_Clk_CountZ0Z_5 ));
    LocalMux I__5885 (
            .O(N__23878),
            .I(\b2v_inst1.r_Clk_CountZ0Z_5 ));
    LocalMux I__5884 (
            .O(N__23873),
            .I(\b2v_inst1.r_Clk_CountZ0Z_5 ));
    Odrv4 I__5883 (
            .O(N__23870),
            .I(\b2v_inst1.r_Clk_CountZ0Z_5 ));
    LocalMux I__5882 (
            .O(N__23863),
            .I(\b2v_inst1.r_Clk_CountZ0Z_5 ));
    LocalMux I__5881 (
            .O(N__23858),
            .I(\b2v_inst1.r_Clk_CountZ0Z_5 ));
    InMux I__5880 (
            .O(N__23837),
            .I(N__23824));
    InMux I__5879 (
            .O(N__23836),
            .I(N__23824));
    InMux I__5878 (
            .O(N__23835),
            .I(N__23815));
    InMux I__5877 (
            .O(N__23834),
            .I(N__23815));
    InMux I__5876 (
            .O(N__23833),
            .I(N__23810));
    InMux I__5875 (
            .O(N__23832),
            .I(N__23810));
    InMux I__5874 (
            .O(N__23831),
            .I(N__23804));
    InMux I__5873 (
            .O(N__23830),
            .I(N__23804));
    InMux I__5872 (
            .O(N__23829),
            .I(N__23801));
    LocalMux I__5871 (
            .O(N__23824),
            .I(N__23798));
    InMux I__5870 (
            .O(N__23823),
            .I(N__23793));
    InMux I__5869 (
            .O(N__23822),
            .I(N__23793));
    InMux I__5868 (
            .O(N__23821),
            .I(N__23790));
    InMux I__5867 (
            .O(N__23820),
            .I(N__23787));
    LocalMux I__5866 (
            .O(N__23815),
            .I(N__23782));
    LocalMux I__5865 (
            .O(N__23810),
            .I(N__23782));
    InMux I__5864 (
            .O(N__23809),
            .I(N__23779));
    LocalMux I__5863 (
            .O(N__23804),
            .I(\b2v_inst1.r_Clk_CountZ0Z_2 ));
    LocalMux I__5862 (
            .O(N__23801),
            .I(\b2v_inst1.r_Clk_CountZ0Z_2 ));
    Odrv4 I__5861 (
            .O(N__23798),
            .I(\b2v_inst1.r_Clk_CountZ0Z_2 ));
    LocalMux I__5860 (
            .O(N__23793),
            .I(\b2v_inst1.r_Clk_CountZ0Z_2 ));
    LocalMux I__5859 (
            .O(N__23790),
            .I(\b2v_inst1.r_Clk_CountZ0Z_2 ));
    LocalMux I__5858 (
            .O(N__23787),
            .I(\b2v_inst1.r_Clk_CountZ0Z_2 ));
    Odrv4 I__5857 (
            .O(N__23782),
            .I(\b2v_inst1.r_Clk_CountZ0Z_2 ));
    LocalMux I__5856 (
            .O(N__23779),
            .I(\b2v_inst1.r_Clk_CountZ0Z_2 ));
    InMux I__5855 (
            .O(N__23762),
            .I(N__23759));
    LocalMux I__5854 (
            .O(N__23759),
            .I(\b2v_inst1.g2_1_4 ));
    CascadeMux I__5853 (
            .O(N__23756),
            .I(N__23750));
    InMux I__5852 (
            .O(N__23755),
            .I(N__23743));
    InMux I__5851 (
            .O(N__23754),
            .I(N__23743));
    InMux I__5850 (
            .O(N__23753),
            .I(N__23735));
    InMux I__5849 (
            .O(N__23750),
            .I(N__23730));
    InMux I__5848 (
            .O(N__23749),
            .I(N__23730));
    CascadeMux I__5847 (
            .O(N__23748),
            .I(N__23724));
    LocalMux I__5846 (
            .O(N__23743),
            .I(N__23721));
    CascadeMux I__5845 (
            .O(N__23742),
            .I(N__23718));
    InMux I__5844 (
            .O(N__23741),
            .I(N__23715));
    InMux I__5843 (
            .O(N__23740),
            .I(N__23712));
    InMux I__5842 (
            .O(N__23739),
            .I(N__23709));
    InMux I__5841 (
            .O(N__23738),
            .I(N__23700));
    LocalMux I__5840 (
            .O(N__23735),
            .I(N__23695));
    LocalMux I__5839 (
            .O(N__23730),
            .I(N__23695));
    InMux I__5838 (
            .O(N__23729),
            .I(N__23690));
    InMux I__5837 (
            .O(N__23728),
            .I(N__23690));
    InMux I__5836 (
            .O(N__23727),
            .I(N__23685));
    InMux I__5835 (
            .O(N__23724),
            .I(N__23685));
    Span4Mux_h I__5834 (
            .O(N__23721),
            .I(N__23682));
    InMux I__5833 (
            .O(N__23718),
            .I(N__23679));
    LocalMux I__5832 (
            .O(N__23715),
            .I(N__23672));
    LocalMux I__5831 (
            .O(N__23712),
            .I(N__23672));
    LocalMux I__5830 (
            .O(N__23709),
            .I(N__23672));
    InMux I__5829 (
            .O(N__23708),
            .I(N__23667));
    InMux I__5828 (
            .O(N__23707),
            .I(N__23667));
    InMux I__5827 (
            .O(N__23706),
            .I(N__23664));
    InMux I__5826 (
            .O(N__23705),
            .I(N__23661));
    InMux I__5825 (
            .O(N__23704),
            .I(N__23656));
    InMux I__5824 (
            .O(N__23703),
            .I(N__23656));
    LocalMux I__5823 (
            .O(N__23700),
            .I(N__23647));
    Span4Mux_h I__5822 (
            .O(N__23695),
            .I(N__23647));
    LocalMux I__5821 (
            .O(N__23690),
            .I(N__23647));
    LocalMux I__5820 (
            .O(N__23685),
            .I(N__23647));
    Odrv4 I__5819 (
            .O(N__23682),
            .I(\b2v_inst1.r_SM_MainZ0Z_0 ));
    LocalMux I__5818 (
            .O(N__23679),
            .I(\b2v_inst1.r_SM_MainZ0Z_0 ));
    Odrv4 I__5817 (
            .O(N__23672),
            .I(\b2v_inst1.r_SM_MainZ0Z_0 ));
    LocalMux I__5816 (
            .O(N__23667),
            .I(\b2v_inst1.r_SM_MainZ0Z_0 ));
    LocalMux I__5815 (
            .O(N__23664),
            .I(\b2v_inst1.r_SM_MainZ0Z_0 ));
    LocalMux I__5814 (
            .O(N__23661),
            .I(\b2v_inst1.r_SM_MainZ0Z_0 ));
    LocalMux I__5813 (
            .O(N__23656),
            .I(\b2v_inst1.r_SM_MainZ0Z_0 ));
    Odrv4 I__5812 (
            .O(N__23647),
            .I(\b2v_inst1.r_SM_MainZ0Z_0 ));
    InMux I__5811 (
            .O(N__23630),
            .I(N__23626));
    InMux I__5810 (
            .O(N__23629),
            .I(N__23614));
    LocalMux I__5809 (
            .O(N__23626),
            .I(N__23609));
    CascadeMux I__5808 (
            .O(N__23625),
            .I(N__23604));
    InMux I__5807 (
            .O(N__23624),
            .I(N__23600));
    CascadeMux I__5806 (
            .O(N__23623),
            .I(N__23595));
    InMux I__5805 (
            .O(N__23622),
            .I(N__23583));
    InMux I__5804 (
            .O(N__23621),
            .I(N__23583));
    InMux I__5803 (
            .O(N__23620),
            .I(N__23574));
    InMux I__5802 (
            .O(N__23619),
            .I(N__23574));
    InMux I__5801 (
            .O(N__23618),
            .I(N__23574));
    InMux I__5800 (
            .O(N__23617),
            .I(N__23574));
    LocalMux I__5799 (
            .O(N__23614),
            .I(N__23571));
    InMux I__5798 (
            .O(N__23613),
            .I(N__23566));
    InMux I__5797 (
            .O(N__23612),
            .I(N__23566));
    Span4Mux_v I__5796 (
            .O(N__23609),
            .I(N__23563));
    InMux I__5795 (
            .O(N__23608),
            .I(N__23558));
    InMux I__5794 (
            .O(N__23607),
            .I(N__23558));
    InMux I__5793 (
            .O(N__23604),
            .I(N__23553));
    InMux I__5792 (
            .O(N__23603),
            .I(N__23553));
    LocalMux I__5791 (
            .O(N__23600),
            .I(N__23550));
    InMux I__5790 (
            .O(N__23599),
            .I(N__23545));
    InMux I__5789 (
            .O(N__23598),
            .I(N__23545));
    InMux I__5788 (
            .O(N__23595),
            .I(N__23540));
    InMux I__5787 (
            .O(N__23594),
            .I(N__23540));
    InMux I__5786 (
            .O(N__23593),
            .I(N__23533));
    InMux I__5785 (
            .O(N__23592),
            .I(N__23533));
    InMux I__5784 (
            .O(N__23591),
            .I(N__23533));
    InMux I__5783 (
            .O(N__23590),
            .I(N__23526));
    InMux I__5782 (
            .O(N__23589),
            .I(N__23526));
    InMux I__5781 (
            .O(N__23588),
            .I(N__23526));
    LocalMux I__5780 (
            .O(N__23583),
            .I(N__23519));
    LocalMux I__5779 (
            .O(N__23574),
            .I(N__23519));
    Span4Mux_h I__5778 (
            .O(N__23571),
            .I(N__23519));
    LocalMux I__5777 (
            .O(N__23566),
            .I(\b2v_inst1.r_SM_MainZ0Z_1 ));
    Odrv4 I__5776 (
            .O(N__23563),
            .I(\b2v_inst1.r_SM_MainZ0Z_1 ));
    LocalMux I__5775 (
            .O(N__23558),
            .I(\b2v_inst1.r_SM_MainZ0Z_1 ));
    LocalMux I__5774 (
            .O(N__23553),
            .I(\b2v_inst1.r_SM_MainZ0Z_1 ));
    Odrv4 I__5773 (
            .O(N__23550),
            .I(\b2v_inst1.r_SM_MainZ0Z_1 ));
    LocalMux I__5772 (
            .O(N__23545),
            .I(\b2v_inst1.r_SM_MainZ0Z_1 ));
    LocalMux I__5771 (
            .O(N__23540),
            .I(\b2v_inst1.r_SM_MainZ0Z_1 ));
    LocalMux I__5770 (
            .O(N__23533),
            .I(\b2v_inst1.r_SM_MainZ0Z_1 ));
    LocalMux I__5769 (
            .O(N__23526),
            .I(\b2v_inst1.r_SM_MainZ0Z_1 ));
    Odrv4 I__5768 (
            .O(N__23519),
            .I(\b2v_inst1.r_SM_MainZ0Z_1 ));
    CascadeMux I__5767 (
            .O(N__23498),
            .I(N__23491));
    InMux I__5766 (
            .O(N__23497),
            .I(N__23485));
    CascadeMux I__5765 (
            .O(N__23496),
            .I(N__23479));
    CascadeMux I__5764 (
            .O(N__23495),
            .I(N__23476));
    InMux I__5763 (
            .O(N__23494),
            .I(N__23471));
    InMux I__5762 (
            .O(N__23491),
            .I(N__23468));
    InMux I__5761 (
            .O(N__23490),
            .I(N__23465));
    InMux I__5760 (
            .O(N__23489),
            .I(N__23462));
    InMux I__5759 (
            .O(N__23488),
            .I(N__23459));
    LocalMux I__5758 (
            .O(N__23485),
            .I(N__23456));
    CascadeMux I__5757 (
            .O(N__23484),
            .I(N__23452));
    InMux I__5756 (
            .O(N__23483),
            .I(N__23449));
    InMux I__5755 (
            .O(N__23482),
            .I(N__23446));
    InMux I__5754 (
            .O(N__23479),
            .I(N__23442));
    InMux I__5753 (
            .O(N__23476),
            .I(N__23439));
    CascadeMux I__5752 (
            .O(N__23475),
            .I(N__23436));
    CascadeMux I__5751 (
            .O(N__23474),
            .I(N__23433));
    LocalMux I__5750 (
            .O(N__23471),
            .I(N__23430));
    LocalMux I__5749 (
            .O(N__23468),
            .I(N__23427));
    LocalMux I__5748 (
            .O(N__23465),
            .I(N__23420));
    LocalMux I__5747 (
            .O(N__23462),
            .I(N__23420));
    LocalMux I__5746 (
            .O(N__23459),
            .I(N__23420));
    Span4Mux_v I__5745 (
            .O(N__23456),
            .I(N__23417));
    InMux I__5744 (
            .O(N__23455),
            .I(N__23412));
    InMux I__5743 (
            .O(N__23452),
            .I(N__23412));
    LocalMux I__5742 (
            .O(N__23449),
            .I(N__23409));
    LocalMux I__5741 (
            .O(N__23446),
            .I(N__23406));
    InMux I__5740 (
            .O(N__23445),
            .I(N__23403));
    LocalMux I__5739 (
            .O(N__23442),
            .I(N__23398));
    LocalMux I__5738 (
            .O(N__23439),
            .I(N__23398));
    InMux I__5737 (
            .O(N__23436),
            .I(N__23395));
    InMux I__5736 (
            .O(N__23433),
            .I(N__23392));
    Span4Mux_v I__5735 (
            .O(N__23430),
            .I(N__23379));
    Span4Mux_v I__5734 (
            .O(N__23427),
            .I(N__23379));
    Span4Mux_v I__5733 (
            .O(N__23420),
            .I(N__23379));
    Span4Mux_h I__5732 (
            .O(N__23417),
            .I(N__23379));
    LocalMux I__5731 (
            .O(N__23412),
            .I(N__23379));
    Span4Mux_v I__5730 (
            .O(N__23409),
            .I(N__23379));
    Odrv4 I__5729 (
            .O(N__23406),
            .I(\b2v_inst1.r_SM_MainZ0Z_2 ));
    LocalMux I__5728 (
            .O(N__23403),
            .I(\b2v_inst1.r_SM_MainZ0Z_2 ));
    Odrv4 I__5727 (
            .O(N__23398),
            .I(\b2v_inst1.r_SM_MainZ0Z_2 ));
    LocalMux I__5726 (
            .O(N__23395),
            .I(\b2v_inst1.r_SM_MainZ0Z_2 ));
    LocalMux I__5725 (
            .O(N__23392),
            .I(\b2v_inst1.r_SM_MainZ0Z_2 ));
    Odrv4 I__5724 (
            .O(N__23379),
            .I(\b2v_inst1.r_SM_MainZ0Z_2 ));
    InMux I__5723 (
            .O(N__23366),
            .I(N__23362));
    InMux I__5722 (
            .O(N__23365),
            .I(N__23359));
    LocalMux I__5721 (
            .O(N__23362),
            .I(\b2v_inst1.N_11_1 ));
    LocalMux I__5720 (
            .O(N__23359),
            .I(\b2v_inst1.N_11_1 ));
    CascadeMux I__5719 (
            .O(N__23354),
            .I(\b2v_inst1.g0_0_i_a6_2_0_cascade_ ));
    CascadeMux I__5718 (
            .O(N__23351),
            .I(N__23348));
    InMux I__5717 (
            .O(N__23348),
            .I(N__23336));
    InMux I__5716 (
            .O(N__23347),
            .I(N__23336));
    CascadeMux I__5715 (
            .O(N__23346),
            .I(N__23333));
    CascadeMux I__5714 (
            .O(N__23345),
            .I(N__23330));
    CascadeMux I__5713 (
            .O(N__23344),
            .I(N__23327));
    InMux I__5712 (
            .O(N__23343),
            .I(N__23324));
    InMux I__5711 (
            .O(N__23342),
            .I(N__23321));
    CascadeMux I__5710 (
            .O(N__23341),
            .I(N__23317));
    LocalMux I__5709 (
            .O(N__23336),
            .I(N__23310));
    InMux I__5708 (
            .O(N__23333),
            .I(N__23305));
    InMux I__5707 (
            .O(N__23330),
            .I(N__23305));
    InMux I__5706 (
            .O(N__23327),
            .I(N__23302));
    LocalMux I__5705 (
            .O(N__23324),
            .I(N__23296));
    LocalMux I__5704 (
            .O(N__23321),
            .I(N__23296));
    CascadeMux I__5703 (
            .O(N__23320),
            .I(N__23291));
    InMux I__5702 (
            .O(N__23317),
            .I(N__23286));
    InMux I__5701 (
            .O(N__23316),
            .I(N__23286));
    InMux I__5700 (
            .O(N__23315),
            .I(N__23282));
    InMux I__5699 (
            .O(N__23314),
            .I(N__23279));
    InMux I__5698 (
            .O(N__23313),
            .I(N__23276));
    Span4Mux_v I__5697 (
            .O(N__23310),
            .I(N__23271));
    LocalMux I__5696 (
            .O(N__23305),
            .I(N__23271));
    LocalMux I__5695 (
            .O(N__23302),
            .I(N__23268));
    InMux I__5694 (
            .O(N__23301),
            .I(N__23265));
    Span4Mux_h I__5693 (
            .O(N__23296),
            .I(N__23262));
    InMux I__5692 (
            .O(N__23295),
            .I(N__23255));
    InMux I__5691 (
            .O(N__23294),
            .I(N__23255));
    InMux I__5690 (
            .O(N__23291),
            .I(N__23255));
    LocalMux I__5689 (
            .O(N__23286),
            .I(N__23252));
    InMux I__5688 (
            .O(N__23285),
            .I(N__23249));
    LocalMux I__5687 (
            .O(N__23282),
            .I(N__23238));
    LocalMux I__5686 (
            .O(N__23279),
            .I(N__23238));
    LocalMux I__5685 (
            .O(N__23276),
            .I(N__23238));
    Span4Mux_h I__5684 (
            .O(N__23271),
            .I(N__23238));
    Span4Mux_h I__5683 (
            .O(N__23268),
            .I(N__23238));
    LocalMux I__5682 (
            .O(N__23265),
            .I(\b2v_inst1.r_Clk_CountZ0Z_4 ));
    Odrv4 I__5681 (
            .O(N__23262),
            .I(\b2v_inst1.r_Clk_CountZ0Z_4 ));
    LocalMux I__5680 (
            .O(N__23255),
            .I(\b2v_inst1.r_Clk_CountZ0Z_4 ));
    Odrv4 I__5679 (
            .O(N__23252),
            .I(\b2v_inst1.r_Clk_CountZ0Z_4 ));
    LocalMux I__5678 (
            .O(N__23249),
            .I(\b2v_inst1.r_Clk_CountZ0Z_4 ));
    Odrv4 I__5677 (
            .O(N__23238),
            .I(\b2v_inst1.r_Clk_CountZ0Z_4 ));
    InMux I__5676 (
            .O(N__23225),
            .I(N__23222));
    LocalMux I__5675 (
            .O(N__23222),
            .I(\b2v_inst1.g0_0_i_0_0 ));
    CascadeMux I__5674 (
            .O(N__23219),
            .I(N__23212));
    InMux I__5673 (
            .O(N__23218),
            .I(N__23207));
    CascadeMux I__5672 (
            .O(N__23217),
            .I(N__23203));
    CascadeMux I__5671 (
            .O(N__23216),
            .I(N__23196));
    CascadeMux I__5670 (
            .O(N__23215),
            .I(N__23192));
    InMux I__5669 (
            .O(N__23212),
            .I(N__23185));
    InMux I__5668 (
            .O(N__23211),
            .I(N__23185));
    InMux I__5667 (
            .O(N__23210),
            .I(N__23185));
    LocalMux I__5666 (
            .O(N__23207),
            .I(N__23182));
    InMux I__5665 (
            .O(N__23206),
            .I(N__23177));
    InMux I__5664 (
            .O(N__23203),
            .I(N__23177));
    InMux I__5663 (
            .O(N__23202),
            .I(N__23168));
    InMux I__5662 (
            .O(N__23201),
            .I(N__23168));
    InMux I__5661 (
            .O(N__23200),
            .I(N__23163));
    InMux I__5660 (
            .O(N__23199),
            .I(N__23158));
    InMux I__5659 (
            .O(N__23196),
            .I(N__23158));
    InMux I__5658 (
            .O(N__23195),
            .I(N__23153));
    InMux I__5657 (
            .O(N__23192),
            .I(N__23153));
    LocalMux I__5656 (
            .O(N__23185),
            .I(N__23149));
    Span4Mux_v I__5655 (
            .O(N__23182),
            .I(N__23144));
    LocalMux I__5654 (
            .O(N__23177),
            .I(N__23144));
    InMux I__5653 (
            .O(N__23176),
            .I(N__23135));
    InMux I__5652 (
            .O(N__23175),
            .I(N__23135));
    InMux I__5651 (
            .O(N__23174),
            .I(N__23135));
    InMux I__5650 (
            .O(N__23173),
            .I(N__23135));
    LocalMux I__5649 (
            .O(N__23168),
            .I(N__23131));
    InMux I__5648 (
            .O(N__23167),
            .I(N__23126));
    InMux I__5647 (
            .O(N__23166),
            .I(N__23126));
    LocalMux I__5646 (
            .O(N__23163),
            .I(N__23119));
    LocalMux I__5645 (
            .O(N__23158),
            .I(N__23119));
    LocalMux I__5644 (
            .O(N__23153),
            .I(N__23119));
    InMux I__5643 (
            .O(N__23152),
            .I(N__23116));
    Span12Mux_v I__5642 (
            .O(N__23149),
            .I(N__23113));
    Span4Mux_h I__5641 (
            .O(N__23144),
            .I(N__23110));
    LocalMux I__5640 (
            .O(N__23135),
            .I(N__23107));
    InMux I__5639 (
            .O(N__23134),
            .I(N__23104));
    Span4Mux_v I__5638 (
            .O(N__23131),
            .I(N__23097));
    LocalMux I__5637 (
            .O(N__23126),
            .I(N__23097));
    Span4Mux_h I__5636 (
            .O(N__23119),
            .I(N__23097));
    LocalMux I__5635 (
            .O(N__23116),
            .I(\b2v_inst.indiceZ0Z_0 ));
    Odrv12 I__5634 (
            .O(N__23113),
            .I(\b2v_inst.indiceZ0Z_0 ));
    Odrv4 I__5633 (
            .O(N__23110),
            .I(\b2v_inst.indiceZ0Z_0 ));
    Odrv12 I__5632 (
            .O(N__23107),
            .I(\b2v_inst.indiceZ0Z_0 ));
    LocalMux I__5631 (
            .O(N__23104),
            .I(\b2v_inst.indiceZ0Z_0 ));
    Odrv4 I__5630 (
            .O(N__23097),
            .I(\b2v_inst.indiceZ0Z_0 ));
    InMux I__5629 (
            .O(N__23084),
            .I(N__23078));
    InMux I__5628 (
            .O(N__23083),
            .I(N__23071));
    InMux I__5627 (
            .O(N__23082),
            .I(N__23071));
    InMux I__5626 (
            .O(N__23081),
            .I(N__23068));
    LocalMux I__5625 (
            .O(N__23078),
            .I(N__23065));
    CascadeMux I__5624 (
            .O(N__23077),
            .I(N__23060));
    CascadeMux I__5623 (
            .O(N__23076),
            .I(N__23055));
    LocalMux I__5622 (
            .O(N__23071),
            .I(N__23051));
    LocalMux I__5621 (
            .O(N__23068),
            .I(N__23048));
    Span4Mux_v I__5620 (
            .O(N__23065),
            .I(N__23045));
    InMux I__5619 (
            .O(N__23064),
            .I(N__23038));
    InMux I__5618 (
            .O(N__23063),
            .I(N__23038));
    InMux I__5617 (
            .O(N__23060),
            .I(N__23038));
    InMux I__5616 (
            .O(N__23059),
            .I(N__23029));
    InMux I__5615 (
            .O(N__23058),
            .I(N__23029));
    InMux I__5614 (
            .O(N__23055),
            .I(N__23029));
    CascadeMux I__5613 (
            .O(N__23054),
            .I(N__23024));
    Span4Mux_v I__5612 (
            .O(N__23051),
            .I(N__23012));
    Span4Mux_h I__5611 (
            .O(N__23048),
            .I(N__23012));
    Span4Mux_v I__5610 (
            .O(N__23045),
            .I(N__23012));
    LocalMux I__5609 (
            .O(N__23038),
            .I(N__23012));
    InMux I__5608 (
            .O(N__23037),
            .I(N__23007));
    InMux I__5607 (
            .O(N__23036),
            .I(N__23007));
    LocalMux I__5606 (
            .O(N__23029),
            .I(N__23004));
    InMux I__5605 (
            .O(N__23028),
            .I(N__22997));
    InMux I__5604 (
            .O(N__23027),
            .I(N__22997));
    InMux I__5603 (
            .O(N__23024),
            .I(N__22997));
    InMux I__5602 (
            .O(N__23023),
            .I(N__22991));
    InMux I__5601 (
            .O(N__23022),
            .I(N__22991));
    InMux I__5600 (
            .O(N__23021),
            .I(N__22988));
    Span4Mux_h I__5599 (
            .O(N__23012),
            .I(N__22985));
    LocalMux I__5598 (
            .O(N__23007),
            .I(N__22982));
    Span4Mux_v I__5597 (
            .O(N__23004),
            .I(N__22977));
    LocalMux I__5596 (
            .O(N__22997),
            .I(N__22977));
    InMux I__5595 (
            .O(N__22996),
            .I(N__22974));
    LocalMux I__5594 (
            .O(N__22991),
            .I(N__22969));
    LocalMux I__5593 (
            .O(N__22988),
            .I(N__22969));
    Span4Mux_h I__5592 (
            .O(N__22985),
            .I(N__22966));
    Span4Mux_v I__5591 (
            .O(N__22982),
            .I(N__22961));
    Span4Mux_h I__5590 (
            .O(N__22977),
            .I(N__22961));
    LocalMux I__5589 (
            .O(N__22974),
            .I(\b2v_inst.indiceZ0Z_1 ));
    Odrv4 I__5588 (
            .O(N__22969),
            .I(\b2v_inst.indiceZ0Z_1 ));
    Odrv4 I__5587 (
            .O(N__22966),
            .I(\b2v_inst.indiceZ0Z_1 ));
    Odrv4 I__5586 (
            .O(N__22961),
            .I(\b2v_inst.indiceZ0Z_1 ));
    CEMux I__5585 (
            .O(N__22952),
            .I(N__22928));
    CEMux I__5584 (
            .O(N__22951),
            .I(N__22928));
    CEMux I__5583 (
            .O(N__22950),
            .I(N__22928));
    CEMux I__5582 (
            .O(N__22949),
            .I(N__22928));
    CEMux I__5581 (
            .O(N__22948),
            .I(N__22928));
    CEMux I__5580 (
            .O(N__22947),
            .I(N__22928));
    CEMux I__5579 (
            .O(N__22946),
            .I(N__22928));
    CEMux I__5578 (
            .O(N__22945),
            .I(N__22928));
    GlobalMux I__5577 (
            .O(N__22928),
            .I(N__22925));
    gio2CtrlBuf I__5576 (
            .O(N__22925),
            .I(\b2v_inst.state_g_2 ));
    SRMux I__5575 (
            .O(N__22922),
            .I(N__22778));
    SRMux I__5574 (
            .O(N__22921),
            .I(N__22778));
    SRMux I__5573 (
            .O(N__22920),
            .I(N__22778));
    SRMux I__5572 (
            .O(N__22919),
            .I(N__22778));
    SRMux I__5571 (
            .O(N__22918),
            .I(N__22778));
    SRMux I__5570 (
            .O(N__22917),
            .I(N__22778));
    SRMux I__5569 (
            .O(N__22916),
            .I(N__22778));
    SRMux I__5568 (
            .O(N__22915),
            .I(N__22778));
    SRMux I__5567 (
            .O(N__22914),
            .I(N__22778));
    SRMux I__5566 (
            .O(N__22913),
            .I(N__22778));
    SRMux I__5565 (
            .O(N__22912),
            .I(N__22778));
    SRMux I__5564 (
            .O(N__22911),
            .I(N__22778));
    SRMux I__5563 (
            .O(N__22910),
            .I(N__22778));
    SRMux I__5562 (
            .O(N__22909),
            .I(N__22778));
    SRMux I__5561 (
            .O(N__22908),
            .I(N__22778));
    SRMux I__5560 (
            .O(N__22907),
            .I(N__22778));
    SRMux I__5559 (
            .O(N__22906),
            .I(N__22778));
    SRMux I__5558 (
            .O(N__22905),
            .I(N__22778));
    SRMux I__5557 (
            .O(N__22904),
            .I(N__22778));
    SRMux I__5556 (
            .O(N__22903),
            .I(N__22778));
    SRMux I__5555 (
            .O(N__22902),
            .I(N__22778));
    SRMux I__5554 (
            .O(N__22901),
            .I(N__22778));
    SRMux I__5553 (
            .O(N__22900),
            .I(N__22778));
    SRMux I__5552 (
            .O(N__22899),
            .I(N__22778));
    SRMux I__5551 (
            .O(N__22898),
            .I(N__22778));
    SRMux I__5550 (
            .O(N__22897),
            .I(N__22778));
    SRMux I__5549 (
            .O(N__22896),
            .I(N__22778));
    SRMux I__5548 (
            .O(N__22895),
            .I(N__22778));
    SRMux I__5547 (
            .O(N__22894),
            .I(N__22778));
    SRMux I__5546 (
            .O(N__22893),
            .I(N__22778));
    SRMux I__5545 (
            .O(N__22892),
            .I(N__22778));
    SRMux I__5544 (
            .O(N__22891),
            .I(N__22778));
    SRMux I__5543 (
            .O(N__22890),
            .I(N__22778));
    SRMux I__5542 (
            .O(N__22889),
            .I(N__22778));
    SRMux I__5541 (
            .O(N__22888),
            .I(N__22778));
    SRMux I__5540 (
            .O(N__22887),
            .I(N__22778));
    SRMux I__5539 (
            .O(N__22886),
            .I(N__22778));
    SRMux I__5538 (
            .O(N__22885),
            .I(N__22778));
    SRMux I__5537 (
            .O(N__22884),
            .I(N__22778));
    SRMux I__5536 (
            .O(N__22883),
            .I(N__22778));
    SRMux I__5535 (
            .O(N__22882),
            .I(N__22778));
    SRMux I__5534 (
            .O(N__22881),
            .I(N__22778));
    SRMux I__5533 (
            .O(N__22880),
            .I(N__22778));
    SRMux I__5532 (
            .O(N__22879),
            .I(N__22778));
    SRMux I__5531 (
            .O(N__22878),
            .I(N__22778));
    SRMux I__5530 (
            .O(N__22877),
            .I(N__22778));
    SRMux I__5529 (
            .O(N__22876),
            .I(N__22778));
    SRMux I__5528 (
            .O(N__22875),
            .I(N__22778));
    GlobalMux I__5527 (
            .O(N__22778),
            .I(N__22775));
    gio2CtrlBuf I__5526 (
            .O(N__22775),
            .I(reset_i_g));
    InMux I__5525 (
            .O(N__22772),
            .I(N__22769));
    LocalMux I__5524 (
            .O(N__22769),
            .I(N__22766));
    Span4Mux_h I__5523 (
            .O(N__22766),
            .I(N__22763));
    Span4Mux_v I__5522 (
            .O(N__22763),
            .I(N__22760));
    Odrv4 I__5521 (
            .O(N__22760),
            .I(uart_rx_i));
    InMux I__5520 (
            .O(N__22757),
            .I(N__22754));
    LocalMux I__5519 (
            .O(N__22754),
            .I(\b2v_inst1.r_RX_Data_RZ0 ));
    CascadeMux I__5518 (
            .O(N__22751),
            .I(N__22743));
    CascadeMux I__5517 (
            .O(N__22750),
            .I(N__22740));
    CascadeMux I__5516 (
            .O(N__22749),
            .I(N__22737));
    CascadeMux I__5515 (
            .O(N__22748),
            .I(N__22734));
    CascadeMux I__5514 (
            .O(N__22747),
            .I(N__22730));
    CascadeMux I__5513 (
            .O(N__22746),
            .I(N__22727));
    InMux I__5512 (
            .O(N__22743),
            .I(N__22724));
    InMux I__5511 (
            .O(N__22740),
            .I(N__22715));
    InMux I__5510 (
            .O(N__22737),
            .I(N__22715));
    InMux I__5509 (
            .O(N__22734),
            .I(N__22715));
    InMux I__5508 (
            .O(N__22733),
            .I(N__22715));
    InMux I__5507 (
            .O(N__22730),
            .I(N__22710));
    InMux I__5506 (
            .O(N__22727),
            .I(N__22710));
    LocalMux I__5505 (
            .O(N__22724),
            .I(N__22705));
    LocalMux I__5504 (
            .O(N__22715),
            .I(N__22700));
    LocalMux I__5503 (
            .O(N__22710),
            .I(N__22700));
    CascadeMux I__5502 (
            .O(N__22709),
            .I(N__22695));
    InMux I__5501 (
            .O(N__22708),
            .I(N__22691));
    Span4Mux_h I__5500 (
            .O(N__22705),
            .I(N__22686));
    Span4Mux_v I__5499 (
            .O(N__22700),
            .I(N__22683));
    CascadeMux I__5498 (
            .O(N__22699),
            .I(N__22680));
    CascadeMux I__5497 (
            .O(N__22698),
            .I(N__22676));
    InMux I__5496 (
            .O(N__22695),
            .I(N__22673));
    InMux I__5495 (
            .O(N__22694),
            .I(N__22670));
    LocalMux I__5494 (
            .O(N__22691),
            .I(N__22667));
    InMux I__5493 (
            .O(N__22690),
            .I(N__22664));
    CascadeMux I__5492 (
            .O(N__22689),
            .I(N__22661));
    Span4Mux_h I__5491 (
            .O(N__22686),
            .I(N__22658));
    Span4Mux_v I__5490 (
            .O(N__22683),
            .I(N__22655));
    InMux I__5489 (
            .O(N__22680),
            .I(N__22650));
    InMux I__5488 (
            .O(N__22679),
            .I(N__22650));
    InMux I__5487 (
            .O(N__22676),
            .I(N__22647));
    LocalMux I__5486 (
            .O(N__22673),
            .I(N__22642));
    LocalMux I__5485 (
            .O(N__22670),
            .I(N__22642));
    Span4Mux_v I__5484 (
            .O(N__22667),
            .I(N__22637));
    LocalMux I__5483 (
            .O(N__22664),
            .I(N__22637));
    InMux I__5482 (
            .O(N__22661),
            .I(N__22634));
    Span4Mux_h I__5481 (
            .O(N__22658),
            .I(N__22631));
    Span4Mux_h I__5480 (
            .O(N__22655),
            .I(N__22624));
    LocalMux I__5479 (
            .O(N__22650),
            .I(N__22624));
    LocalMux I__5478 (
            .O(N__22647),
            .I(N__22624));
    Span4Mux_h I__5477 (
            .O(N__22642),
            .I(N__22621));
    Span4Mux_h I__5476 (
            .O(N__22637),
            .I(N__22618));
    LocalMux I__5475 (
            .O(N__22634),
            .I(\b2v_inst1.r_RX_DataZ0 ));
    Odrv4 I__5474 (
            .O(N__22631),
            .I(\b2v_inst1.r_RX_DataZ0 ));
    Odrv4 I__5473 (
            .O(N__22624),
            .I(\b2v_inst1.r_RX_DataZ0 ));
    Odrv4 I__5472 (
            .O(N__22621),
            .I(\b2v_inst1.r_RX_DataZ0 ));
    Odrv4 I__5471 (
            .O(N__22618),
            .I(\b2v_inst1.r_RX_DataZ0 ));
    ClkMux I__5470 (
            .O(N__22607),
            .I(N__22602));
    ClkMux I__5469 (
            .O(N__22606),
            .I(N__22599));
    ClkMux I__5468 (
            .O(N__22605),
            .I(N__22590));
    LocalMux I__5467 (
            .O(N__22602),
            .I(N__22582));
    LocalMux I__5466 (
            .O(N__22599),
            .I(N__22582));
    ClkMux I__5465 (
            .O(N__22598),
            .I(N__22579));
    ClkMux I__5464 (
            .O(N__22597),
            .I(N__22574));
    ClkMux I__5463 (
            .O(N__22596),
            .I(N__22566));
    ClkMux I__5462 (
            .O(N__22595),
            .I(N__22558));
    ClkMux I__5461 (
            .O(N__22594),
            .I(N__22555));
    ClkMux I__5460 (
            .O(N__22593),
            .I(N__22551));
    LocalMux I__5459 (
            .O(N__22590),
            .I(N__22547));
    ClkMux I__5458 (
            .O(N__22589),
            .I(N__22544));
    ClkMux I__5457 (
            .O(N__22588),
            .I(N__22541));
    ClkMux I__5456 (
            .O(N__22587),
            .I(N__22538));
    Span4Mux_v I__5455 (
            .O(N__22582),
            .I(N__22533));
    LocalMux I__5454 (
            .O(N__22579),
            .I(N__22533));
    ClkMux I__5453 (
            .O(N__22578),
            .I(N__22530));
    ClkMux I__5452 (
            .O(N__22577),
            .I(N__22527));
    LocalMux I__5451 (
            .O(N__22574),
            .I(N__22524));
    ClkMux I__5450 (
            .O(N__22573),
            .I(N__22521));
    ClkMux I__5449 (
            .O(N__22572),
            .I(N__22518));
    ClkMux I__5448 (
            .O(N__22571),
            .I(N__22511));
    ClkMux I__5447 (
            .O(N__22570),
            .I(N__22506));
    ClkMux I__5446 (
            .O(N__22569),
            .I(N__22503));
    LocalMux I__5445 (
            .O(N__22566),
            .I(N__22497));
    ClkMux I__5444 (
            .O(N__22565),
            .I(N__22493));
    ClkMux I__5443 (
            .O(N__22564),
            .I(N__22490));
    ClkMux I__5442 (
            .O(N__22563),
            .I(N__22487));
    ClkMux I__5441 (
            .O(N__22562),
            .I(N__22484));
    ClkMux I__5440 (
            .O(N__22561),
            .I(N__22477));
    LocalMux I__5439 (
            .O(N__22558),
            .I(N__22472));
    LocalMux I__5438 (
            .O(N__22555),
            .I(N__22472));
    ClkMux I__5437 (
            .O(N__22554),
            .I(N__22469));
    LocalMux I__5436 (
            .O(N__22551),
            .I(N__22465));
    ClkMux I__5435 (
            .O(N__22550),
            .I(N__22462));
    Span4Mux_v I__5434 (
            .O(N__22547),
            .I(N__22456));
    LocalMux I__5433 (
            .O(N__22544),
            .I(N__22456));
    LocalMux I__5432 (
            .O(N__22541),
            .I(N__22448));
    LocalMux I__5431 (
            .O(N__22538),
            .I(N__22448));
    Span4Mux_v I__5430 (
            .O(N__22533),
            .I(N__22444));
    LocalMux I__5429 (
            .O(N__22530),
            .I(N__22439));
    LocalMux I__5428 (
            .O(N__22527),
            .I(N__22439));
    Span4Mux_h I__5427 (
            .O(N__22524),
            .I(N__22432));
    LocalMux I__5426 (
            .O(N__22521),
            .I(N__22432));
    LocalMux I__5425 (
            .O(N__22518),
            .I(N__22432));
    ClkMux I__5424 (
            .O(N__22517),
            .I(N__22429));
    ClkMux I__5423 (
            .O(N__22516),
            .I(N__22426));
    ClkMux I__5422 (
            .O(N__22515),
            .I(N__22423));
    ClkMux I__5421 (
            .O(N__22514),
            .I(N__22420));
    LocalMux I__5420 (
            .O(N__22511),
            .I(N__22416));
    ClkMux I__5419 (
            .O(N__22510),
            .I(N__22413));
    ClkMux I__5418 (
            .O(N__22509),
            .I(N__22407));
    LocalMux I__5417 (
            .O(N__22506),
            .I(N__22402));
    LocalMux I__5416 (
            .O(N__22503),
            .I(N__22399));
    ClkMux I__5415 (
            .O(N__22502),
            .I(N__22396));
    ClkMux I__5414 (
            .O(N__22501),
            .I(N__22393));
    ClkMux I__5413 (
            .O(N__22500),
            .I(N__22389));
    Span4Mux_v I__5412 (
            .O(N__22497),
            .I(N__22385));
    ClkMux I__5411 (
            .O(N__22496),
            .I(N__22382));
    LocalMux I__5410 (
            .O(N__22493),
            .I(N__22377));
    LocalMux I__5409 (
            .O(N__22490),
            .I(N__22374));
    LocalMux I__5408 (
            .O(N__22487),
            .I(N__22371));
    LocalMux I__5407 (
            .O(N__22484),
            .I(N__22368));
    ClkMux I__5406 (
            .O(N__22483),
            .I(N__22365));
    ClkMux I__5405 (
            .O(N__22482),
            .I(N__22362));
    ClkMux I__5404 (
            .O(N__22481),
            .I(N__22359));
    ClkMux I__5403 (
            .O(N__22480),
            .I(N__22356));
    LocalMux I__5402 (
            .O(N__22477),
            .I(N__22348));
    Span4Mux_v I__5401 (
            .O(N__22472),
            .I(N__22343));
    LocalMux I__5400 (
            .O(N__22469),
            .I(N__22343));
    ClkMux I__5399 (
            .O(N__22468),
            .I(N__22340));
    Span4Mux_h I__5398 (
            .O(N__22465),
            .I(N__22335));
    LocalMux I__5397 (
            .O(N__22462),
            .I(N__22335));
    ClkMux I__5396 (
            .O(N__22461),
            .I(N__22332));
    Span4Mux_h I__5395 (
            .O(N__22456),
            .I(N__22329));
    ClkMux I__5394 (
            .O(N__22455),
            .I(N__22326));
    ClkMux I__5393 (
            .O(N__22454),
            .I(N__22323));
    ClkMux I__5392 (
            .O(N__22453),
            .I(N__22320));
    Span4Mux_v I__5391 (
            .O(N__22448),
            .I(N__22315));
    ClkMux I__5390 (
            .O(N__22447),
            .I(N__22312));
    Span4Mux_h I__5389 (
            .O(N__22444),
            .I(N__22297));
    Span4Mux_h I__5388 (
            .O(N__22439),
            .I(N__22297));
    Span4Mux_v I__5387 (
            .O(N__22432),
            .I(N__22297));
    LocalMux I__5386 (
            .O(N__22429),
            .I(N__22297));
    LocalMux I__5385 (
            .O(N__22426),
            .I(N__22297));
    LocalMux I__5384 (
            .O(N__22423),
            .I(N__22297));
    LocalMux I__5383 (
            .O(N__22420),
            .I(N__22297));
    ClkMux I__5382 (
            .O(N__22419),
            .I(N__22294));
    Span4Mux_v I__5381 (
            .O(N__22416),
            .I(N__22291));
    LocalMux I__5380 (
            .O(N__22413),
            .I(N__22288));
    ClkMux I__5379 (
            .O(N__22412),
            .I(N__22285));
    ClkMux I__5378 (
            .O(N__22411),
            .I(N__22282));
    ClkMux I__5377 (
            .O(N__22410),
            .I(N__22277));
    LocalMux I__5376 (
            .O(N__22407),
            .I(N__22274));
    ClkMux I__5375 (
            .O(N__22406),
            .I(N__22271));
    ClkMux I__5374 (
            .O(N__22405),
            .I(N__22268));
    Span4Mux_v I__5373 (
            .O(N__22402),
            .I(N__22264));
    Span4Mux_v I__5372 (
            .O(N__22399),
            .I(N__22256));
    LocalMux I__5371 (
            .O(N__22396),
            .I(N__22256));
    LocalMux I__5370 (
            .O(N__22393),
            .I(N__22256));
    ClkMux I__5369 (
            .O(N__22392),
            .I(N__22253));
    LocalMux I__5368 (
            .O(N__22389),
            .I(N__22248));
    ClkMux I__5367 (
            .O(N__22388),
            .I(N__22245));
    Span4Mux_v I__5366 (
            .O(N__22385),
            .I(N__22237));
    LocalMux I__5365 (
            .O(N__22382),
            .I(N__22237));
    ClkMux I__5364 (
            .O(N__22381),
            .I(N__22234));
    ClkMux I__5363 (
            .O(N__22380),
            .I(N__22231));
    Span4Mux_v I__5362 (
            .O(N__22377),
            .I(N__22219));
    Span4Mux_h I__5361 (
            .O(N__22374),
            .I(N__22219));
    Span4Mux_h I__5360 (
            .O(N__22371),
            .I(N__22219));
    Span4Mux_h I__5359 (
            .O(N__22368),
            .I(N__22219));
    LocalMux I__5358 (
            .O(N__22365),
            .I(N__22219));
    LocalMux I__5357 (
            .O(N__22362),
            .I(N__22216));
    LocalMux I__5356 (
            .O(N__22359),
            .I(N__22213));
    LocalMux I__5355 (
            .O(N__22356),
            .I(N__22210));
    ClkMux I__5354 (
            .O(N__22355),
            .I(N__22207));
    ClkMux I__5353 (
            .O(N__22354),
            .I(N__22204));
    ClkMux I__5352 (
            .O(N__22353),
            .I(N__22201));
    ClkMux I__5351 (
            .O(N__22352),
            .I(N__22198));
    ClkMux I__5350 (
            .O(N__22351),
            .I(N__22195));
    Span4Mux_v I__5349 (
            .O(N__22348),
            .I(N__22188));
    Span4Mux_v I__5348 (
            .O(N__22343),
            .I(N__22188));
    LocalMux I__5347 (
            .O(N__22340),
            .I(N__22188));
    Span4Mux_v I__5346 (
            .O(N__22335),
            .I(N__22182));
    LocalMux I__5345 (
            .O(N__22332),
            .I(N__22182));
    Span4Mux_h I__5344 (
            .O(N__22329),
            .I(N__22177));
    LocalMux I__5343 (
            .O(N__22326),
            .I(N__22177));
    LocalMux I__5342 (
            .O(N__22323),
            .I(N__22174));
    LocalMux I__5341 (
            .O(N__22320),
            .I(N__22171));
    ClkMux I__5340 (
            .O(N__22319),
            .I(N__22168));
    ClkMux I__5339 (
            .O(N__22318),
            .I(N__22165));
    Span4Mux_h I__5338 (
            .O(N__22315),
            .I(N__22162));
    LocalMux I__5337 (
            .O(N__22312),
            .I(N__22155));
    Span4Mux_v I__5336 (
            .O(N__22297),
            .I(N__22155));
    LocalMux I__5335 (
            .O(N__22294),
            .I(N__22155));
    Span4Mux_h I__5334 (
            .O(N__22291),
            .I(N__22150));
    Span4Mux_h I__5333 (
            .O(N__22288),
            .I(N__22150));
    LocalMux I__5332 (
            .O(N__22285),
            .I(N__22145));
    LocalMux I__5331 (
            .O(N__22282),
            .I(N__22145));
    ClkMux I__5330 (
            .O(N__22281),
            .I(N__22142));
    ClkMux I__5329 (
            .O(N__22280),
            .I(N__22139));
    LocalMux I__5328 (
            .O(N__22277),
            .I(N__22136));
    Span4Mux_h I__5327 (
            .O(N__22274),
            .I(N__22129));
    LocalMux I__5326 (
            .O(N__22271),
            .I(N__22129));
    LocalMux I__5325 (
            .O(N__22268),
            .I(N__22129));
    ClkMux I__5324 (
            .O(N__22267),
            .I(N__22126));
    Span4Mux_h I__5323 (
            .O(N__22264),
            .I(N__22123));
    ClkMux I__5322 (
            .O(N__22263),
            .I(N__22120));
    Span4Mux_v I__5321 (
            .O(N__22256),
            .I(N__22115));
    LocalMux I__5320 (
            .O(N__22253),
            .I(N__22115));
    ClkMux I__5319 (
            .O(N__22252),
            .I(N__22111));
    ClkMux I__5318 (
            .O(N__22251),
            .I(N__22108));
    Span4Mux_v I__5317 (
            .O(N__22248),
            .I(N__22103));
    LocalMux I__5316 (
            .O(N__22245),
            .I(N__22103));
    ClkMux I__5315 (
            .O(N__22244),
            .I(N__22099));
    ClkMux I__5314 (
            .O(N__22243),
            .I(N__22096));
    ClkMux I__5313 (
            .O(N__22242),
            .I(N__22093));
    Span4Mux_v I__5312 (
            .O(N__22237),
            .I(N__22090));
    LocalMux I__5311 (
            .O(N__22234),
            .I(N__22085));
    LocalMux I__5310 (
            .O(N__22231),
            .I(N__22085));
    ClkMux I__5309 (
            .O(N__22230),
            .I(N__22078));
    Span4Mux_v I__5308 (
            .O(N__22219),
            .I(N__22075));
    Span4Mux_h I__5307 (
            .O(N__22216),
            .I(N__22072));
    Span4Mux_v I__5306 (
            .O(N__22213),
            .I(N__22069));
    Span4Mux_v I__5305 (
            .O(N__22210),
            .I(N__22064));
    LocalMux I__5304 (
            .O(N__22207),
            .I(N__22064));
    LocalMux I__5303 (
            .O(N__22204),
            .I(N__22053));
    LocalMux I__5302 (
            .O(N__22201),
            .I(N__22053));
    LocalMux I__5301 (
            .O(N__22198),
            .I(N__22053));
    LocalMux I__5300 (
            .O(N__22195),
            .I(N__22053));
    Span4Mux_h I__5299 (
            .O(N__22188),
            .I(N__22053));
    ClkMux I__5298 (
            .O(N__22187),
            .I(N__22050));
    Span4Mux_h I__5297 (
            .O(N__22182),
            .I(N__22047));
    Span4Mux_v I__5296 (
            .O(N__22177),
            .I(N__22044));
    Span4Mux_h I__5295 (
            .O(N__22174),
            .I(N__22035));
    Span4Mux_v I__5294 (
            .O(N__22171),
            .I(N__22035));
    LocalMux I__5293 (
            .O(N__22168),
            .I(N__22035));
    LocalMux I__5292 (
            .O(N__22165),
            .I(N__22035));
    Span4Mux_h I__5291 (
            .O(N__22162),
            .I(N__22030));
    Span4Mux_v I__5290 (
            .O(N__22155),
            .I(N__22030));
    Span4Mux_v I__5289 (
            .O(N__22150),
            .I(N__22021));
    Span4Mux_v I__5288 (
            .O(N__22145),
            .I(N__22021));
    LocalMux I__5287 (
            .O(N__22142),
            .I(N__22021));
    LocalMux I__5286 (
            .O(N__22139),
            .I(N__22021));
    Span4Mux_h I__5285 (
            .O(N__22136),
            .I(N__22014));
    Span4Mux_v I__5284 (
            .O(N__22129),
            .I(N__22014));
    LocalMux I__5283 (
            .O(N__22126),
            .I(N__22014));
    Span4Mux_v I__5282 (
            .O(N__22123),
            .I(N__22009));
    LocalMux I__5281 (
            .O(N__22120),
            .I(N__22009));
    Span4Mux_v I__5280 (
            .O(N__22115),
            .I(N__22006));
    ClkMux I__5279 (
            .O(N__22114),
            .I(N__22003));
    LocalMux I__5278 (
            .O(N__22111),
            .I(N__21998));
    LocalMux I__5277 (
            .O(N__22108),
            .I(N__21998));
    Span4Mux_v I__5276 (
            .O(N__22103),
            .I(N__21995));
    ClkMux I__5275 (
            .O(N__22102),
            .I(N__21992));
    LocalMux I__5274 (
            .O(N__22099),
            .I(N__21989));
    LocalMux I__5273 (
            .O(N__22096),
            .I(N__21986));
    LocalMux I__5272 (
            .O(N__22093),
            .I(N__21983));
    Span4Mux_h I__5271 (
            .O(N__22090),
            .I(N__21978));
    Span4Mux_v I__5270 (
            .O(N__22085),
            .I(N__21978));
    ClkMux I__5269 (
            .O(N__22084),
            .I(N__21975));
    ClkMux I__5268 (
            .O(N__22083),
            .I(N__21972));
    ClkMux I__5267 (
            .O(N__22082),
            .I(N__21968));
    ClkMux I__5266 (
            .O(N__22081),
            .I(N__21965));
    LocalMux I__5265 (
            .O(N__22078),
            .I(N__21961));
    Span4Mux_h I__5264 (
            .O(N__22075),
            .I(N__21948));
    Span4Mux_h I__5263 (
            .O(N__22072),
            .I(N__21948));
    Span4Mux_h I__5262 (
            .O(N__22069),
            .I(N__21948));
    Span4Mux_v I__5261 (
            .O(N__22064),
            .I(N__21948));
    Span4Mux_v I__5260 (
            .O(N__22053),
            .I(N__21948));
    LocalMux I__5259 (
            .O(N__22050),
            .I(N__21948));
    Span4Mux_v I__5258 (
            .O(N__22047),
            .I(N__21940));
    Span4Mux_h I__5257 (
            .O(N__22044),
            .I(N__21940));
    Span4Mux_v I__5256 (
            .O(N__22035),
            .I(N__21937));
    Span4Mux_h I__5255 (
            .O(N__22030),
            .I(N__21932));
    Span4Mux_v I__5254 (
            .O(N__22021),
            .I(N__21932));
    Span4Mux_h I__5253 (
            .O(N__22014),
            .I(N__21923));
    Span4Mux_h I__5252 (
            .O(N__22009),
            .I(N__21923));
    Span4Mux_v I__5251 (
            .O(N__22006),
            .I(N__21923));
    LocalMux I__5250 (
            .O(N__22003),
            .I(N__21923));
    Span4Mux_v I__5249 (
            .O(N__21998),
            .I(N__21916));
    Span4Mux_v I__5248 (
            .O(N__21995),
            .I(N__21916));
    LocalMux I__5247 (
            .O(N__21992),
            .I(N__21916));
    Span4Mux_v I__5246 (
            .O(N__21989),
            .I(N__21905));
    Span4Mux_v I__5245 (
            .O(N__21986),
            .I(N__21905));
    Span4Mux_v I__5244 (
            .O(N__21983),
            .I(N__21905));
    Span4Mux_h I__5243 (
            .O(N__21978),
            .I(N__21905));
    LocalMux I__5242 (
            .O(N__21975),
            .I(N__21905));
    LocalMux I__5241 (
            .O(N__21972),
            .I(N__21902));
    ClkMux I__5240 (
            .O(N__21971),
            .I(N__21899));
    LocalMux I__5239 (
            .O(N__21968),
            .I(N__21894));
    LocalMux I__5238 (
            .O(N__21965),
            .I(N__21894));
    ClkMux I__5237 (
            .O(N__21964),
            .I(N__21891));
    Span4Mux_h I__5236 (
            .O(N__21961),
            .I(N__21885));
    Span4Mux_v I__5235 (
            .O(N__21948),
            .I(N__21885));
    ClkMux I__5234 (
            .O(N__21947),
            .I(N__21881));
    ClkMux I__5233 (
            .O(N__21946),
            .I(N__21878));
    ClkMux I__5232 (
            .O(N__21945),
            .I(N__21875));
    Span4Mux_h I__5231 (
            .O(N__21940),
            .I(N__21871));
    Span4Mux_h I__5230 (
            .O(N__21937),
            .I(N__21866));
    Span4Mux_h I__5229 (
            .O(N__21932),
            .I(N__21866));
    Span4Mux_h I__5228 (
            .O(N__21923),
            .I(N__21861));
    Span4Mux_v I__5227 (
            .O(N__21916),
            .I(N__21861));
    Span4Mux_v I__5226 (
            .O(N__21905),
            .I(N__21850));
    Span4Mux_v I__5225 (
            .O(N__21902),
            .I(N__21850));
    LocalMux I__5224 (
            .O(N__21899),
            .I(N__21850));
    Span4Mux_v I__5223 (
            .O(N__21894),
            .I(N__21850));
    LocalMux I__5222 (
            .O(N__21891),
            .I(N__21850));
    ClkMux I__5221 (
            .O(N__21890),
            .I(N__21847));
    Span4Mux_h I__5220 (
            .O(N__21885),
            .I(N__21844));
    ClkMux I__5219 (
            .O(N__21884),
            .I(N__21841));
    LocalMux I__5218 (
            .O(N__21881),
            .I(N__21838));
    LocalMux I__5217 (
            .O(N__21878),
            .I(N__21833));
    LocalMux I__5216 (
            .O(N__21875),
            .I(N__21833));
    ClkMux I__5215 (
            .O(N__21874),
            .I(N__21830));
    Span4Mux_h I__5214 (
            .O(N__21871),
            .I(N__21827));
    Span4Mux_h I__5213 (
            .O(N__21866),
            .I(N__21824));
    Span4Mux_h I__5212 (
            .O(N__21861),
            .I(N__21821));
    Sp12to4 I__5211 (
            .O(N__21850),
            .I(N__21818));
    LocalMux I__5210 (
            .O(N__21847),
            .I(N__21811));
    Sp12to4 I__5209 (
            .O(N__21844),
            .I(N__21811));
    LocalMux I__5208 (
            .O(N__21841),
            .I(N__21811));
    Span4Mux_h I__5207 (
            .O(N__21838),
            .I(N__21804));
    Span4Mux_v I__5206 (
            .O(N__21833),
            .I(N__21804));
    LocalMux I__5205 (
            .O(N__21830),
            .I(N__21804));
    Span4Mux_h I__5204 (
            .O(N__21827),
            .I(N__21801));
    Span4Mux_h I__5203 (
            .O(N__21824),
            .I(N__21798));
    Sp12to4 I__5202 (
            .O(N__21821),
            .I(N__21793));
    Span12Mux_h I__5201 (
            .O(N__21818),
            .I(N__21793));
    Span12Mux_v I__5200 (
            .O(N__21811),
            .I(N__21788));
    Sp12to4 I__5199 (
            .O(N__21804),
            .I(N__21788));
    IoSpan4Mux I__5198 (
            .O(N__21801),
            .I(N__21785));
    Span4Mux_h I__5197 (
            .O(N__21798),
            .I(N__21782));
    Span12Mux_h I__5196 (
            .O(N__21793),
            .I(N__21779));
    Span12Mux_h I__5195 (
            .O(N__21788),
            .I(N__21776));
    Odrv4 I__5194 (
            .O(N__21785),
            .I(clk));
    Odrv4 I__5193 (
            .O(N__21782),
            .I(clk));
    Odrv12 I__5192 (
            .O(N__21779),
            .I(clk));
    Odrv12 I__5191 (
            .O(N__21776),
            .I(clk));
    InMux I__5190 (
            .O(N__21767),
            .I(N__21763));
    InMux I__5189 (
            .O(N__21766),
            .I(N__21760));
    LocalMux I__5188 (
            .O(N__21763),
            .I(N__21757));
    LocalMux I__5187 (
            .O(N__21760),
            .I(\b2v_inst1.N_29_mux ));
    Odrv4 I__5186 (
            .O(N__21757),
            .I(\b2v_inst1.N_29_mux ));
    CascadeMux I__5185 (
            .O(N__21752),
            .I(\b2v_inst1.r_SM_Main_1_sqmuxa_1_cascade_ ));
    InMux I__5184 (
            .O(N__21749),
            .I(N__21742));
    InMux I__5183 (
            .O(N__21748),
            .I(N__21742));
    InMux I__5182 (
            .O(N__21747),
            .I(N__21739));
    LocalMux I__5181 (
            .O(N__21742),
            .I(\b2v_inst1.un1_r_SM_Main_1_sqmuxa_0 ));
    LocalMux I__5180 (
            .O(N__21739),
            .I(\b2v_inst1.un1_r_SM_Main_1_sqmuxa_0 ));
    InMux I__5179 (
            .O(N__21734),
            .I(N__21729));
    InMux I__5178 (
            .O(N__21733),
            .I(N__21726));
    InMux I__5177 (
            .O(N__21732),
            .I(N__21720));
    LocalMux I__5176 (
            .O(N__21729),
            .I(N__21715));
    LocalMux I__5175 (
            .O(N__21726),
            .I(N__21715));
    InMux I__5174 (
            .O(N__21725),
            .I(N__21712));
    InMux I__5173 (
            .O(N__21724),
            .I(N__21709));
    InMux I__5172 (
            .O(N__21723),
            .I(N__21706));
    LocalMux I__5171 (
            .O(N__21720),
            .I(\b2v_inst1.un1_r_Clk_Count_ac0_1_out ));
    Odrv4 I__5170 (
            .O(N__21715),
            .I(\b2v_inst1.un1_r_Clk_Count_ac0_1_out ));
    LocalMux I__5169 (
            .O(N__21712),
            .I(\b2v_inst1.un1_r_Clk_Count_ac0_1_out ));
    LocalMux I__5168 (
            .O(N__21709),
            .I(\b2v_inst1.un1_r_Clk_Count_ac0_1_out ));
    LocalMux I__5167 (
            .O(N__21706),
            .I(\b2v_inst1.un1_r_Clk_Count_ac0_1_out ));
    CascadeMux I__5166 (
            .O(N__21695),
            .I(N__21686));
    InMux I__5165 (
            .O(N__21694),
            .I(N__21681));
    InMux I__5164 (
            .O(N__21693),
            .I(N__21681));
    CascadeMux I__5163 (
            .O(N__21692),
            .I(N__21678));
    CascadeMux I__5162 (
            .O(N__21691),
            .I(N__21675));
    InMux I__5161 (
            .O(N__21690),
            .I(N__21670));
    InMux I__5160 (
            .O(N__21689),
            .I(N__21670));
    InMux I__5159 (
            .O(N__21686),
            .I(N__21667));
    LocalMux I__5158 (
            .O(N__21681),
            .I(N__21663));
    InMux I__5157 (
            .O(N__21678),
            .I(N__21653));
    InMux I__5156 (
            .O(N__21675),
            .I(N__21650));
    LocalMux I__5155 (
            .O(N__21670),
            .I(N__21647));
    LocalMux I__5154 (
            .O(N__21667),
            .I(N__21644));
    CascadeMux I__5153 (
            .O(N__21666),
            .I(N__21640));
    Span4Mux_h I__5152 (
            .O(N__21663),
            .I(N__21636));
    InMux I__5151 (
            .O(N__21662),
            .I(N__21633));
    InMux I__5150 (
            .O(N__21661),
            .I(N__21626));
    InMux I__5149 (
            .O(N__21660),
            .I(N__21626));
    InMux I__5148 (
            .O(N__21659),
            .I(N__21626));
    InMux I__5147 (
            .O(N__21658),
            .I(N__21623));
    InMux I__5146 (
            .O(N__21657),
            .I(N__21620));
    InMux I__5145 (
            .O(N__21656),
            .I(N__21617));
    LocalMux I__5144 (
            .O(N__21653),
            .I(N__21612));
    LocalMux I__5143 (
            .O(N__21650),
            .I(N__21612));
    Span4Mux_h I__5142 (
            .O(N__21647),
            .I(N__21607));
    Span4Mux_h I__5141 (
            .O(N__21644),
            .I(N__21607));
    InMux I__5140 (
            .O(N__21643),
            .I(N__21600));
    InMux I__5139 (
            .O(N__21640),
            .I(N__21600));
    InMux I__5138 (
            .O(N__21639),
            .I(N__21600));
    Odrv4 I__5137 (
            .O(N__21636),
            .I(\b2v_inst1.r_Clk_CountZ0Z_3 ));
    LocalMux I__5136 (
            .O(N__21633),
            .I(\b2v_inst1.r_Clk_CountZ0Z_3 ));
    LocalMux I__5135 (
            .O(N__21626),
            .I(\b2v_inst1.r_Clk_CountZ0Z_3 ));
    LocalMux I__5134 (
            .O(N__21623),
            .I(\b2v_inst1.r_Clk_CountZ0Z_3 ));
    LocalMux I__5133 (
            .O(N__21620),
            .I(\b2v_inst1.r_Clk_CountZ0Z_3 ));
    LocalMux I__5132 (
            .O(N__21617),
            .I(\b2v_inst1.r_Clk_CountZ0Z_3 ));
    Odrv4 I__5131 (
            .O(N__21612),
            .I(\b2v_inst1.r_Clk_CountZ0Z_3 ));
    Odrv4 I__5130 (
            .O(N__21607),
            .I(\b2v_inst1.r_Clk_CountZ0Z_3 ));
    LocalMux I__5129 (
            .O(N__21600),
            .I(\b2v_inst1.r_Clk_CountZ0Z_3 ));
    CascadeMux I__5128 (
            .O(N__21581),
            .I(\b2v_inst1.g0_3_1_cascade_ ));
    InMux I__5127 (
            .O(N__21578),
            .I(N__21575));
    LocalMux I__5126 (
            .O(N__21575),
            .I(\b2v_inst1.N_14_0_0 ));
    CascadeMux I__5125 (
            .O(N__21572),
            .I(\b2v_inst1.N_14_0_0_cascade_ ));
    InMux I__5124 (
            .O(N__21569),
            .I(N__21566));
    LocalMux I__5123 (
            .O(N__21566),
            .I(\b2v_inst1.N_29_mux_0 ));
    InMux I__5122 (
            .O(N__21563),
            .I(N__21556));
    CascadeMux I__5121 (
            .O(N__21562),
            .I(N__21553));
    InMux I__5120 (
            .O(N__21561),
            .I(N__21549));
    InMux I__5119 (
            .O(N__21560),
            .I(N__21544));
    InMux I__5118 (
            .O(N__21559),
            .I(N__21544));
    LocalMux I__5117 (
            .O(N__21556),
            .I(N__21539));
    InMux I__5116 (
            .O(N__21553),
            .I(N__21534));
    InMux I__5115 (
            .O(N__21552),
            .I(N__21534));
    LocalMux I__5114 (
            .O(N__21549),
            .I(N__21522));
    LocalMux I__5113 (
            .O(N__21544),
            .I(N__21522));
    InMux I__5112 (
            .O(N__21543),
            .I(N__21517));
    InMux I__5111 (
            .O(N__21542),
            .I(N__21517));
    Span4Mux_v I__5110 (
            .O(N__21539),
            .I(N__21512));
    LocalMux I__5109 (
            .O(N__21534),
            .I(N__21512));
    InMux I__5108 (
            .O(N__21533),
            .I(N__21507));
    InMux I__5107 (
            .O(N__21532),
            .I(N__21507));
    InMux I__5106 (
            .O(N__21531),
            .I(N__21500));
    InMux I__5105 (
            .O(N__21530),
            .I(N__21500));
    InMux I__5104 (
            .O(N__21529),
            .I(N__21500));
    InMux I__5103 (
            .O(N__21528),
            .I(N__21495));
    InMux I__5102 (
            .O(N__21527),
            .I(N__21495));
    Odrv4 I__5101 (
            .O(N__21522),
            .I(\b2v_inst1.r_Clk_CountZ0Z_0 ));
    LocalMux I__5100 (
            .O(N__21517),
            .I(\b2v_inst1.r_Clk_CountZ0Z_0 ));
    Odrv4 I__5099 (
            .O(N__21512),
            .I(\b2v_inst1.r_Clk_CountZ0Z_0 ));
    LocalMux I__5098 (
            .O(N__21507),
            .I(\b2v_inst1.r_Clk_CountZ0Z_0 ));
    LocalMux I__5097 (
            .O(N__21500),
            .I(\b2v_inst1.r_Clk_CountZ0Z_0 ));
    LocalMux I__5096 (
            .O(N__21495),
            .I(\b2v_inst1.r_Clk_CountZ0Z_0 ));
    CascadeMux I__5095 (
            .O(N__21482),
            .I(\b2v_inst1.g3_1_cascade_ ));
    InMux I__5094 (
            .O(N__21479),
            .I(N__21473));
    InMux I__5093 (
            .O(N__21478),
            .I(N__21468));
    InMux I__5092 (
            .O(N__21477),
            .I(N__21468));
    CascadeMux I__5091 (
            .O(N__21476),
            .I(N__21464));
    LocalMux I__5090 (
            .O(N__21473),
            .I(N__21457));
    LocalMux I__5089 (
            .O(N__21468),
            .I(N__21457));
    InMux I__5088 (
            .O(N__21467),
            .I(N__21450));
    InMux I__5087 (
            .O(N__21464),
            .I(N__21445));
    InMux I__5086 (
            .O(N__21463),
            .I(N__21445));
    CascadeMux I__5085 (
            .O(N__21462),
            .I(N__21440));
    Span4Mux_v I__5084 (
            .O(N__21457),
            .I(N__21436));
    InMux I__5083 (
            .O(N__21456),
            .I(N__21431));
    InMux I__5082 (
            .O(N__21455),
            .I(N__21431));
    InMux I__5081 (
            .O(N__21454),
            .I(N__21426));
    InMux I__5080 (
            .O(N__21453),
            .I(N__21426));
    LocalMux I__5079 (
            .O(N__21450),
            .I(N__21421));
    LocalMux I__5078 (
            .O(N__21445),
            .I(N__21421));
    InMux I__5077 (
            .O(N__21444),
            .I(N__21416));
    InMux I__5076 (
            .O(N__21443),
            .I(N__21416));
    InMux I__5075 (
            .O(N__21440),
            .I(N__21411));
    InMux I__5074 (
            .O(N__21439),
            .I(N__21411));
    Span4Mux_h I__5073 (
            .O(N__21436),
            .I(N__21404));
    LocalMux I__5072 (
            .O(N__21431),
            .I(N__21404));
    LocalMux I__5071 (
            .O(N__21426),
            .I(N__21404));
    Odrv4 I__5070 (
            .O(N__21421),
            .I(\b2v_inst1.r_Clk_CountZ0Z_1 ));
    LocalMux I__5069 (
            .O(N__21416),
            .I(\b2v_inst1.r_Clk_CountZ0Z_1 ));
    LocalMux I__5068 (
            .O(N__21411),
            .I(\b2v_inst1.r_Clk_CountZ0Z_1 ));
    Odrv4 I__5067 (
            .O(N__21404),
            .I(\b2v_inst1.r_Clk_CountZ0Z_1 ));
    InMux I__5066 (
            .O(N__21395),
            .I(N__21392));
    LocalMux I__5065 (
            .O(N__21392),
            .I(N__21389));
    Odrv4 I__5064 (
            .O(N__21389),
            .I(\b2v_inst1.g3 ));
    InMux I__5063 (
            .O(N__21386),
            .I(N__21383));
    LocalMux I__5062 (
            .O(N__21383),
            .I(N__21380));
    Odrv4 I__5061 (
            .O(N__21380),
            .I(\b2v_inst1.N_9_0 ));
    CascadeMux I__5060 (
            .O(N__21377),
            .I(\b2v_inst1.N_13_cascade_ ));
    InMux I__5059 (
            .O(N__21374),
            .I(N__21371));
    LocalMux I__5058 (
            .O(N__21371),
            .I(N__21368));
    Span4Mux_h I__5057 (
            .O(N__21368),
            .I(N__21365));
    Odrv4 I__5056 (
            .O(N__21365),
            .I(\b2v_inst1.g0_0_i_a6_3_0 ));
    CascadeMux I__5055 (
            .O(N__21362),
            .I(\b2v_inst1.g0_1_4_cascade_ ));
    InMux I__5054 (
            .O(N__21359),
            .I(N__21356));
    LocalMux I__5053 (
            .O(N__21356),
            .I(N__21348));
    CascadeMux I__5052 (
            .O(N__21355),
            .I(N__21345));
    CascadeMux I__5051 (
            .O(N__21354),
            .I(N__21342));
    InMux I__5050 (
            .O(N__21353),
            .I(N__21339));
    InMux I__5049 (
            .O(N__21352),
            .I(N__21336));
    InMux I__5048 (
            .O(N__21351),
            .I(N__21333));
    Span4Mux_h I__5047 (
            .O(N__21348),
            .I(N__21330));
    InMux I__5046 (
            .O(N__21345),
            .I(N__21327));
    InMux I__5045 (
            .O(N__21342),
            .I(N__21324));
    LocalMux I__5044 (
            .O(N__21339),
            .I(\b2v_inst1.N_28_mux ));
    LocalMux I__5043 (
            .O(N__21336),
            .I(\b2v_inst1.N_28_mux ));
    LocalMux I__5042 (
            .O(N__21333),
            .I(\b2v_inst1.N_28_mux ));
    Odrv4 I__5041 (
            .O(N__21330),
            .I(\b2v_inst1.N_28_mux ));
    LocalMux I__5040 (
            .O(N__21327),
            .I(\b2v_inst1.N_28_mux ));
    LocalMux I__5039 (
            .O(N__21324),
            .I(\b2v_inst1.N_28_mux ));
    InMux I__5038 (
            .O(N__21311),
            .I(N__21305));
    InMux I__5037 (
            .O(N__21310),
            .I(N__21305));
    LocalMux I__5036 (
            .O(N__21305),
            .I(N__21302));
    Odrv4 I__5035 (
            .O(N__21302),
            .I(\b2v_inst1.un1_r_SM_Main_3_0 ));
    CascadeMux I__5034 (
            .O(N__21299),
            .I(\b2v_inst1.g0_1_cascade_ ));
    InMux I__5033 (
            .O(N__21296),
            .I(N__21293));
    LocalMux I__5032 (
            .O(N__21293),
            .I(\b2v_inst1.N_29_mux_1 ));
    CascadeMux I__5031 (
            .O(N__21290),
            .I(\b2v_inst1.N_14_0_1_cascade_ ));
    CascadeMux I__5030 (
            .O(N__21287),
            .I(\b2v_inst1.g0_0_i_a6_1_5_cascade_ ));
    InMux I__5029 (
            .O(N__21284),
            .I(N__21281));
    LocalMux I__5028 (
            .O(N__21281),
            .I(\b2v_inst1.g0_0_i_a6_1_1 ));
    CascadeMux I__5027 (
            .O(N__21278),
            .I(N__21275));
    InMux I__5026 (
            .O(N__21275),
            .I(N__21272));
    LocalMux I__5025 (
            .O(N__21272),
            .I(\b2v_inst1.un1_r_Clk_Count_ac0_3_out ));
    CascadeMux I__5024 (
            .O(N__21269),
            .I(\b2v_inst.un8_dir_mem_3_ac0_9_0_cascade_ ));
    InMux I__5023 (
            .O(N__21266),
            .I(N__21262));
    InMux I__5022 (
            .O(N__21265),
            .I(N__21258));
    LocalMux I__5021 (
            .O(N__21262),
            .I(N__21255));
    InMux I__5020 (
            .O(N__21261),
            .I(N__21252));
    LocalMux I__5019 (
            .O(N__21258),
            .I(N__21248));
    Span4Mux_v I__5018 (
            .O(N__21255),
            .I(N__21243));
    LocalMux I__5017 (
            .O(N__21252),
            .I(N__21243));
    InMux I__5016 (
            .O(N__21251),
            .I(N__21240));
    Odrv4 I__5015 (
            .O(N__21248),
            .I(\b2v_inst.un10_indice ));
    Odrv4 I__5014 (
            .O(N__21243),
            .I(\b2v_inst.un10_indice ));
    LocalMux I__5013 (
            .O(N__21240),
            .I(\b2v_inst.un10_indice ));
    InMux I__5012 (
            .O(N__21233),
            .I(N__21229));
    InMux I__5011 (
            .O(N__21232),
            .I(N__21226));
    LocalMux I__5010 (
            .O(N__21229),
            .I(N__21215));
    LocalMux I__5009 (
            .O(N__21226),
            .I(N__21215));
    InMux I__5008 (
            .O(N__21225),
            .I(N__21210));
    InMux I__5007 (
            .O(N__21224),
            .I(N__21210));
    InMux I__5006 (
            .O(N__21223),
            .I(N__21207));
    InMux I__5005 (
            .O(N__21222),
            .I(N__21197));
    InMux I__5004 (
            .O(N__21221),
            .I(N__21197));
    InMux I__5003 (
            .O(N__21220),
            .I(N__21197));
    Span4Mux_h I__5002 (
            .O(N__21215),
            .I(N__21190));
    LocalMux I__5001 (
            .O(N__21210),
            .I(N__21190));
    LocalMux I__5000 (
            .O(N__21207),
            .I(N__21190));
    InMux I__4999 (
            .O(N__21206),
            .I(N__21183));
    InMux I__4998 (
            .O(N__21205),
            .I(N__21183));
    InMux I__4997 (
            .O(N__21204),
            .I(N__21183));
    LocalMux I__4996 (
            .O(N__21197),
            .I(\b2v_inst.indice_4_repZ0Z1 ));
    Odrv4 I__4995 (
            .O(N__21190),
            .I(\b2v_inst.indice_4_repZ0Z1 ));
    LocalMux I__4994 (
            .O(N__21183),
            .I(\b2v_inst.indice_4_repZ0Z1 ));
    InMux I__4993 (
            .O(N__21176),
            .I(N__21165));
    InMux I__4992 (
            .O(N__21175),
            .I(N__21165));
    InMux I__4991 (
            .O(N__21174),
            .I(N__21165));
    InMux I__4990 (
            .O(N__21173),
            .I(N__21162));
    InMux I__4989 (
            .O(N__21172),
            .I(N__21159));
    LocalMux I__4988 (
            .O(N__21165),
            .I(N__21152));
    LocalMux I__4987 (
            .O(N__21162),
            .I(N__21147));
    LocalMux I__4986 (
            .O(N__21159),
            .I(N__21147));
    InMux I__4985 (
            .O(N__21158),
            .I(N__21142));
    InMux I__4984 (
            .O(N__21157),
            .I(N__21135));
    InMux I__4983 (
            .O(N__21156),
            .I(N__21135));
    InMux I__4982 (
            .O(N__21155),
            .I(N__21135));
    Span4Mux_v I__4981 (
            .O(N__21152),
            .I(N__21128));
    Span4Mux_h I__4980 (
            .O(N__21147),
            .I(N__21128));
    InMux I__4979 (
            .O(N__21146),
            .I(N__21125));
    InMux I__4978 (
            .O(N__21145),
            .I(N__21122));
    LocalMux I__4977 (
            .O(N__21142),
            .I(N__21119));
    LocalMux I__4976 (
            .O(N__21135),
            .I(N__21116));
    InMux I__4975 (
            .O(N__21134),
            .I(N__21111));
    InMux I__4974 (
            .O(N__21133),
            .I(N__21111));
    Span4Mux_v I__4973 (
            .O(N__21128),
            .I(N__21106));
    LocalMux I__4972 (
            .O(N__21125),
            .I(N__21106));
    LocalMux I__4971 (
            .O(N__21122),
            .I(\b2v_inst.indice_1_repZ0Z2 ));
    Odrv12 I__4970 (
            .O(N__21119),
            .I(\b2v_inst.indice_1_repZ0Z2 ));
    Odrv4 I__4969 (
            .O(N__21116),
            .I(\b2v_inst.indice_1_repZ0Z2 ));
    LocalMux I__4968 (
            .O(N__21111),
            .I(\b2v_inst.indice_1_repZ0Z2 ));
    Odrv4 I__4967 (
            .O(N__21106),
            .I(\b2v_inst.indice_1_repZ0Z2 ));
    CascadeMux I__4966 (
            .O(N__21095),
            .I(N__21087));
    InMux I__4965 (
            .O(N__21094),
            .I(N__21080));
    InMux I__4964 (
            .O(N__21093),
            .I(N__21077));
    InMux I__4963 (
            .O(N__21092),
            .I(N__21072));
    InMux I__4962 (
            .O(N__21091),
            .I(N__21072));
    InMux I__4961 (
            .O(N__21090),
            .I(N__21069));
    InMux I__4960 (
            .O(N__21087),
            .I(N__21066));
    InMux I__4959 (
            .O(N__21086),
            .I(N__21063));
    CascadeMux I__4958 (
            .O(N__21085),
            .I(N__21060));
    InMux I__4957 (
            .O(N__21084),
            .I(N__21053));
    InMux I__4956 (
            .O(N__21083),
            .I(N__21053));
    LocalMux I__4955 (
            .O(N__21080),
            .I(N__21046));
    LocalMux I__4954 (
            .O(N__21077),
            .I(N__21046));
    LocalMux I__4953 (
            .O(N__21072),
            .I(N__21046));
    LocalMux I__4952 (
            .O(N__21069),
            .I(N__21039));
    LocalMux I__4951 (
            .O(N__21066),
            .I(N__21039));
    LocalMux I__4950 (
            .O(N__21063),
            .I(N__21039));
    InMux I__4949 (
            .O(N__21060),
            .I(N__21035));
    InMux I__4948 (
            .O(N__21059),
            .I(N__21032));
    InMux I__4947 (
            .O(N__21058),
            .I(N__21029));
    LocalMux I__4946 (
            .O(N__21053),
            .I(N__21024));
    Span4Mux_v I__4945 (
            .O(N__21046),
            .I(N__21024));
    Span4Mux_v I__4944 (
            .O(N__21039),
            .I(N__21021));
    InMux I__4943 (
            .O(N__21038),
            .I(N__21018));
    LocalMux I__4942 (
            .O(N__21035),
            .I(\b2v_inst.indice_0_repZ0Z2 ));
    LocalMux I__4941 (
            .O(N__21032),
            .I(\b2v_inst.indice_0_repZ0Z2 ));
    LocalMux I__4940 (
            .O(N__21029),
            .I(\b2v_inst.indice_0_repZ0Z2 ));
    Odrv4 I__4939 (
            .O(N__21024),
            .I(\b2v_inst.indice_0_repZ0Z2 ));
    Odrv4 I__4938 (
            .O(N__21021),
            .I(\b2v_inst.indice_0_repZ0Z2 ));
    LocalMux I__4937 (
            .O(N__21018),
            .I(\b2v_inst.indice_0_repZ0Z2 ));
    InMux I__4936 (
            .O(N__21005),
            .I(N__20997));
    InMux I__4935 (
            .O(N__21004),
            .I(N__20997));
    InMux I__4934 (
            .O(N__21003),
            .I(N__20994));
    CascadeMux I__4933 (
            .O(N__21002),
            .I(N__20991));
    LocalMux I__4932 (
            .O(N__20997),
            .I(N__20987));
    LocalMux I__4931 (
            .O(N__20994),
            .I(N__20984));
    InMux I__4930 (
            .O(N__20991),
            .I(N__20981));
    InMux I__4929 (
            .O(N__20990),
            .I(N__20978));
    Span4Mux_h I__4928 (
            .O(N__20987),
            .I(N__20975));
    Span4Mux_h I__4927 (
            .O(N__20984),
            .I(N__20972));
    LocalMux I__4926 (
            .O(N__20981),
            .I(N__20969));
    LocalMux I__4925 (
            .O(N__20978),
            .I(N__20966));
    Odrv4 I__4924 (
            .O(N__20975),
            .I(\b2v_inst.un10_indice_2_0 ));
    Odrv4 I__4923 (
            .O(N__20972),
            .I(\b2v_inst.un10_indice_2_0 ));
    Odrv4 I__4922 (
            .O(N__20969),
            .I(\b2v_inst.un10_indice_2_0 ));
    Odrv4 I__4921 (
            .O(N__20966),
            .I(\b2v_inst.un10_indice_2_0 ));
    InMux I__4920 (
            .O(N__20957),
            .I(N__20954));
    LocalMux I__4919 (
            .O(N__20954),
            .I(N__20950));
    CascadeMux I__4918 (
            .O(N__20953),
            .I(N__20947));
    Span4Mux_h I__4917 (
            .O(N__20950),
            .I(N__20944));
    InMux I__4916 (
            .O(N__20947),
            .I(N__20941));
    Odrv4 I__4915 (
            .O(N__20944),
            .I(\b2v_inst.un8_dir_mem_3_ac0_9_0 ));
    LocalMux I__4914 (
            .O(N__20941),
            .I(\b2v_inst.un8_dir_mem_3_ac0_9_0 ));
    InMux I__4913 (
            .O(N__20936),
            .I(N__20929));
    InMux I__4912 (
            .O(N__20935),
            .I(N__20924));
    InMux I__4911 (
            .O(N__20934),
            .I(N__20921));
    InMux I__4910 (
            .O(N__20933),
            .I(N__20918));
    InMux I__4909 (
            .O(N__20932),
            .I(N__20915));
    LocalMux I__4908 (
            .O(N__20929),
            .I(N__20909));
    InMux I__4907 (
            .O(N__20928),
            .I(N__20906));
    InMux I__4906 (
            .O(N__20927),
            .I(N__20903));
    LocalMux I__4905 (
            .O(N__20924),
            .I(N__20900));
    LocalMux I__4904 (
            .O(N__20921),
            .I(N__20890));
    LocalMux I__4903 (
            .O(N__20918),
            .I(N__20890));
    LocalMux I__4902 (
            .O(N__20915),
            .I(N__20890));
    InMux I__4901 (
            .O(N__20914),
            .I(N__20883));
    InMux I__4900 (
            .O(N__20913),
            .I(N__20883));
    InMux I__4899 (
            .O(N__20912),
            .I(N__20883));
    Span4Mux_v I__4898 (
            .O(N__20909),
            .I(N__20878));
    LocalMux I__4897 (
            .O(N__20906),
            .I(N__20878));
    LocalMux I__4896 (
            .O(N__20903),
            .I(N__20873));
    Span4Mux_h I__4895 (
            .O(N__20900),
            .I(N__20873));
    CascadeMux I__4894 (
            .O(N__20899),
            .I(N__20869));
    InMux I__4893 (
            .O(N__20898),
            .I(N__20862));
    InMux I__4892 (
            .O(N__20897),
            .I(N__20862));
    Span4Mux_v I__4891 (
            .O(N__20890),
            .I(N__20857));
    LocalMux I__4890 (
            .O(N__20883),
            .I(N__20857));
    Span4Mux_h I__4889 (
            .O(N__20878),
            .I(N__20852));
    Span4Mux_v I__4888 (
            .O(N__20873),
            .I(N__20852));
    InMux I__4887 (
            .O(N__20872),
            .I(N__20847));
    InMux I__4886 (
            .O(N__20869),
            .I(N__20847));
    InMux I__4885 (
            .O(N__20868),
            .I(N__20842));
    InMux I__4884 (
            .O(N__20867),
            .I(N__20842));
    LocalMux I__4883 (
            .O(N__20862),
            .I(\b2v_inst.indiceZ0Z_7 ));
    Odrv4 I__4882 (
            .O(N__20857),
            .I(\b2v_inst.indiceZ0Z_7 ));
    Odrv4 I__4881 (
            .O(N__20852),
            .I(\b2v_inst.indiceZ0Z_7 ));
    LocalMux I__4880 (
            .O(N__20847),
            .I(\b2v_inst.indiceZ0Z_7 ));
    LocalMux I__4879 (
            .O(N__20842),
            .I(\b2v_inst.indiceZ0Z_7 ));
    CascadeMux I__4878 (
            .O(N__20831),
            .I(N__20828));
    InMux I__4877 (
            .O(N__20828),
            .I(N__20815));
    InMux I__4876 (
            .O(N__20827),
            .I(N__20815));
    InMux I__4875 (
            .O(N__20826),
            .I(N__20815));
    InMux I__4874 (
            .O(N__20825),
            .I(N__20812));
    InMux I__4873 (
            .O(N__20824),
            .I(N__20809));
    InMux I__4872 (
            .O(N__20823),
            .I(N__20804));
    InMux I__4871 (
            .O(N__20822),
            .I(N__20804));
    LocalMux I__4870 (
            .O(N__20815),
            .I(N__20801));
    LocalMux I__4869 (
            .O(N__20812),
            .I(N__20798));
    LocalMux I__4868 (
            .O(N__20809),
            .I(N__20792));
    LocalMux I__4867 (
            .O(N__20804),
            .I(N__20792));
    Span4Mux_v I__4866 (
            .O(N__20801),
            .I(N__20789));
    Span4Mux_h I__4865 (
            .O(N__20798),
            .I(N__20786));
    InMux I__4864 (
            .O(N__20797),
            .I(N__20783));
    Span4Mux_v I__4863 (
            .O(N__20792),
            .I(N__20780));
    Span4Mux_h I__4862 (
            .O(N__20789),
            .I(N__20777));
    Odrv4 I__4861 (
            .O(N__20786),
            .I(\b2v_inst.un8_dir_mem_3_c4 ));
    LocalMux I__4860 (
            .O(N__20783),
            .I(\b2v_inst.un8_dir_mem_3_c4 ));
    Odrv4 I__4859 (
            .O(N__20780),
            .I(\b2v_inst.un8_dir_mem_3_c4 ));
    Odrv4 I__4858 (
            .O(N__20777),
            .I(\b2v_inst.un8_dir_mem_3_c4 ));
    CascadeMux I__4857 (
            .O(N__20768),
            .I(N__20765));
    InMux I__4856 (
            .O(N__20765),
            .I(N__20760));
    CascadeMux I__4855 (
            .O(N__20764),
            .I(N__20757));
    CascadeMux I__4854 (
            .O(N__20763),
            .I(N__20751));
    LocalMux I__4853 (
            .O(N__20760),
            .I(N__20748));
    InMux I__4852 (
            .O(N__20757),
            .I(N__20745));
    InMux I__4851 (
            .O(N__20756),
            .I(N__20742));
    InMux I__4850 (
            .O(N__20755),
            .I(N__20737));
    InMux I__4849 (
            .O(N__20754),
            .I(N__20737));
    InMux I__4848 (
            .O(N__20751),
            .I(N__20734));
    Odrv4 I__4847 (
            .O(N__20748),
            .I(\b2v_inst.indice_fastZ0Z_4 ));
    LocalMux I__4846 (
            .O(N__20745),
            .I(\b2v_inst.indice_fastZ0Z_4 ));
    LocalMux I__4845 (
            .O(N__20742),
            .I(\b2v_inst.indice_fastZ0Z_4 ));
    LocalMux I__4844 (
            .O(N__20737),
            .I(\b2v_inst.indice_fastZ0Z_4 ));
    LocalMux I__4843 (
            .O(N__20734),
            .I(\b2v_inst.indice_fastZ0Z_4 ));
    InMux I__4842 (
            .O(N__20723),
            .I(N__20719));
    InMux I__4841 (
            .O(N__20722),
            .I(N__20716));
    LocalMux I__4840 (
            .O(N__20719),
            .I(N__20713));
    LocalMux I__4839 (
            .O(N__20716),
            .I(N__20707));
    Span4Mux_h I__4838 (
            .O(N__20713),
            .I(N__20704));
    InMux I__4837 (
            .O(N__20712),
            .I(N__20699));
    InMux I__4836 (
            .O(N__20711),
            .I(N__20699));
    InMux I__4835 (
            .O(N__20710),
            .I(N__20696));
    Odrv12 I__4834 (
            .O(N__20707),
            .I(\b2v_inst.indice_fastZ0Z_3 ));
    Odrv4 I__4833 (
            .O(N__20704),
            .I(\b2v_inst.indice_fastZ0Z_3 ));
    LocalMux I__4832 (
            .O(N__20699),
            .I(\b2v_inst.indice_fastZ0Z_3 ));
    LocalMux I__4831 (
            .O(N__20696),
            .I(\b2v_inst.indice_fastZ0Z_3 ));
    InMux I__4830 (
            .O(N__20687),
            .I(N__20682));
    InMux I__4829 (
            .O(N__20686),
            .I(N__20677));
    InMux I__4828 (
            .O(N__20685),
            .I(N__20677));
    LocalMux I__4827 (
            .O(N__20682),
            .I(N__20674));
    LocalMux I__4826 (
            .O(N__20677),
            .I(N__20671));
    Odrv12 I__4825 (
            .O(N__20674),
            .I(\b2v_inst.un8_dir_mem_1_ac0_7_out ));
    Odrv4 I__4824 (
            .O(N__20671),
            .I(\b2v_inst.un8_dir_mem_1_ac0_7_out ));
    CascadeMux I__4823 (
            .O(N__20666),
            .I(N__20661));
    InMux I__4822 (
            .O(N__20665),
            .I(N__20658));
    InMux I__4821 (
            .O(N__20664),
            .I(N__20653));
    InMux I__4820 (
            .O(N__20661),
            .I(N__20653));
    LocalMux I__4819 (
            .O(N__20658),
            .I(N__20650));
    LocalMux I__4818 (
            .O(N__20653),
            .I(N__20647));
    Span4Mux_v I__4817 (
            .O(N__20650),
            .I(N__20642));
    Span4Mux_v I__4816 (
            .O(N__20647),
            .I(N__20642));
    Odrv4 I__4815 (
            .O(N__20642),
            .I(\b2v_inst.un8_dir_mem_2_c4 ));
    InMux I__4814 (
            .O(N__20639),
            .I(N__20627));
    InMux I__4813 (
            .O(N__20638),
            .I(N__20624));
    InMux I__4812 (
            .O(N__20637),
            .I(N__20621));
    InMux I__4811 (
            .O(N__20636),
            .I(N__20618));
    InMux I__4810 (
            .O(N__20635),
            .I(N__20614));
    InMux I__4809 (
            .O(N__20634),
            .I(N__20611));
    InMux I__4808 (
            .O(N__20633),
            .I(N__20605));
    InMux I__4807 (
            .O(N__20632),
            .I(N__20605));
    InMux I__4806 (
            .O(N__20631),
            .I(N__20600));
    InMux I__4805 (
            .O(N__20630),
            .I(N__20597));
    LocalMux I__4804 (
            .O(N__20627),
            .I(N__20588));
    LocalMux I__4803 (
            .O(N__20624),
            .I(N__20588));
    LocalMux I__4802 (
            .O(N__20621),
            .I(N__20588));
    LocalMux I__4801 (
            .O(N__20618),
            .I(N__20588));
    InMux I__4800 (
            .O(N__20617),
            .I(N__20585));
    LocalMux I__4799 (
            .O(N__20614),
            .I(N__20580));
    LocalMux I__4798 (
            .O(N__20611),
            .I(N__20580));
    InMux I__4797 (
            .O(N__20610),
            .I(N__20573));
    LocalMux I__4796 (
            .O(N__20605),
            .I(N__20570));
    InMux I__4795 (
            .O(N__20604),
            .I(N__20565));
    InMux I__4794 (
            .O(N__20603),
            .I(N__20565));
    LocalMux I__4793 (
            .O(N__20600),
            .I(N__20562));
    LocalMux I__4792 (
            .O(N__20597),
            .I(N__20558));
    Span4Mux_v I__4791 (
            .O(N__20588),
            .I(N__20550));
    LocalMux I__4790 (
            .O(N__20585),
            .I(N__20550));
    Span4Mux_v I__4789 (
            .O(N__20580),
            .I(N__20550));
    InMux I__4788 (
            .O(N__20579),
            .I(N__20547));
    InMux I__4787 (
            .O(N__20578),
            .I(N__20540));
    InMux I__4786 (
            .O(N__20577),
            .I(N__20540));
    InMux I__4785 (
            .O(N__20576),
            .I(N__20540));
    LocalMux I__4784 (
            .O(N__20573),
            .I(N__20531));
    Span12Mux_s11_v I__4783 (
            .O(N__20570),
            .I(N__20531));
    LocalMux I__4782 (
            .O(N__20565),
            .I(N__20531));
    Span12Mux_v I__4781 (
            .O(N__20562),
            .I(N__20531));
    InMux I__4780 (
            .O(N__20561),
            .I(N__20528));
    Span4Mux_v I__4779 (
            .O(N__20558),
            .I(N__20525));
    InMux I__4778 (
            .O(N__20557),
            .I(N__20522));
    Span4Mux_h I__4777 (
            .O(N__20550),
            .I(N__20519));
    LocalMux I__4776 (
            .O(N__20547),
            .I(\b2v_inst.indiceZ0Z_6 ));
    LocalMux I__4775 (
            .O(N__20540),
            .I(\b2v_inst.indiceZ0Z_6 ));
    Odrv12 I__4774 (
            .O(N__20531),
            .I(\b2v_inst.indiceZ0Z_6 ));
    LocalMux I__4773 (
            .O(N__20528),
            .I(\b2v_inst.indiceZ0Z_6 ));
    Odrv4 I__4772 (
            .O(N__20525),
            .I(\b2v_inst.indiceZ0Z_6 ));
    LocalMux I__4771 (
            .O(N__20522),
            .I(\b2v_inst.indiceZ0Z_6 ));
    Odrv4 I__4770 (
            .O(N__20519),
            .I(\b2v_inst.indiceZ0Z_6 ));
    InMux I__4769 (
            .O(N__20504),
            .I(N__20495));
    InMux I__4768 (
            .O(N__20503),
            .I(N__20495));
    InMux I__4767 (
            .O(N__20502),
            .I(N__20489));
    InMux I__4766 (
            .O(N__20501),
            .I(N__20486));
    CascadeMux I__4765 (
            .O(N__20500),
            .I(N__20479));
    LocalMux I__4764 (
            .O(N__20495),
            .I(N__20473));
    InMux I__4763 (
            .O(N__20494),
            .I(N__20468));
    InMux I__4762 (
            .O(N__20493),
            .I(N__20468));
    InMux I__4761 (
            .O(N__20492),
            .I(N__20465));
    LocalMux I__4760 (
            .O(N__20489),
            .I(N__20462));
    LocalMux I__4759 (
            .O(N__20486),
            .I(N__20459));
    InMux I__4758 (
            .O(N__20485),
            .I(N__20454));
    InMux I__4757 (
            .O(N__20484),
            .I(N__20454));
    InMux I__4756 (
            .O(N__20483),
            .I(N__20448));
    InMux I__4755 (
            .O(N__20482),
            .I(N__20448));
    InMux I__4754 (
            .O(N__20479),
            .I(N__20445));
    InMux I__4753 (
            .O(N__20478),
            .I(N__20442));
    InMux I__4752 (
            .O(N__20477),
            .I(N__20436));
    InMux I__4751 (
            .O(N__20476),
            .I(N__20436));
    Span4Mux_h I__4750 (
            .O(N__20473),
            .I(N__20425));
    LocalMux I__4749 (
            .O(N__20468),
            .I(N__20425));
    LocalMux I__4748 (
            .O(N__20465),
            .I(N__20425));
    Span4Mux_v I__4747 (
            .O(N__20462),
            .I(N__20425));
    Span4Mux_v I__4746 (
            .O(N__20459),
            .I(N__20425));
    LocalMux I__4745 (
            .O(N__20454),
            .I(N__20422));
    InMux I__4744 (
            .O(N__20453),
            .I(N__20419));
    LocalMux I__4743 (
            .O(N__20448),
            .I(N__20416));
    LocalMux I__4742 (
            .O(N__20445),
            .I(N__20411));
    LocalMux I__4741 (
            .O(N__20442),
            .I(N__20411));
    InMux I__4740 (
            .O(N__20441),
            .I(N__20408));
    LocalMux I__4739 (
            .O(N__20436),
            .I(N__20399));
    Span4Mux_v I__4738 (
            .O(N__20425),
            .I(N__20394));
    Span4Mux_v I__4737 (
            .O(N__20422),
            .I(N__20394));
    LocalMux I__4736 (
            .O(N__20419),
            .I(N__20391));
    Span4Mux_h I__4735 (
            .O(N__20416),
            .I(N__20384));
    Span4Mux_h I__4734 (
            .O(N__20411),
            .I(N__20384));
    LocalMux I__4733 (
            .O(N__20408),
            .I(N__20384));
    InMux I__4732 (
            .O(N__20407),
            .I(N__20375));
    InMux I__4731 (
            .O(N__20406),
            .I(N__20375));
    InMux I__4730 (
            .O(N__20405),
            .I(N__20375));
    InMux I__4729 (
            .O(N__20404),
            .I(N__20375));
    InMux I__4728 (
            .O(N__20403),
            .I(N__20370));
    InMux I__4727 (
            .O(N__20402),
            .I(N__20370));
    Span4Mux_h I__4726 (
            .O(N__20399),
            .I(N__20367));
    Odrv4 I__4725 (
            .O(N__20394),
            .I(\b2v_inst.indiceZ0Z_5 ));
    Odrv4 I__4724 (
            .O(N__20391),
            .I(\b2v_inst.indiceZ0Z_5 ));
    Odrv4 I__4723 (
            .O(N__20384),
            .I(\b2v_inst.indiceZ0Z_5 ));
    LocalMux I__4722 (
            .O(N__20375),
            .I(\b2v_inst.indiceZ0Z_5 ));
    LocalMux I__4721 (
            .O(N__20370),
            .I(\b2v_inst.indiceZ0Z_5 ));
    Odrv4 I__4720 (
            .O(N__20367),
            .I(\b2v_inst.indiceZ0Z_5 ));
    InMux I__4719 (
            .O(N__20354),
            .I(N__20351));
    LocalMux I__4718 (
            .O(N__20351),
            .I(N__20348));
    Span4Mux_h I__4717 (
            .O(N__20348),
            .I(N__20345));
    Span4Mux_h I__4716 (
            .O(N__20345),
            .I(N__20342));
    Odrv4 I__4715 (
            .O(N__20342),
            .I(\b2v_inst.dir_mem_2_RNO_1Z0Z_6 ));
    InMux I__4714 (
            .O(N__20339),
            .I(N__20336));
    LocalMux I__4713 (
            .O(N__20336),
            .I(\b2v_inst1.g0_i_o5_0_2 ));
    CascadeMux I__4712 (
            .O(N__20333),
            .I(N__20320));
    InMux I__4711 (
            .O(N__20332),
            .I(N__20317));
    InMux I__4710 (
            .O(N__20331),
            .I(N__20312));
    InMux I__4709 (
            .O(N__20330),
            .I(N__20312));
    CascadeMux I__4708 (
            .O(N__20329),
            .I(N__20309));
    InMux I__4707 (
            .O(N__20328),
            .I(N__20304));
    InMux I__4706 (
            .O(N__20327),
            .I(N__20304));
    InMux I__4705 (
            .O(N__20326),
            .I(N__20299));
    InMux I__4704 (
            .O(N__20325),
            .I(N__20299));
    CascadeMux I__4703 (
            .O(N__20324),
            .I(N__20291));
    InMux I__4702 (
            .O(N__20323),
            .I(N__20286));
    InMux I__4701 (
            .O(N__20320),
            .I(N__20286));
    LocalMux I__4700 (
            .O(N__20317),
            .I(N__20281));
    LocalMux I__4699 (
            .O(N__20312),
            .I(N__20281));
    InMux I__4698 (
            .O(N__20309),
            .I(N__20278));
    LocalMux I__4697 (
            .O(N__20304),
            .I(N__20271));
    LocalMux I__4696 (
            .O(N__20299),
            .I(N__20271));
    InMux I__4695 (
            .O(N__20298),
            .I(N__20266));
    InMux I__4694 (
            .O(N__20297),
            .I(N__20266));
    InMux I__4693 (
            .O(N__20296),
            .I(N__20257));
    InMux I__4692 (
            .O(N__20295),
            .I(N__20257));
    InMux I__4691 (
            .O(N__20294),
            .I(N__20257));
    InMux I__4690 (
            .O(N__20291),
            .I(N__20257));
    LocalMux I__4689 (
            .O(N__20286),
            .I(N__20254));
    Span4Mux_h I__4688 (
            .O(N__20281),
            .I(N__20249));
    LocalMux I__4687 (
            .O(N__20278),
            .I(N__20249));
    InMux I__4686 (
            .O(N__20277),
            .I(N__20246));
    CascadeMux I__4685 (
            .O(N__20276),
            .I(N__20243));
    Span4Mux_v I__4684 (
            .O(N__20271),
            .I(N__20239));
    LocalMux I__4683 (
            .O(N__20266),
            .I(N__20234));
    LocalMux I__4682 (
            .O(N__20257),
            .I(N__20234));
    Span4Mux_v I__4681 (
            .O(N__20254),
            .I(N__20227));
    Span4Mux_v I__4680 (
            .O(N__20249),
            .I(N__20227));
    LocalMux I__4679 (
            .O(N__20246),
            .I(N__20227));
    InMux I__4678 (
            .O(N__20243),
            .I(N__20222));
    InMux I__4677 (
            .O(N__20242),
            .I(N__20222));
    Odrv4 I__4676 (
            .O(N__20239),
            .I(\b2v_inst.indiceZ0Z_3 ));
    Odrv12 I__4675 (
            .O(N__20234),
            .I(\b2v_inst.indiceZ0Z_3 ));
    Odrv4 I__4674 (
            .O(N__20227),
            .I(\b2v_inst.indiceZ0Z_3 ));
    LocalMux I__4673 (
            .O(N__20222),
            .I(\b2v_inst.indiceZ0Z_3 ));
    CascadeMux I__4672 (
            .O(N__20213),
            .I(\b2v_inst.dir_mem_1_RNO_0Z0Z_3_cascade_ ));
    CascadeMux I__4671 (
            .O(N__20210),
            .I(N__20207));
    InMux I__4670 (
            .O(N__20207),
            .I(N__20204));
    LocalMux I__4669 (
            .O(N__20204),
            .I(N__20201));
    Odrv12 I__4668 (
            .O(N__20201),
            .I(\b2v_inst.dir_mem_1Z0Z_3 ));
    InMux I__4667 (
            .O(N__20198),
            .I(N__20195));
    LocalMux I__4666 (
            .O(N__20195),
            .I(\b2v_inst.indice_fast_RNIF91EZ0Z_0 ));
    InMux I__4665 (
            .O(N__20192),
            .I(N__20189));
    LocalMux I__4664 (
            .O(N__20189),
            .I(\b2v_inst.dir_mem_115lto8_1 ));
    InMux I__4663 (
            .O(N__20186),
            .I(N__20183));
    LocalMux I__4662 (
            .O(N__20183),
            .I(\b2v_inst.dir_mem_115lto6_1 ));
    InMux I__4661 (
            .O(N__20180),
            .I(N__20176));
    InMux I__4660 (
            .O(N__20179),
            .I(N__20173));
    LocalMux I__4659 (
            .O(N__20176),
            .I(\b2v_inst.un8_dir_mem_1_c7 ));
    LocalMux I__4658 (
            .O(N__20173),
            .I(\b2v_inst.un8_dir_mem_1_c7 ));
    CascadeMux I__4657 (
            .O(N__20168),
            .I(\b2v_inst.dir_mem_115lto8_1_cascade_ ));
    CascadeMux I__4656 (
            .O(N__20165),
            .I(\b2v_inst.dir_mem_115_0_cascade_ ));
    InMux I__4655 (
            .O(N__20162),
            .I(N__20159));
    LocalMux I__4654 (
            .O(N__20159),
            .I(N__20156));
    Span4Mux_v I__4653 (
            .O(N__20156),
            .I(N__20153));
    Span4Mux_h I__4652 (
            .O(N__20153),
            .I(N__20150));
    Odrv4 I__4651 (
            .O(N__20150),
            .I(\b2v_inst.dir_mem_1Z0Z_0 ));
    InMux I__4650 (
            .O(N__20147),
            .I(N__20143));
    CascadeMux I__4649 (
            .O(N__20146),
            .I(N__20136));
    LocalMux I__4648 (
            .O(N__20143),
            .I(N__20133));
    InMux I__4647 (
            .O(N__20142),
            .I(N__20128));
    InMux I__4646 (
            .O(N__20141),
            .I(N__20128));
    InMux I__4645 (
            .O(N__20140),
            .I(N__20125));
    InMux I__4644 (
            .O(N__20139),
            .I(N__20118));
    InMux I__4643 (
            .O(N__20136),
            .I(N__20118));
    Span4Mux_v I__4642 (
            .O(N__20133),
            .I(N__20110));
    LocalMux I__4641 (
            .O(N__20128),
            .I(N__20107));
    LocalMux I__4640 (
            .O(N__20125),
            .I(N__20103));
    InMux I__4639 (
            .O(N__20124),
            .I(N__20098));
    InMux I__4638 (
            .O(N__20123),
            .I(N__20098));
    LocalMux I__4637 (
            .O(N__20118),
            .I(N__20090));
    InMux I__4636 (
            .O(N__20117),
            .I(N__20085));
    InMux I__4635 (
            .O(N__20116),
            .I(N__20085));
    InMux I__4634 (
            .O(N__20115),
            .I(N__20082));
    InMux I__4633 (
            .O(N__20114),
            .I(N__20077));
    InMux I__4632 (
            .O(N__20113),
            .I(N__20077));
    Span4Mux_h I__4631 (
            .O(N__20110),
            .I(N__20072));
    Span4Mux_v I__4630 (
            .O(N__20107),
            .I(N__20072));
    InMux I__4629 (
            .O(N__20106),
            .I(N__20069));
    Span4Mux_h I__4628 (
            .O(N__20103),
            .I(N__20064));
    LocalMux I__4627 (
            .O(N__20098),
            .I(N__20064));
    InMux I__4626 (
            .O(N__20097),
            .I(N__20059));
    InMux I__4625 (
            .O(N__20096),
            .I(N__20059));
    InMux I__4624 (
            .O(N__20095),
            .I(N__20054));
    InMux I__4623 (
            .O(N__20094),
            .I(N__20054));
    InMux I__4622 (
            .O(N__20093),
            .I(N__20051));
    Span4Mux_h I__4621 (
            .O(N__20090),
            .I(N__20048));
    LocalMux I__4620 (
            .O(N__20085),
            .I(\b2v_inst.indiceZ0Z_2 ));
    LocalMux I__4619 (
            .O(N__20082),
            .I(\b2v_inst.indiceZ0Z_2 ));
    LocalMux I__4618 (
            .O(N__20077),
            .I(\b2v_inst.indiceZ0Z_2 ));
    Odrv4 I__4617 (
            .O(N__20072),
            .I(\b2v_inst.indiceZ0Z_2 ));
    LocalMux I__4616 (
            .O(N__20069),
            .I(\b2v_inst.indiceZ0Z_2 ));
    Odrv4 I__4615 (
            .O(N__20064),
            .I(\b2v_inst.indiceZ0Z_2 ));
    LocalMux I__4614 (
            .O(N__20059),
            .I(\b2v_inst.indiceZ0Z_2 ));
    LocalMux I__4613 (
            .O(N__20054),
            .I(\b2v_inst.indiceZ0Z_2 ));
    LocalMux I__4612 (
            .O(N__20051),
            .I(\b2v_inst.indiceZ0Z_2 ));
    Odrv4 I__4611 (
            .O(N__20048),
            .I(\b2v_inst.indiceZ0Z_2 ));
    CascadeMux I__4610 (
            .O(N__20027),
            .I(N__20024));
    InMux I__4609 (
            .O(N__20024),
            .I(N__20021));
    LocalMux I__4608 (
            .O(N__20021),
            .I(N__20016));
    InMux I__4607 (
            .O(N__20020),
            .I(N__20013));
    InMux I__4606 (
            .O(N__20019),
            .I(N__20010));
    Span4Mux_v I__4605 (
            .O(N__20016),
            .I(N__20007));
    LocalMux I__4604 (
            .O(N__20013),
            .I(\b2v_inst.un2_dir_mem_2_c2 ));
    LocalMux I__4603 (
            .O(N__20010),
            .I(\b2v_inst.un2_dir_mem_2_c2 ));
    Odrv4 I__4602 (
            .O(N__20007),
            .I(\b2v_inst.un2_dir_mem_2_c2 ));
    InMux I__4601 (
            .O(N__20000),
            .I(N__19997));
    LocalMux I__4600 (
            .O(N__19997),
            .I(N__19994));
    Span4Mux_v I__4599 (
            .O(N__19994),
            .I(N__19991));
    Span4Mux_h I__4598 (
            .O(N__19991),
            .I(N__19988));
    Odrv4 I__4597 (
            .O(N__19988),
            .I(\b2v_inst.dir_mem_1Z0Z_2 ));
    InMux I__4596 (
            .O(N__19985),
            .I(N__19982));
    LocalMux I__4595 (
            .O(N__19982),
            .I(\b2v_inst.dir_mem_1_RNO_0Z0Z_5 ));
    InMux I__4594 (
            .O(N__19979),
            .I(N__19976));
    LocalMux I__4593 (
            .O(N__19976),
            .I(N__19973));
    Span4Mux_h I__4592 (
            .O(N__19973),
            .I(N__19970));
    Span4Mux_h I__4591 (
            .O(N__19970),
            .I(N__19967));
    Odrv4 I__4590 (
            .O(N__19967),
            .I(\b2v_inst.dir_mem_1Z0Z_5 ));
    InMux I__4589 (
            .O(N__19964),
            .I(N__19952));
    InMux I__4588 (
            .O(N__19963),
            .I(N__19952));
    InMux I__4587 (
            .O(N__19962),
            .I(N__19952));
    InMux I__4586 (
            .O(N__19961),
            .I(N__19952));
    LocalMux I__4585 (
            .O(N__19952),
            .I(\b2v_inst.dir_mem_115_0 ));
    InMux I__4584 (
            .O(N__19949),
            .I(N__19946));
    LocalMux I__4583 (
            .O(N__19946),
            .I(N__19943));
    Span4Mux_h I__4582 (
            .O(N__19943),
            .I(N__19940));
    Span4Mux_h I__4581 (
            .O(N__19940),
            .I(N__19937));
    Odrv4 I__4580 (
            .O(N__19937),
            .I(\b2v_inst.dir_mem_1Z0Z_1 ));
    CEMux I__4579 (
            .O(N__19934),
            .I(N__19930));
    CEMux I__4578 (
            .O(N__19933),
            .I(N__19927));
    LocalMux I__4577 (
            .O(N__19930),
            .I(N__19921));
    LocalMux I__4576 (
            .O(N__19927),
            .I(N__19921));
    CEMux I__4575 (
            .O(N__19926),
            .I(N__19917));
    Span4Mux_v I__4574 (
            .O(N__19921),
            .I(N__19914));
    CEMux I__4573 (
            .O(N__19920),
            .I(N__19911));
    LocalMux I__4572 (
            .O(N__19917),
            .I(N__19908));
    Sp12to4 I__4571 (
            .O(N__19914),
            .I(N__19905));
    LocalMux I__4570 (
            .O(N__19911),
            .I(N__19900));
    Span4Mux_v I__4569 (
            .O(N__19908),
            .I(N__19900));
    Odrv12 I__4568 (
            .O(N__19905),
            .I(\b2v_inst.N_134_i ));
    Odrv4 I__4567 (
            .O(N__19900),
            .I(\b2v_inst.N_134_i ));
    InMux I__4566 (
            .O(N__19895),
            .I(N__19891));
    InMux I__4565 (
            .O(N__19894),
            .I(N__19886));
    LocalMux I__4564 (
            .O(N__19891),
            .I(N__19883));
    InMux I__4563 (
            .O(N__19890),
            .I(N__19880));
    CascadeMux I__4562 (
            .O(N__19889),
            .I(N__19877));
    LocalMux I__4561 (
            .O(N__19886),
            .I(N__19870));
    Span4Mux_h I__4560 (
            .O(N__19883),
            .I(N__19866));
    LocalMux I__4559 (
            .O(N__19880),
            .I(N__19863));
    InMux I__4558 (
            .O(N__19877),
            .I(N__19857));
    InMux I__4557 (
            .O(N__19876),
            .I(N__19857));
    InMux I__4556 (
            .O(N__19875),
            .I(N__19852));
    InMux I__4555 (
            .O(N__19874),
            .I(N__19852));
    InMux I__4554 (
            .O(N__19873),
            .I(N__19849));
    Span4Mux_h I__4553 (
            .O(N__19870),
            .I(N__19846));
    InMux I__4552 (
            .O(N__19869),
            .I(N__19843));
    Span4Mux_h I__4551 (
            .O(N__19866),
            .I(N__19838));
    Span4Mux_h I__4550 (
            .O(N__19863),
            .I(N__19838));
    InMux I__4549 (
            .O(N__19862),
            .I(N__19835));
    LocalMux I__4548 (
            .O(N__19857),
            .I(N__19830));
    LocalMux I__4547 (
            .O(N__19852),
            .I(N__19830));
    LocalMux I__4546 (
            .O(N__19849),
            .I(\b2v_inst.dir_memZ0Z_0 ));
    Odrv4 I__4545 (
            .O(N__19846),
            .I(\b2v_inst.dir_memZ0Z_0 ));
    LocalMux I__4544 (
            .O(N__19843),
            .I(\b2v_inst.dir_memZ0Z_0 ));
    Odrv4 I__4543 (
            .O(N__19838),
            .I(\b2v_inst.dir_memZ0Z_0 ));
    LocalMux I__4542 (
            .O(N__19835),
            .I(\b2v_inst.dir_memZ0Z_0 ));
    Odrv4 I__4541 (
            .O(N__19830),
            .I(\b2v_inst.dir_memZ0Z_0 ));
    InMux I__4540 (
            .O(N__19817),
            .I(N__19812));
    InMux I__4539 (
            .O(N__19816),
            .I(N__19809));
    InMux I__4538 (
            .O(N__19815),
            .I(N__19801));
    LocalMux I__4537 (
            .O(N__19812),
            .I(N__19798));
    LocalMux I__4536 (
            .O(N__19809),
            .I(N__19795));
    InMux I__4535 (
            .O(N__19808),
            .I(N__19792));
    InMux I__4534 (
            .O(N__19807),
            .I(N__19789));
    InMux I__4533 (
            .O(N__19806),
            .I(N__19786));
    InMux I__4532 (
            .O(N__19805),
            .I(N__19781));
    InMux I__4531 (
            .O(N__19804),
            .I(N__19781));
    LocalMux I__4530 (
            .O(N__19801),
            .I(N__19778));
    Span4Mux_h I__4529 (
            .O(N__19798),
            .I(N__19773));
    Span4Mux_h I__4528 (
            .O(N__19795),
            .I(N__19773));
    LocalMux I__4527 (
            .O(N__19792),
            .I(\b2v_inst.dir_memZ0Z_1 ));
    LocalMux I__4526 (
            .O(N__19789),
            .I(\b2v_inst.dir_memZ0Z_1 ));
    LocalMux I__4525 (
            .O(N__19786),
            .I(\b2v_inst.dir_memZ0Z_1 ));
    LocalMux I__4524 (
            .O(N__19781),
            .I(\b2v_inst.dir_memZ0Z_1 ));
    Odrv4 I__4523 (
            .O(N__19778),
            .I(\b2v_inst.dir_memZ0Z_1 ));
    Odrv4 I__4522 (
            .O(N__19773),
            .I(\b2v_inst.dir_memZ0Z_1 ));
    InMux I__4521 (
            .O(N__19760),
            .I(N__19751));
    InMux I__4520 (
            .O(N__19759),
            .I(N__19744));
    InMux I__4519 (
            .O(N__19758),
            .I(N__19744));
    InMux I__4518 (
            .O(N__19757),
            .I(N__19744));
    InMux I__4517 (
            .O(N__19756),
            .I(N__19741));
    InMux I__4516 (
            .O(N__19755),
            .I(N__19735));
    InMux I__4515 (
            .O(N__19754),
            .I(N__19735));
    LocalMux I__4514 (
            .O(N__19751),
            .I(N__19728));
    LocalMux I__4513 (
            .O(N__19744),
            .I(N__19728));
    LocalMux I__4512 (
            .O(N__19741),
            .I(N__19728));
    InMux I__4511 (
            .O(N__19740),
            .I(N__19718));
    LocalMux I__4510 (
            .O(N__19735),
            .I(N__19713));
    Span4Mux_v I__4509 (
            .O(N__19728),
            .I(N__19713));
    InMux I__4508 (
            .O(N__19727),
            .I(N__19708));
    InMux I__4507 (
            .O(N__19726),
            .I(N__19708));
    InMux I__4506 (
            .O(N__19725),
            .I(N__19703));
    InMux I__4505 (
            .O(N__19724),
            .I(N__19703));
    InMux I__4504 (
            .O(N__19723),
            .I(N__19696));
    InMux I__4503 (
            .O(N__19722),
            .I(N__19696));
    InMux I__4502 (
            .O(N__19721),
            .I(N__19696));
    LocalMux I__4501 (
            .O(N__19718),
            .I(\b2v_inst.N_253 ));
    Odrv4 I__4500 (
            .O(N__19713),
            .I(\b2v_inst.N_253 ));
    LocalMux I__4499 (
            .O(N__19708),
            .I(\b2v_inst.N_253 ));
    LocalMux I__4498 (
            .O(N__19703),
            .I(\b2v_inst.N_253 ));
    LocalMux I__4497 (
            .O(N__19696),
            .I(\b2v_inst.N_253 ));
    CascadeMux I__4496 (
            .O(N__19685),
            .I(N__19682));
    InMux I__4495 (
            .O(N__19682),
            .I(N__19679));
    LocalMux I__4494 (
            .O(N__19679),
            .I(N__19676));
    Odrv4 I__4493 (
            .O(N__19676),
            .I(\b2v_inst.un2_indice_21_s1_1 ));
    InMux I__4492 (
            .O(N__19673),
            .I(N__19668));
    InMux I__4491 (
            .O(N__19672),
            .I(N__19660));
    InMux I__4490 (
            .O(N__19671),
            .I(N__19660));
    LocalMux I__4489 (
            .O(N__19668),
            .I(N__19657));
    InMux I__4488 (
            .O(N__19667),
            .I(N__19652));
    InMux I__4487 (
            .O(N__19666),
            .I(N__19649));
    InMux I__4486 (
            .O(N__19665),
            .I(N__19646));
    LocalMux I__4485 (
            .O(N__19660),
            .I(N__19643));
    Span4Mux_h I__4484 (
            .O(N__19657),
            .I(N__19640));
    InMux I__4483 (
            .O(N__19656),
            .I(N__19637));
    InMux I__4482 (
            .O(N__19655),
            .I(N__19634));
    LocalMux I__4481 (
            .O(N__19652),
            .I(N__19631));
    LocalMux I__4480 (
            .O(N__19649),
            .I(\b2v_inst.un10_indice_2 ));
    LocalMux I__4479 (
            .O(N__19646),
            .I(\b2v_inst.un10_indice_2 ));
    Odrv4 I__4478 (
            .O(N__19643),
            .I(\b2v_inst.un10_indice_2 ));
    Odrv4 I__4477 (
            .O(N__19640),
            .I(\b2v_inst.un10_indice_2 ));
    LocalMux I__4476 (
            .O(N__19637),
            .I(\b2v_inst.un10_indice_2 ));
    LocalMux I__4475 (
            .O(N__19634),
            .I(\b2v_inst.un10_indice_2 ));
    Odrv4 I__4474 (
            .O(N__19631),
            .I(\b2v_inst.un10_indice_2 ));
    CascadeMux I__4473 (
            .O(N__19616),
            .I(N__19610));
    InMux I__4472 (
            .O(N__19615),
            .I(N__19607));
    CascadeMux I__4471 (
            .O(N__19614),
            .I(N__19604));
    InMux I__4470 (
            .O(N__19613),
            .I(N__19598));
    InMux I__4469 (
            .O(N__19610),
            .I(N__19598));
    LocalMux I__4468 (
            .O(N__19607),
            .I(N__19595));
    InMux I__4467 (
            .O(N__19604),
            .I(N__19592));
    InMux I__4466 (
            .O(N__19603),
            .I(N__19589));
    LocalMux I__4465 (
            .O(N__19598),
            .I(N__19584));
    Span4Mux_h I__4464 (
            .O(N__19595),
            .I(N__19581));
    LocalMux I__4463 (
            .O(N__19592),
            .I(N__19576));
    LocalMux I__4462 (
            .O(N__19589),
            .I(N__19576));
    InMux I__4461 (
            .O(N__19588),
            .I(N__19573));
    InMux I__4460 (
            .O(N__19587),
            .I(N__19570));
    Span4Mux_v I__4459 (
            .O(N__19584),
            .I(N__19563));
    Span4Mux_v I__4458 (
            .O(N__19581),
            .I(N__19563));
    Span4Mux_v I__4457 (
            .O(N__19576),
            .I(N__19563));
    LocalMux I__4456 (
            .O(N__19573),
            .I(\b2v_inst.CO1 ));
    LocalMux I__4455 (
            .O(N__19570),
            .I(\b2v_inst.CO1 ));
    Odrv4 I__4454 (
            .O(N__19563),
            .I(\b2v_inst.CO1 ));
    CascadeMux I__4453 (
            .O(N__19556),
            .I(\b2v_inst.CO1_cascade_ ));
    CascadeMux I__4452 (
            .O(N__19553),
            .I(\b2v_inst.un2_dir_mem_2_c2_cascade_ ));
    InMux I__4451 (
            .O(N__19550),
            .I(N__19541));
    InMux I__4450 (
            .O(N__19549),
            .I(N__19541));
    InMux I__4449 (
            .O(N__19548),
            .I(N__19541));
    LocalMux I__4448 (
            .O(N__19541),
            .I(\b2v_inst.indice_fastZ0Z_0 ));
    CascadeMux I__4447 (
            .O(N__19538),
            .I(N__19533));
    CascadeMux I__4446 (
            .O(N__19537),
            .I(N__19530));
    InMux I__4445 (
            .O(N__19536),
            .I(N__19523));
    InMux I__4444 (
            .O(N__19533),
            .I(N__19523));
    InMux I__4443 (
            .O(N__19530),
            .I(N__19523));
    LocalMux I__4442 (
            .O(N__19523),
            .I(\b2v_inst.indice_fastZ0Z_1 ));
    CascadeMux I__4441 (
            .O(N__19520),
            .I(N__19511));
    CascadeMux I__4440 (
            .O(N__19519),
            .I(N__19508));
    CascadeMux I__4439 (
            .O(N__19518),
            .I(N__19505));
    CascadeMux I__4438 (
            .O(N__19517),
            .I(N__19501));
    CascadeMux I__4437 (
            .O(N__19516),
            .I(N__19498));
    CascadeMux I__4436 (
            .O(N__19515),
            .I(N__19495));
    InMux I__4435 (
            .O(N__19514),
            .I(N__19492));
    InMux I__4434 (
            .O(N__19511),
            .I(N__19489));
    InMux I__4433 (
            .O(N__19508),
            .I(N__19486));
    InMux I__4432 (
            .O(N__19505),
            .I(N__19483));
    InMux I__4431 (
            .O(N__19504),
            .I(N__19478));
    InMux I__4430 (
            .O(N__19501),
            .I(N__19478));
    InMux I__4429 (
            .O(N__19498),
            .I(N__19473));
    InMux I__4428 (
            .O(N__19495),
            .I(N__19473));
    LocalMux I__4427 (
            .O(N__19492),
            .I(N__19469));
    LocalMux I__4426 (
            .O(N__19489),
            .I(N__19463));
    LocalMux I__4425 (
            .O(N__19486),
            .I(N__19460));
    LocalMux I__4424 (
            .O(N__19483),
            .I(N__19455));
    LocalMux I__4423 (
            .O(N__19478),
            .I(N__19455));
    LocalMux I__4422 (
            .O(N__19473),
            .I(N__19452));
    InMux I__4421 (
            .O(N__19472),
            .I(N__19449));
    Span4Mux_h I__4420 (
            .O(N__19469),
            .I(N__19446));
    InMux I__4419 (
            .O(N__19468),
            .I(N__19439));
    InMux I__4418 (
            .O(N__19467),
            .I(N__19439));
    InMux I__4417 (
            .O(N__19466),
            .I(N__19439));
    Span4Mux_v I__4416 (
            .O(N__19463),
            .I(N__19432));
    Span4Mux_v I__4415 (
            .O(N__19460),
            .I(N__19432));
    Span4Mux_h I__4414 (
            .O(N__19455),
            .I(N__19432));
    Span4Mux_h I__4413 (
            .O(N__19452),
            .I(N__19429));
    LocalMux I__4412 (
            .O(N__19449),
            .I(\b2v_inst.indice_2_repZ0Z1 ));
    Odrv4 I__4411 (
            .O(N__19446),
            .I(\b2v_inst.indice_2_repZ0Z1 ));
    LocalMux I__4410 (
            .O(N__19439),
            .I(\b2v_inst.indice_2_repZ0Z1 ));
    Odrv4 I__4409 (
            .O(N__19432),
            .I(\b2v_inst.indice_2_repZ0Z1 ));
    Odrv4 I__4408 (
            .O(N__19429),
            .I(\b2v_inst.indice_2_repZ0Z1 ));
    InMux I__4407 (
            .O(N__19418),
            .I(N__19412));
    InMux I__4406 (
            .O(N__19417),
            .I(N__19408));
    InMux I__4405 (
            .O(N__19416),
            .I(N__19405));
    InMux I__4404 (
            .O(N__19415),
            .I(N__19402));
    LocalMux I__4403 (
            .O(N__19412),
            .I(N__19399));
    InMux I__4402 (
            .O(N__19411),
            .I(N__19396));
    LocalMux I__4401 (
            .O(N__19408),
            .I(\b2v_inst1.m6_2 ));
    LocalMux I__4400 (
            .O(N__19405),
            .I(\b2v_inst1.m6_2 ));
    LocalMux I__4399 (
            .O(N__19402),
            .I(\b2v_inst1.m6_2 ));
    Odrv4 I__4398 (
            .O(N__19399),
            .I(\b2v_inst1.m6_2 ));
    LocalMux I__4397 (
            .O(N__19396),
            .I(\b2v_inst1.m6_2 ));
    CascadeMux I__4396 (
            .O(N__19385),
            .I(N__19382));
    InMux I__4395 (
            .O(N__19382),
            .I(N__19379));
    LocalMux I__4394 (
            .O(N__19379),
            .I(N__19376));
    Odrv4 I__4393 (
            .O(N__19376),
            .I(\b2v_inst.un2_indice_0_d1_c5 ));
    InMux I__4392 (
            .O(N__19373),
            .I(N__19369));
    InMux I__4391 (
            .O(N__19372),
            .I(N__19366));
    LocalMux I__4390 (
            .O(N__19369),
            .I(N__19363));
    LocalMux I__4389 (
            .O(N__19366),
            .I(N__19358));
    Span4Mux_v I__4388 (
            .O(N__19363),
            .I(N__19354));
    InMux I__4387 (
            .O(N__19362),
            .I(N__19351));
    InMux I__4386 (
            .O(N__19361),
            .I(N__19348));
    Span4Mux_h I__4385 (
            .O(N__19358),
            .I(N__19345));
    InMux I__4384 (
            .O(N__19357),
            .I(N__19342));
    Odrv4 I__4383 (
            .O(N__19354),
            .I(\b2v_inst.dir_memZ0Z_4 ));
    LocalMux I__4382 (
            .O(N__19351),
            .I(\b2v_inst.dir_memZ0Z_4 ));
    LocalMux I__4381 (
            .O(N__19348),
            .I(\b2v_inst.dir_memZ0Z_4 ));
    Odrv4 I__4380 (
            .O(N__19345),
            .I(\b2v_inst.dir_memZ0Z_4 ));
    LocalMux I__4379 (
            .O(N__19342),
            .I(\b2v_inst.dir_memZ0Z_4 ));
    CascadeMux I__4378 (
            .O(N__19331),
            .I(N__19328));
    InMux I__4377 (
            .O(N__19328),
            .I(N__19325));
    LocalMux I__4376 (
            .O(N__19325),
            .I(\b2v_inst.un2_indice_0_d1_ac0_7_s_0_0 ));
    InMux I__4375 (
            .O(N__19322),
            .I(N__19316));
    CascadeMux I__4374 (
            .O(N__19321),
            .I(N__19312));
    InMux I__4373 (
            .O(N__19320),
            .I(N__19309));
    InMux I__4372 (
            .O(N__19319),
            .I(N__19306));
    LocalMux I__4371 (
            .O(N__19316),
            .I(N__19303));
    InMux I__4370 (
            .O(N__19315),
            .I(N__19296));
    InMux I__4369 (
            .O(N__19312),
            .I(N__19296));
    LocalMux I__4368 (
            .O(N__19309),
            .I(N__19293));
    LocalMux I__4367 (
            .O(N__19306),
            .I(N__19290));
    Span4Mux_v I__4366 (
            .O(N__19303),
            .I(N__19287));
    InMux I__4365 (
            .O(N__19302),
            .I(N__19282));
    InMux I__4364 (
            .O(N__19301),
            .I(N__19282));
    LocalMux I__4363 (
            .O(N__19296),
            .I(N__19277));
    Span4Mux_v I__4362 (
            .O(N__19293),
            .I(N__19277));
    Span4Mux_h I__4361 (
            .O(N__19290),
            .I(N__19274));
    Odrv4 I__4360 (
            .O(N__19287),
            .I(\b2v_inst.dir_memZ0Z_3 ));
    LocalMux I__4359 (
            .O(N__19282),
            .I(\b2v_inst.dir_memZ0Z_3 ));
    Odrv4 I__4358 (
            .O(N__19277),
            .I(\b2v_inst.dir_memZ0Z_3 ));
    Odrv4 I__4357 (
            .O(N__19274),
            .I(\b2v_inst.dir_memZ0Z_3 ));
    InMux I__4356 (
            .O(N__19265),
            .I(N__19261));
    InMux I__4355 (
            .O(N__19264),
            .I(N__19257));
    LocalMux I__4354 (
            .O(N__19261),
            .I(N__19252));
    CascadeMux I__4353 (
            .O(N__19260),
            .I(N__19249));
    LocalMux I__4352 (
            .O(N__19257),
            .I(N__19246));
    InMux I__4351 (
            .O(N__19256),
            .I(N__19243));
    InMux I__4350 (
            .O(N__19255),
            .I(N__19240));
    Span4Mux_v I__4349 (
            .O(N__19252),
            .I(N__19237));
    InMux I__4348 (
            .O(N__19249),
            .I(N__19234));
    Span4Mux_h I__4347 (
            .O(N__19246),
            .I(N__19229));
    LocalMux I__4346 (
            .O(N__19243),
            .I(N__19229));
    LocalMux I__4345 (
            .O(N__19240),
            .I(\b2v_inst.dir_memZ0Z_5 ));
    Odrv4 I__4344 (
            .O(N__19237),
            .I(\b2v_inst.dir_memZ0Z_5 ));
    LocalMux I__4343 (
            .O(N__19234),
            .I(\b2v_inst.dir_memZ0Z_5 ));
    Odrv4 I__4342 (
            .O(N__19229),
            .I(\b2v_inst.dir_memZ0Z_5 ));
    CascadeMux I__4341 (
            .O(N__19220),
            .I(\b2v_inst.un2_indice_0_d1_ac0_7_s_0_0_cascade_ ));
    InMux I__4340 (
            .O(N__19217),
            .I(N__19214));
    LocalMux I__4339 (
            .O(N__19214),
            .I(N__19209));
    InMux I__4338 (
            .O(N__19213),
            .I(N__19206));
    CascadeMux I__4337 (
            .O(N__19212),
            .I(N__19202));
    Span4Mux_h I__4336 (
            .O(N__19209),
            .I(N__19195));
    LocalMux I__4335 (
            .O(N__19206),
            .I(N__19192));
    InMux I__4334 (
            .O(N__19205),
            .I(N__19189));
    InMux I__4333 (
            .O(N__19202),
            .I(N__19186));
    InMux I__4332 (
            .O(N__19201),
            .I(N__19181));
    InMux I__4331 (
            .O(N__19200),
            .I(N__19181));
    InMux I__4330 (
            .O(N__19199),
            .I(N__19176));
    InMux I__4329 (
            .O(N__19198),
            .I(N__19176));
    Span4Mux_v I__4328 (
            .O(N__19195),
            .I(N__19169));
    Span4Mux_v I__4327 (
            .O(N__19192),
            .I(N__19169));
    LocalMux I__4326 (
            .O(N__19189),
            .I(N__19169));
    LocalMux I__4325 (
            .O(N__19186),
            .I(\b2v_inst.dir_memZ0Z_2 ));
    LocalMux I__4324 (
            .O(N__19181),
            .I(\b2v_inst.dir_memZ0Z_2 ));
    LocalMux I__4323 (
            .O(N__19176),
            .I(\b2v_inst.dir_memZ0Z_2 ));
    Odrv4 I__4322 (
            .O(N__19169),
            .I(\b2v_inst.dir_memZ0Z_2 ));
    InMux I__4321 (
            .O(N__19160),
            .I(N__19156));
    CascadeMux I__4320 (
            .O(N__19159),
            .I(N__19153));
    LocalMux I__4319 (
            .O(N__19156),
            .I(N__19150));
    InMux I__4318 (
            .O(N__19153),
            .I(N__19146));
    Span4Mux_v I__4317 (
            .O(N__19150),
            .I(N__19143));
    InMux I__4316 (
            .O(N__19149),
            .I(N__19140));
    LocalMux I__4315 (
            .O(N__19146),
            .I(N__19137));
    Odrv4 I__4314 (
            .O(N__19143),
            .I(\b2v_inst.dir_memZ0Z_7 ));
    LocalMux I__4313 (
            .O(N__19140),
            .I(\b2v_inst.dir_memZ0Z_7 ));
    Odrv4 I__4312 (
            .O(N__19137),
            .I(\b2v_inst.dir_memZ0Z_7 ));
    CascadeMux I__4311 (
            .O(N__19130),
            .I(\b2v_inst.un2_indice_0_d1_ac0_9_0_cascade_ ));
    InMux I__4310 (
            .O(N__19127),
            .I(N__19123));
    InMux I__4309 (
            .O(N__19126),
            .I(N__19120));
    LocalMux I__4308 (
            .O(N__19123),
            .I(N__19116));
    LocalMux I__4307 (
            .O(N__19120),
            .I(N__19113));
    CascadeMux I__4306 (
            .O(N__19119),
            .I(N__19109));
    Span4Mux_v I__4305 (
            .O(N__19116),
            .I(N__19106));
    Span4Mux_h I__4304 (
            .O(N__19113),
            .I(N__19103));
    InMux I__4303 (
            .O(N__19112),
            .I(N__19098));
    InMux I__4302 (
            .O(N__19109),
            .I(N__19098));
    Odrv4 I__4301 (
            .O(N__19106),
            .I(\b2v_inst.dir_memZ0Z_6 ));
    Odrv4 I__4300 (
            .O(N__19103),
            .I(\b2v_inst.dir_memZ0Z_6 ));
    LocalMux I__4299 (
            .O(N__19098),
            .I(\b2v_inst.dir_memZ0Z_6 ));
    InMux I__4298 (
            .O(N__19091),
            .I(N__19088));
    LocalMux I__4297 (
            .O(N__19088),
            .I(N__19085));
    Odrv4 I__4296 (
            .O(N__19085),
            .I(\b2v_inst.un2_indice_21_s1_7 ));
    InMux I__4295 (
            .O(N__19082),
            .I(N__19077));
    InMux I__4294 (
            .O(N__19081),
            .I(N__19072));
    InMux I__4293 (
            .O(N__19080),
            .I(N__19067));
    LocalMux I__4292 (
            .O(N__19077),
            .I(N__19063));
    InMux I__4291 (
            .O(N__19076),
            .I(N__19059));
    InMux I__4290 (
            .O(N__19075),
            .I(N__19056));
    LocalMux I__4289 (
            .O(N__19072),
            .I(N__19053));
    InMux I__4288 (
            .O(N__19071),
            .I(N__19049));
    InMux I__4287 (
            .O(N__19070),
            .I(N__19045));
    LocalMux I__4286 (
            .O(N__19067),
            .I(N__19042));
    InMux I__4285 (
            .O(N__19066),
            .I(N__19039));
    Span4Mux_h I__4284 (
            .O(N__19063),
            .I(N__19036));
    InMux I__4283 (
            .O(N__19062),
            .I(N__19033));
    LocalMux I__4282 (
            .O(N__19059),
            .I(N__19026));
    LocalMux I__4281 (
            .O(N__19056),
            .I(N__19026));
    Span4Mux_v I__4280 (
            .O(N__19053),
            .I(N__19026));
    InMux I__4279 (
            .O(N__19052),
            .I(N__19023));
    LocalMux I__4278 (
            .O(N__19049),
            .I(N__19020));
    InMux I__4277 (
            .O(N__19048),
            .I(N__19017));
    LocalMux I__4276 (
            .O(N__19045),
            .I(\b2v_inst.state_17_repZ0Z1 ));
    Odrv4 I__4275 (
            .O(N__19042),
            .I(\b2v_inst.state_17_repZ0Z1 ));
    LocalMux I__4274 (
            .O(N__19039),
            .I(\b2v_inst.state_17_repZ0Z1 ));
    Odrv4 I__4273 (
            .O(N__19036),
            .I(\b2v_inst.state_17_repZ0Z1 ));
    LocalMux I__4272 (
            .O(N__19033),
            .I(\b2v_inst.state_17_repZ0Z1 ));
    Odrv4 I__4271 (
            .O(N__19026),
            .I(\b2v_inst.state_17_repZ0Z1 ));
    LocalMux I__4270 (
            .O(N__19023),
            .I(\b2v_inst.state_17_repZ0Z1 ));
    Odrv12 I__4269 (
            .O(N__19020),
            .I(\b2v_inst.state_17_repZ0Z1 ));
    LocalMux I__4268 (
            .O(N__19017),
            .I(\b2v_inst.state_17_repZ0Z1 ));
    InMux I__4267 (
            .O(N__18998),
            .I(N__18994));
    InMux I__4266 (
            .O(N__18997),
            .I(N__18991));
    LocalMux I__4265 (
            .O(N__18994),
            .I(N__18987));
    LocalMux I__4264 (
            .O(N__18991),
            .I(N__18978));
    InMux I__4263 (
            .O(N__18990),
            .I(N__18975));
    Span4Mux_v I__4262 (
            .O(N__18987),
            .I(N__18972));
    InMux I__4261 (
            .O(N__18986),
            .I(N__18969));
    InMux I__4260 (
            .O(N__18985),
            .I(N__18962));
    InMux I__4259 (
            .O(N__18984),
            .I(N__18962));
    InMux I__4258 (
            .O(N__18983),
            .I(N__18962));
    InMux I__4257 (
            .O(N__18982),
            .I(N__18957));
    InMux I__4256 (
            .O(N__18981),
            .I(N__18957));
    Span4Mux_v I__4255 (
            .O(N__18978),
            .I(N__18952));
    LocalMux I__4254 (
            .O(N__18975),
            .I(N__18952));
    Odrv4 I__4253 (
            .O(N__18972),
            .I(\b2v_inst.stateZ0Z_15 ));
    LocalMux I__4252 (
            .O(N__18969),
            .I(\b2v_inst.stateZ0Z_15 ));
    LocalMux I__4251 (
            .O(N__18962),
            .I(\b2v_inst.stateZ0Z_15 ));
    LocalMux I__4250 (
            .O(N__18957),
            .I(\b2v_inst.stateZ0Z_15 ));
    Odrv4 I__4249 (
            .O(N__18952),
            .I(\b2v_inst.stateZ0Z_15 ));
    CascadeMux I__4248 (
            .O(N__18941),
            .I(N__18934));
    CascadeMux I__4247 (
            .O(N__18940),
            .I(N__18928));
    CascadeMux I__4246 (
            .O(N__18939),
            .I(N__18924));
    InMux I__4245 (
            .O(N__18938),
            .I(N__18919));
    InMux I__4244 (
            .O(N__18937),
            .I(N__18911));
    InMux I__4243 (
            .O(N__18934),
            .I(N__18908));
    InMux I__4242 (
            .O(N__18933),
            .I(N__18905));
    InMux I__4241 (
            .O(N__18932),
            .I(N__18900));
    InMux I__4240 (
            .O(N__18931),
            .I(N__18900));
    InMux I__4239 (
            .O(N__18928),
            .I(N__18897));
    InMux I__4238 (
            .O(N__18927),
            .I(N__18892));
    InMux I__4237 (
            .O(N__18924),
            .I(N__18892));
    InMux I__4236 (
            .O(N__18923),
            .I(N__18887));
    InMux I__4235 (
            .O(N__18922),
            .I(N__18887));
    LocalMux I__4234 (
            .O(N__18919),
            .I(N__18884));
    InMux I__4233 (
            .O(N__18918),
            .I(N__18881));
    InMux I__4232 (
            .O(N__18917),
            .I(N__18876));
    InMux I__4231 (
            .O(N__18916),
            .I(N__18876));
    InMux I__4230 (
            .O(N__18915),
            .I(N__18873));
    InMux I__4229 (
            .O(N__18914),
            .I(N__18870));
    LocalMux I__4228 (
            .O(N__18911),
            .I(N__18867));
    LocalMux I__4227 (
            .O(N__18908),
            .I(N__18864));
    LocalMux I__4226 (
            .O(N__18905),
            .I(N__18860));
    LocalMux I__4225 (
            .O(N__18900),
            .I(N__18857));
    LocalMux I__4224 (
            .O(N__18897),
            .I(N__18854));
    LocalMux I__4223 (
            .O(N__18892),
            .I(N__18849));
    LocalMux I__4222 (
            .O(N__18887),
            .I(N__18849));
    Span4Mux_v I__4221 (
            .O(N__18884),
            .I(N__18842));
    LocalMux I__4220 (
            .O(N__18881),
            .I(N__18842));
    LocalMux I__4219 (
            .O(N__18876),
            .I(N__18842));
    LocalMux I__4218 (
            .O(N__18873),
            .I(N__18836));
    LocalMux I__4217 (
            .O(N__18870),
            .I(N__18836));
    Span4Mux_h I__4216 (
            .O(N__18867),
            .I(N__18831));
    Span4Mux_v I__4215 (
            .O(N__18864),
            .I(N__18831));
    InMux I__4214 (
            .O(N__18863),
            .I(N__18828));
    Span4Mux_h I__4213 (
            .O(N__18860),
            .I(N__18825));
    Span4Mux_v I__4212 (
            .O(N__18857),
            .I(N__18822));
    Span4Mux_v I__4211 (
            .O(N__18854),
            .I(N__18817));
    Span4Mux_v I__4210 (
            .O(N__18849),
            .I(N__18817));
    Span4Mux_v I__4209 (
            .O(N__18842),
            .I(N__18814));
    InMux I__4208 (
            .O(N__18841),
            .I(N__18811));
    Span4Mux_v I__4207 (
            .O(N__18836),
            .I(N__18808));
    Span4Mux_v I__4206 (
            .O(N__18831),
            .I(N__18803));
    LocalMux I__4205 (
            .O(N__18828),
            .I(N__18803));
    Sp12to4 I__4204 (
            .O(N__18825),
            .I(N__18800));
    Sp12to4 I__4203 (
            .O(N__18822),
            .I(N__18787));
    Sp12to4 I__4202 (
            .O(N__18817),
            .I(N__18787));
    Sp12to4 I__4201 (
            .O(N__18814),
            .I(N__18787));
    LocalMux I__4200 (
            .O(N__18811),
            .I(N__18787));
    Sp12to4 I__4199 (
            .O(N__18808),
            .I(N__18787));
    Sp12to4 I__4198 (
            .O(N__18803),
            .I(N__18787));
    Span12Mux_v I__4197 (
            .O(N__18800),
            .I(N__18782));
    Span12Mux_h I__4196 (
            .O(N__18787),
            .I(N__18782));
    Span12Mux_v I__4195 (
            .O(N__18782),
            .I(N__18779));
    Odrv12 I__4194 (
            .O(N__18779),
            .I(reset));
    InMux I__4193 (
            .O(N__18776),
            .I(N__18759));
    InMux I__4192 (
            .O(N__18775),
            .I(N__18756));
    InMux I__4191 (
            .O(N__18774),
            .I(N__18753));
    InMux I__4190 (
            .O(N__18773),
            .I(N__18750));
    InMux I__4189 (
            .O(N__18772),
            .I(N__18746));
    InMux I__4188 (
            .O(N__18771),
            .I(N__18742));
    InMux I__4187 (
            .O(N__18770),
            .I(N__18735));
    InMux I__4186 (
            .O(N__18769),
            .I(N__18735));
    InMux I__4185 (
            .O(N__18768),
            .I(N__18735));
    InMux I__4184 (
            .O(N__18767),
            .I(N__18730));
    InMux I__4183 (
            .O(N__18766),
            .I(N__18730));
    InMux I__4182 (
            .O(N__18765),
            .I(N__18727));
    InMux I__4181 (
            .O(N__18764),
            .I(N__18724));
    InMux I__4180 (
            .O(N__18763),
            .I(N__18719));
    InMux I__4179 (
            .O(N__18762),
            .I(N__18719));
    LocalMux I__4178 (
            .O(N__18759),
            .I(N__18716));
    LocalMux I__4177 (
            .O(N__18756),
            .I(N__18713));
    LocalMux I__4176 (
            .O(N__18753),
            .I(N__18710));
    LocalMux I__4175 (
            .O(N__18750),
            .I(N__18704));
    InMux I__4174 (
            .O(N__18749),
            .I(N__18700));
    LocalMux I__4173 (
            .O(N__18746),
            .I(N__18696));
    InMux I__4172 (
            .O(N__18745),
            .I(N__18693));
    LocalMux I__4171 (
            .O(N__18742),
            .I(N__18686));
    LocalMux I__4170 (
            .O(N__18735),
            .I(N__18686));
    LocalMux I__4169 (
            .O(N__18730),
            .I(N__18686));
    LocalMux I__4168 (
            .O(N__18727),
            .I(N__18683));
    LocalMux I__4167 (
            .O(N__18724),
            .I(N__18678));
    LocalMux I__4166 (
            .O(N__18719),
            .I(N__18678));
    Span4Mux_h I__4165 (
            .O(N__18716),
            .I(N__18675));
    Span4Mux_v I__4164 (
            .O(N__18713),
            .I(N__18670));
    Span4Mux_v I__4163 (
            .O(N__18710),
            .I(N__18670));
    InMux I__4162 (
            .O(N__18709),
            .I(N__18667));
    InMux I__4161 (
            .O(N__18708),
            .I(N__18662));
    InMux I__4160 (
            .O(N__18707),
            .I(N__18662));
    Span4Mux_h I__4159 (
            .O(N__18704),
            .I(N__18659));
    InMux I__4158 (
            .O(N__18703),
            .I(N__18656));
    LocalMux I__4157 (
            .O(N__18700),
            .I(N__18653));
    InMux I__4156 (
            .O(N__18699),
            .I(N__18650));
    Span4Mux_h I__4155 (
            .O(N__18696),
            .I(N__18639));
    LocalMux I__4154 (
            .O(N__18693),
            .I(N__18639));
    Span4Mux_v I__4153 (
            .O(N__18686),
            .I(N__18639));
    Span4Mux_h I__4152 (
            .O(N__18683),
            .I(N__18639));
    Span4Mux_v I__4151 (
            .O(N__18678),
            .I(N__18639));
    Odrv4 I__4150 (
            .O(N__18675),
            .I(\b2v_inst.N_351_0 ));
    Odrv4 I__4149 (
            .O(N__18670),
            .I(\b2v_inst.N_351_0 ));
    LocalMux I__4148 (
            .O(N__18667),
            .I(\b2v_inst.N_351_0 ));
    LocalMux I__4147 (
            .O(N__18662),
            .I(\b2v_inst.N_351_0 ));
    Odrv4 I__4146 (
            .O(N__18659),
            .I(\b2v_inst.N_351_0 ));
    LocalMux I__4145 (
            .O(N__18656),
            .I(\b2v_inst.N_351_0 ));
    Odrv4 I__4144 (
            .O(N__18653),
            .I(\b2v_inst.N_351_0 ));
    LocalMux I__4143 (
            .O(N__18650),
            .I(\b2v_inst.N_351_0 ));
    Odrv4 I__4142 (
            .O(N__18639),
            .I(\b2v_inst.N_351_0 ));
    SRMux I__4141 (
            .O(N__18620),
            .I(N__18617));
    LocalMux I__4140 (
            .O(N__18617),
            .I(N__18614));
    Span4Mux_v I__4139 (
            .O(N__18614),
            .I(N__18610));
    SRMux I__4138 (
            .O(N__18613),
            .I(N__18607));
    Span4Mux_v I__4137 (
            .O(N__18610),
            .I(N__18596));
    LocalMux I__4136 (
            .O(N__18607),
            .I(N__18596));
    CascadeMux I__4135 (
            .O(N__18606),
            .I(N__18593));
    CascadeMux I__4134 (
            .O(N__18605),
            .I(N__18590));
    CascadeMux I__4133 (
            .O(N__18604),
            .I(N__18587));
    CascadeMux I__4132 (
            .O(N__18603),
            .I(N__18584));
    CascadeMux I__4131 (
            .O(N__18602),
            .I(N__18581));
    CascadeMux I__4130 (
            .O(N__18601),
            .I(N__18578));
    Span4Mux_h I__4129 (
            .O(N__18596),
            .I(N__18575));
    InMux I__4128 (
            .O(N__18593),
            .I(N__18568));
    InMux I__4127 (
            .O(N__18590),
            .I(N__18568));
    InMux I__4126 (
            .O(N__18587),
            .I(N__18568));
    InMux I__4125 (
            .O(N__18584),
            .I(N__18561));
    InMux I__4124 (
            .O(N__18581),
            .I(N__18561));
    InMux I__4123 (
            .O(N__18578),
            .I(N__18561));
    Sp12to4 I__4122 (
            .O(N__18575),
            .I(N__18558));
    LocalMux I__4121 (
            .O(N__18568),
            .I(N__18553));
    LocalMux I__4120 (
            .O(N__18561),
            .I(N__18553));
    Span12Mux_v I__4119 (
            .O(N__18558),
            .I(N__18547));
    Span12Mux_s11_h I__4118 (
            .O(N__18553),
            .I(N__18547));
    InMux I__4117 (
            .O(N__18552),
            .I(N__18544));
    Odrv12 I__4116 (
            .O(N__18547),
            .I(CONSTANT_ONE_NET));
    LocalMux I__4115 (
            .O(N__18544),
            .I(CONSTANT_ONE_NET));
    CascadeMux I__4114 (
            .O(N__18539),
            .I(\b2v_inst.N_384_cascade_ ));
    InMux I__4113 (
            .O(N__18536),
            .I(N__18533));
    LocalMux I__4112 (
            .O(N__18533),
            .I(\b2v_inst.state_17_rep1_RNIN75CZ0Z3 ));
    InMux I__4111 (
            .O(N__18530),
            .I(N__18520));
    InMux I__4110 (
            .O(N__18529),
            .I(N__18520));
    InMux I__4109 (
            .O(N__18528),
            .I(N__18520));
    InMux I__4108 (
            .O(N__18527),
            .I(N__18517));
    LocalMux I__4107 (
            .O(N__18520),
            .I(\b2v_inst.un2_indice_3_0_iv_0_0_2 ));
    LocalMux I__4106 (
            .O(N__18517),
            .I(\b2v_inst.un2_indice_3_0_iv_0_0_2 ));
    CascadeMux I__4105 (
            .O(N__18512),
            .I(\b2v_inst1.m6_2_cascade_ ));
    InMux I__4104 (
            .O(N__18509),
            .I(N__18506));
    LocalMux I__4103 (
            .O(N__18506),
            .I(N__18503));
    Odrv4 I__4102 (
            .O(N__18503),
            .I(\b2v_inst1.N_10_0 ));
    InMux I__4101 (
            .O(N__18500),
            .I(N__18497));
    LocalMux I__4100 (
            .O(N__18497),
            .I(N__18494));
    Span4Mux_h I__4099 (
            .O(N__18494),
            .I(N__18491));
    Odrv4 I__4098 (
            .O(N__18491),
            .I(\b2v_inst1.g0_7_1 ));
    CascadeMux I__4097 (
            .O(N__18488),
            .I(\b2v_inst1.g0_i_1_cascade_ ));
    InMux I__4096 (
            .O(N__18485),
            .I(N__18482));
    LocalMux I__4095 (
            .O(N__18482),
            .I(N__18479));
    Odrv4 I__4094 (
            .O(N__18479),
            .I(\b2v_inst1.N_11_0 ));
    InMux I__4093 (
            .O(N__18476),
            .I(N__18473));
    LocalMux I__4092 (
            .O(N__18473),
            .I(N__18470));
    Odrv4 I__4091 (
            .O(N__18470),
            .I(\b2v_inst1.N_32_mux ));
    CascadeMux I__4090 (
            .O(N__18467),
            .I(\b2v_inst1.N_10_cascade_ ));
    CascadeMux I__4089 (
            .O(N__18464),
            .I(\b2v_inst1.g2_1_cascade_ ));
    InMux I__4088 (
            .O(N__18461),
            .I(N__18458));
    LocalMux I__4087 (
            .O(N__18458),
            .I(\b2v_inst1.g2_0 ));
    InMux I__4086 (
            .O(N__18455),
            .I(N__18452));
    LocalMux I__4085 (
            .O(N__18452),
            .I(\b2v_inst1.N_11_0_0 ));
    InMux I__4084 (
            .O(N__18449),
            .I(N__18445));
    InMux I__4083 (
            .O(N__18448),
            .I(N__18442));
    LocalMux I__4082 (
            .O(N__18445),
            .I(\b2v_inst1.N_9 ));
    LocalMux I__4081 (
            .O(N__18442),
            .I(\b2v_inst1.N_9 ));
    CascadeMux I__4080 (
            .O(N__18437),
            .I(\b2v_inst1.un1_r_Clk_Count_ac0_1_out_cascade_ ));
    InMux I__4079 (
            .O(N__18434),
            .I(N__18431));
    LocalMux I__4078 (
            .O(N__18431),
            .I(\b2v_inst1.m22_ns_1 ));
    CascadeMux I__4077 (
            .O(N__18428),
            .I(\b2v_inst1.N_29_mux_cascade_ ));
    CascadeMux I__4076 (
            .O(N__18425),
            .I(\b2v_inst1.N_11_cascade_ ));
    InMux I__4075 (
            .O(N__18422),
            .I(N__18419));
    LocalMux I__4074 (
            .O(N__18419),
            .I(N__18416));
    Odrv4 I__4073 (
            .O(N__18416),
            .I(\b2v_inst1.g0_0_i_1 ));
    InMux I__4072 (
            .O(N__18413),
            .I(N__18410));
    LocalMux I__4071 (
            .O(N__18410),
            .I(\b2v_inst1.N_14_0 ));
    CascadeMux I__4070 (
            .O(N__18407),
            .I(N__18404));
    InMux I__4069 (
            .O(N__18404),
            .I(N__18401));
    LocalMux I__4068 (
            .O(N__18401),
            .I(N__18398));
    Odrv4 I__4067 (
            .O(N__18398),
            .I(\b2v_inst1.g0_0_i_0 ));
    CascadeMux I__4066 (
            .O(N__18395),
            .I(N__18386));
    CascadeMux I__4065 (
            .O(N__18394),
            .I(N__18383));
    CascadeMux I__4064 (
            .O(N__18393),
            .I(N__18378));
    InMux I__4063 (
            .O(N__18392),
            .I(N__18375));
    InMux I__4062 (
            .O(N__18391),
            .I(N__18372));
    InMux I__4061 (
            .O(N__18390),
            .I(N__18367));
    InMux I__4060 (
            .O(N__18389),
            .I(N__18367));
    InMux I__4059 (
            .O(N__18386),
            .I(N__18364));
    InMux I__4058 (
            .O(N__18383),
            .I(N__18361));
    InMux I__4057 (
            .O(N__18382),
            .I(N__18356));
    InMux I__4056 (
            .O(N__18381),
            .I(N__18356));
    InMux I__4055 (
            .O(N__18378),
            .I(N__18353));
    LocalMux I__4054 (
            .O(N__18375),
            .I(\b2v_inst.indice_1_repZ0Z1 ));
    LocalMux I__4053 (
            .O(N__18372),
            .I(\b2v_inst.indice_1_repZ0Z1 ));
    LocalMux I__4052 (
            .O(N__18367),
            .I(\b2v_inst.indice_1_repZ0Z1 ));
    LocalMux I__4051 (
            .O(N__18364),
            .I(\b2v_inst.indice_1_repZ0Z1 ));
    LocalMux I__4050 (
            .O(N__18361),
            .I(\b2v_inst.indice_1_repZ0Z1 ));
    LocalMux I__4049 (
            .O(N__18356),
            .I(\b2v_inst.indice_1_repZ0Z1 ));
    LocalMux I__4048 (
            .O(N__18353),
            .I(\b2v_inst.indice_1_repZ0Z1 ));
    InMux I__4047 (
            .O(N__18338),
            .I(N__18333));
    InMux I__4046 (
            .O(N__18337),
            .I(N__18327));
    InMux I__4045 (
            .O(N__18336),
            .I(N__18324));
    LocalMux I__4044 (
            .O(N__18333),
            .I(N__18321));
    InMux I__4043 (
            .O(N__18332),
            .I(N__18316));
    InMux I__4042 (
            .O(N__18331),
            .I(N__18316));
    InMux I__4041 (
            .O(N__18330),
            .I(N__18313));
    LocalMux I__4040 (
            .O(N__18327),
            .I(\b2v_inst.indice_fastZ0Z_2 ));
    LocalMux I__4039 (
            .O(N__18324),
            .I(\b2v_inst.indice_fastZ0Z_2 ));
    Odrv4 I__4038 (
            .O(N__18321),
            .I(\b2v_inst.indice_fastZ0Z_2 ));
    LocalMux I__4037 (
            .O(N__18316),
            .I(\b2v_inst.indice_fastZ0Z_2 ));
    LocalMux I__4036 (
            .O(N__18313),
            .I(\b2v_inst.indice_fastZ0Z_2 ));
    CascadeMux I__4035 (
            .O(N__18302),
            .I(\b2v_inst.dir_mem_215lt6_0_cascade_ ));
    InMux I__4034 (
            .O(N__18299),
            .I(N__18296));
    LocalMux I__4033 (
            .O(N__18296),
            .I(N__18293));
    Span4Mux_h I__4032 (
            .O(N__18293),
            .I(N__18290));
    Odrv4 I__4031 (
            .O(N__18290),
            .I(\b2v_inst.dir_mem_215lt8 ));
    InMux I__4030 (
            .O(N__18287),
            .I(N__18284));
    LocalMux I__4029 (
            .O(N__18284),
            .I(N__18281));
    Odrv4 I__4028 (
            .O(N__18281),
            .I(\b2v_inst1.g0_0_i_a6_3_4 ));
    InMux I__4027 (
            .O(N__18278),
            .I(N__18275));
    LocalMux I__4026 (
            .O(N__18275),
            .I(N__18272));
    Span4Mux_v I__4025 (
            .O(N__18272),
            .I(N__18269));
    Span4Mux_h I__4024 (
            .O(N__18269),
            .I(N__18266));
    Odrv4 I__4023 (
            .O(N__18266),
            .I(\b2v_inst1.r_rx_byteZ0Z_7 ));
    CascadeMux I__4022 (
            .O(N__18263),
            .I(\b2v_inst1.r_rx_byteZ0Z_7_cascade_ ));
    InMux I__4021 (
            .O(N__18260),
            .I(N__18256));
    CascadeMux I__4020 (
            .O(N__18259),
            .I(N__18252));
    LocalMux I__4019 (
            .O(N__18256),
            .I(N__18248));
    InMux I__4018 (
            .O(N__18255),
            .I(N__18245));
    InMux I__4017 (
            .O(N__18252),
            .I(N__18240));
    InMux I__4016 (
            .O(N__18251),
            .I(N__18240));
    Span4Mux_h I__4015 (
            .O(N__18248),
            .I(N__18236));
    LocalMux I__4014 (
            .O(N__18245),
            .I(N__18231));
    LocalMux I__4013 (
            .O(N__18240),
            .I(N__18231));
    InMux I__4012 (
            .O(N__18239),
            .I(N__18228));
    Span4Mux_h I__4011 (
            .O(N__18236),
            .I(N__18221));
    Span4Mux_v I__4010 (
            .O(N__18231),
            .I(N__18218));
    LocalMux I__4009 (
            .O(N__18228),
            .I(N__18215));
    InMux I__4008 (
            .O(N__18227),
            .I(N__18210));
    InMux I__4007 (
            .O(N__18226),
            .I(N__18210));
    InMux I__4006 (
            .O(N__18225),
            .I(N__18205));
    InMux I__4005 (
            .O(N__18224),
            .I(N__18205));
    Odrv4 I__4004 (
            .O(N__18221),
            .I(\b2v_inst1.r_Bit_IndexZ0Z_2 ));
    Odrv4 I__4003 (
            .O(N__18218),
            .I(\b2v_inst1.r_Bit_IndexZ0Z_2 ));
    Odrv12 I__4002 (
            .O(N__18215),
            .I(\b2v_inst1.r_Bit_IndexZ0Z_2 ));
    LocalMux I__4001 (
            .O(N__18210),
            .I(\b2v_inst1.r_Bit_IndexZ0Z_2 ));
    LocalMux I__4000 (
            .O(N__18205),
            .I(\b2v_inst1.r_Bit_IndexZ0Z_2 ));
    CascadeMux I__3999 (
            .O(N__18194),
            .I(N__18188));
    InMux I__3998 (
            .O(N__18193),
            .I(N__18179));
    InMux I__3997 (
            .O(N__18192),
            .I(N__18179));
    InMux I__3996 (
            .O(N__18191),
            .I(N__18176));
    InMux I__3995 (
            .O(N__18188),
            .I(N__18169));
    InMux I__3994 (
            .O(N__18187),
            .I(N__18169));
    InMux I__3993 (
            .O(N__18186),
            .I(N__18169));
    CascadeMux I__3992 (
            .O(N__18185),
            .I(N__18166));
    InMux I__3991 (
            .O(N__18184),
            .I(N__18160));
    LocalMux I__3990 (
            .O(N__18179),
            .I(N__18153));
    LocalMux I__3989 (
            .O(N__18176),
            .I(N__18153));
    LocalMux I__3988 (
            .O(N__18169),
            .I(N__18153));
    InMux I__3987 (
            .O(N__18166),
            .I(N__18150));
    InMux I__3986 (
            .O(N__18165),
            .I(N__18147));
    InMux I__3985 (
            .O(N__18164),
            .I(N__18142));
    InMux I__3984 (
            .O(N__18163),
            .I(N__18142));
    LocalMux I__3983 (
            .O(N__18160),
            .I(N__18139));
    Span4Mux_h I__3982 (
            .O(N__18153),
            .I(N__18136));
    LocalMux I__3981 (
            .O(N__18150),
            .I(\b2v_inst1.r_Bit_IndexZ0Z_0 ));
    LocalMux I__3980 (
            .O(N__18147),
            .I(\b2v_inst1.r_Bit_IndexZ0Z_0 ));
    LocalMux I__3979 (
            .O(N__18142),
            .I(\b2v_inst1.r_Bit_IndexZ0Z_0 ));
    Odrv4 I__3978 (
            .O(N__18139),
            .I(\b2v_inst1.r_Bit_IndexZ0Z_0 ));
    Odrv4 I__3977 (
            .O(N__18136),
            .I(\b2v_inst1.r_Bit_IndexZ0Z_0 ));
    InMux I__3976 (
            .O(N__18125),
            .I(N__18120));
    InMux I__3975 (
            .O(N__18124),
            .I(N__18114));
    InMux I__3974 (
            .O(N__18123),
            .I(N__18114));
    LocalMux I__3973 (
            .O(N__18120),
            .I(N__18111));
    InMux I__3972 (
            .O(N__18119),
            .I(N__18108));
    LocalMux I__3971 (
            .O(N__18114),
            .I(N__18105));
    Span4Mux_h I__3970 (
            .O(N__18111),
            .I(N__18099));
    LocalMux I__3969 (
            .O(N__18108),
            .I(N__18094));
    Sp12to4 I__3968 (
            .O(N__18105),
            .I(N__18094));
    InMux I__3967 (
            .O(N__18104),
            .I(N__18091));
    InMux I__3966 (
            .O(N__18103),
            .I(N__18083));
    InMux I__3965 (
            .O(N__18102),
            .I(N__18083));
    Span4Mux_h I__3964 (
            .O(N__18099),
            .I(N__18080));
    Span12Mux_s10_v I__3963 (
            .O(N__18094),
            .I(N__18075));
    LocalMux I__3962 (
            .O(N__18091),
            .I(N__18075));
    InMux I__3961 (
            .O(N__18090),
            .I(N__18070));
    InMux I__3960 (
            .O(N__18089),
            .I(N__18070));
    InMux I__3959 (
            .O(N__18088),
            .I(N__18067));
    LocalMux I__3958 (
            .O(N__18083),
            .I(\b2v_inst1.r_Bit_IndexZ0Z_1 ));
    Odrv4 I__3957 (
            .O(N__18080),
            .I(\b2v_inst1.r_Bit_IndexZ0Z_1 ));
    Odrv12 I__3956 (
            .O(N__18075),
            .I(\b2v_inst1.r_Bit_IndexZ0Z_1 ));
    LocalMux I__3955 (
            .O(N__18070),
            .I(\b2v_inst1.r_Bit_IndexZ0Z_1 ));
    LocalMux I__3954 (
            .O(N__18067),
            .I(\b2v_inst1.r_Bit_IndexZ0Z_1 ));
    CascadeMux I__3953 (
            .O(N__18056),
            .I(\b2v_inst.un10_indice_2_cascade_ ));
    InMux I__3952 (
            .O(N__18053),
            .I(N__18050));
    LocalMux I__3951 (
            .O(N__18050),
            .I(\b2v_inst.indice_fast_RNIDAJGZ0Z_2 ));
    CascadeMux I__3950 (
            .O(N__18047),
            .I(\b2v_inst.dir_mem_115lto6_1_cascade_ ));
    CascadeMux I__3949 (
            .O(N__18044),
            .I(\b2v_inst.un1_dir_mem_1_mb_1_7_cascade_ ));
    InMux I__3948 (
            .O(N__18041),
            .I(N__18038));
    LocalMux I__3947 (
            .O(N__18038),
            .I(N__18035));
    Span4Mux_h I__3946 (
            .O(N__18035),
            .I(N__18032));
    Odrv4 I__3945 (
            .O(N__18032),
            .I(\b2v_inst.dir_mem_1Z0Z_7 ));
    InMux I__3944 (
            .O(N__18029),
            .I(N__18023));
    InMux I__3943 (
            .O(N__18028),
            .I(N__18020));
    InMux I__3942 (
            .O(N__18027),
            .I(N__18013));
    InMux I__3941 (
            .O(N__18026),
            .I(N__18013));
    LocalMux I__3940 (
            .O(N__18023),
            .I(N__18008));
    LocalMux I__3939 (
            .O(N__18020),
            .I(N__18008));
    CascadeMux I__3938 (
            .O(N__18019),
            .I(N__17999));
    InMux I__3937 (
            .O(N__18018),
            .I(N__17996));
    LocalMux I__3936 (
            .O(N__18013),
            .I(N__17991));
    Span4Mux_v I__3935 (
            .O(N__18008),
            .I(N__17991));
    InMux I__3934 (
            .O(N__18007),
            .I(N__17984));
    InMux I__3933 (
            .O(N__18006),
            .I(N__17984));
    InMux I__3932 (
            .O(N__18005),
            .I(N__17984));
    InMux I__3931 (
            .O(N__18004),
            .I(N__17975));
    InMux I__3930 (
            .O(N__18003),
            .I(N__17975));
    InMux I__3929 (
            .O(N__18002),
            .I(N__17975));
    InMux I__3928 (
            .O(N__17999),
            .I(N__17975));
    LocalMux I__3927 (
            .O(N__17996),
            .I(N__17970));
    Span4Mux_h I__3926 (
            .O(N__17991),
            .I(N__17963));
    LocalMux I__3925 (
            .O(N__17984),
            .I(N__17963));
    LocalMux I__3924 (
            .O(N__17975),
            .I(N__17963));
    CascadeMux I__3923 (
            .O(N__17974),
            .I(N__17959));
    CascadeMux I__3922 (
            .O(N__17973),
            .I(N__17955));
    Span4Mux_v I__3921 (
            .O(N__17970),
            .I(N__17952));
    Span4Mux_v I__3920 (
            .O(N__17963),
            .I(N__17949));
    InMux I__3919 (
            .O(N__17962),
            .I(N__17946));
    InMux I__3918 (
            .O(N__17959),
            .I(N__17939));
    InMux I__3917 (
            .O(N__17958),
            .I(N__17939));
    InMux I__3916 (
            .O(N__17955),
            .I(N__17939));
    Odrv4 I__3915 (
            .O(N__17952),
            .I(\b2v_inst.indiceZ0Z_4 ));
    Odrv4 I__3914 (
            .O(N__17949),
            .I(\b2v_inst.indiceZ0Z_4 ));
    LocalMux I__3913 (
            .O(N__17946),
            .I(\b2v_inst.indiceZ0Z_4 ));
    LocalMux I__3912 (
            .O(N__17939),
            .I(\b2v_inst.indiceZ0Z_4 ));
    CascadeMux I__3911 (
            .O(N__17930),
            .I(N__17927));
    InMux I__3910 (
            .O(N__17927),
            .I(N__17924));
    LocalMux I__3909 (
            .O(N__17924),
            .I(N__17921));
    Span4Mux_h I__3908 (
            .O(N__17921),
            .I(N__17918));
    Odrv4 I__3907 (
            .O(N__17918),
            .I(\b2v_inst.un2_dir_mem_2_c5 ));
    CascadeMux I__3906 (
            .O(N__17915),
            .I(\b2v_inst.N_4_0_0_cascade_ ));
    InMux I__3905 (
            .O(N__17912),
            .I(N__17909));
    LocalMux I__3904 (
            .O(N__17909),
            .I(N__17906));
    Odrv4 I__3903 (
            .O(N__17906),
            .I(\b2v_inst.N_8_0 ));
    CascadeMux I__3902 (
            .O(N__17903),
            .I(\b2v_inst.dir_mem_315lto8_a0_1_cascade_ ));
    CascadeMux I__3901 (
            .O(N__17900),
            .I(N__17897));
    InMux I__3900 (
            .O(N__17897),
            .I(N__17894));
    LocalMux I__3899 (
            .O(N__17894),
            .I(N__17891));
    Span4Mux_v I__3898 (
            .O(N__17891),
            .I(N__17888));
    Span4Mux_h I__3897 (
            .O(N__17888),
            .I(N__17885));
    Odrv4 I__3896 (
            .O(N__17885),
            .I(\b2v_inst.indice_fast_RNIRFV61Z0Z_3 ));
    InMux I__3895 (
            .O(N__17882),
            .I(N__17879));
    LocalMux I__3894 (
            .O(N__17879),
            .I(N__17876));
    Span4Mux_h I__3893 (
            .O(N__17876),
            .I(N__17865));
    InMux I__3892 (
            .O(N__17875),
            .I(N__17858));
    InMux I__3891 (
            .O(N__17874),
            .I(N__17858));
    InMux I__3890 (
            .O(N__17873),
            .I(N__17858));
    InMux I__3889 (
            .O(N__17872),
            .I(N__17853));
    InMux I__3888 (
            .O(N__17871),
            .I(N__17853));
    InMux I__3887 (
            .O(N__17870),
            .I(N__17848));
    InMux I__3886 (
            .O(N__17869),
            .I(N__17848));
    InMux I__3885 (
            .O(N__17868),
            .I(N__17845));
    Odrv4 I__3884 (
            .O(N__17865),
            .I(\b2v_inst.indice_0_repZ0Z1 ));
    LocalMux I__3883 (
            .O(N__17858),
            .I(\b2v_inst.indice_0_repZ0Z1 ));
    LocalMux I__3882 (
            .O(N__17853),
            .I(\b2v_inst.indice_0_repZ0Z1 ));
    LocalMux I__3881 (
            .O(N__17848),
            .I(\b2v_inst.indice_0_repZ0Z1 ));
    LocalMux I__3880 (
            .O(N__17845),
            .I(\b2v_inst.indice_0_repZ0Z1 ));
    InMux I__3879 (
            .O(N__17834),
            .I(N__17831));
    LocalMux I__3878 (
            .O(N__17831),
            .I(\b2v_inst.indice_0_rep1_RNIFJJGZ0 ));
    InMux I__3877 (
            .O(N__17828),
            .I(N__17825));
    LocalMux I__3876 (
            .O(N__17825),
            .I(N__17820));
    InMux I__3875 (
            .O(N__17824),
            .I(N__17815));
    InMux I__3874 (
            .O(N__17823),
            .I(N__17815));
    Span4Mux_v I__3873 (
            .O(N__17820),
            .I(N__17810));
    LocalMux I__3872 (
            .O(N__17815),
            .I(N__17810));
    Span4Mux_h I__3871 (
            .O(N__17810),
            .I(N__17807));
    Odrv4 I__3870 (
            .O(N__17807),
            .I(\b2v_inst.N_410 ));
    InMux I__3869 (
            .O(N__17804),
            .I(N__17801));
    LocalMux I__3868 (
            .O(N__17801),
            .I(\b2v_inst.un2_indice_3_iv_0_0_1 ));
    InMux I__3867 (
            .O(N__17798),
            .I(N__17795));
    LocalMux I__3866 (
            .O(N__17795),
            .I(N__17787));
    CascadeMux I__3865 (
            .O(N__17794),
            .I(N__17783));
    CascadeMux I__3864 (
            .O(N__17793),
            .I(N__17777));
    CascadeMux I__3863 (
            .O(N__17792),
            .I(N__17774));
    CascadeMux I__3862 (
            .O(N__17791),
            .I(N__17770));
    CascadeMux I__3861 (
            .O(N__17790),
            .I(N__17765));
    Span4Mux_h I__3860 (
            .O(N__17787),
            .I(N__17761));
    InMux I__3859 (
            .O(N__17786),
            .I(N__17756));
    InMux I__3858 (
            .O(N__17783),
            .I(N__17756));
    InMux I__3857 (
            .O(N__17782),
            .I(N__17753));
    InMux I__3856 (
            .O(N__17781),
            .I(N__17742));
    InMux I__3855 (
            .O(N__17780),
            .I(N__17742));
    InMux I__3854 (
            .O(N__17777),
            .I(N__17742));
    InMux I__3853 (
            .O(N__17774),
            .I(N__17742));
    InMux I__3852 (
            .O(N__17773),
            .I(N__17742));
    InMux I__3851 (
            .O(N__17770),
            .I(N__17737));
    InMux I__3850 (
            .O(N__17769),
            .I(N__17737));
    InMux I__3849 (
            .O(N__17768),
            .I(N__17730));
    InMux I__3848 (
            .O(N__17765),
            .I(N__17730));
    InMux I__3847 (
            .O(N__17764),
            .I(N__17730));
    Odrv4 I__3846 (
            .O(N__17761),
            .I(\b2v_inst.N_253_i ));
    LocalMux I__3845 (
            .O(N__17756),
            .I(\b2v_inst.N_253_i ));
    LocalMux I__3844 (
            .O(N__17753),
            .I(\b2v_inst.N_253_i ));
    LocalMux I__3843 (
            .O(N__17742),
            .I(\b2v_inst.N_253_i ));
    LocalMux I__3842 (
            .O(N__17737),
            .I(\b2v_inst.N_253_i ));
    LocalMux I__3841 (
            .O(N__17730),
            .I(\b2v_inst.N_253_i ));
    InMux I__3840 (
            .O(N__17717),
            .I(N__17707));
    InMux I__3839 (
            .O(N__17716),
            .I(N__17707));
    InMux I__3838 (
            .O(N__17715),
            .I(N__17707));
    InMux I__3837 (
            .O(N__17714),
            .I(N__17704));
    LocalMux I__3836 (
            .O(N__17707),
            .I(N__17693));
    LocalMux I__3835 (
            .O(N__17704),
            .I(N__17693));
    InMux I__3834 (
            .O(N__17703),
            .I(N__17687));
    InMux I__3833 (
            .O(N__17702),
            .I(N__17687));
    CascadeMux I__3832 (
            .O(N__17701),
            .I(N__17684));
    CascadeMux I__3831 (
            .O(N__17700),
            .I(N__17680));
    InMux I__3830 (
            .O(N__17699),
            .I(N__17676));
    InMux I__3829 (
            .O(N__17698),
            .I(N__17673));
    Span4Mux_v I__3828 (
            .O(N__17693),
            .I(N__17670));
    CascadeMux I__3827 (
            .O(N__17692),
            .I(N__17663));
    LocalMux I__3826 (
            .O(N__17687),
            .I(N__17660));
    InMux I__3825 (
            .O(N__17684),
            .I(N__17657));
    InMux I__3824 (
            .O(N__17683),
            .I(N__17654));
    InMux I__3823 (
            .O(N__17680),
            .I(N__17651));
    InMux I__3822 (
            .O(N__17679),
            .I(N__17648));
    LocalMux I__3821 (
            .O(N__17676),
            .I(N__17645));
    LocalMux I__3820 (
            .O(N__17673),
            .I(N__17640));
    Span4Mux_h I__3819 (
            .O(N__17670),
            .I(N__17640));
    InMux I__3818 (
            .O(N__17669),
            .I(N__17636));
    InMux I__3817 (
            .O(N__17668),
            .I(N__17633));
    InMux I__3816 (
            .O(N__17667),
            .I(N__17628));
    InMux I__3815 (
            .O(N__17666),
            .I(N__17628));
    InMux I__3814 (
            .O(N__17663),
            .I(N__17625));
    Span4Mux_h I__3813 (
            .O(N__17660),
            .I(N__17622));
    LocalMux I__3812 (
            .O(N__17657),
            .I(N__17613));
    LocalMux I__3811 (
            .O(N__17654),
            .I(N__17613));
    LocalMux I__3810 (
            .O(N__17651),
            .I(N__17613));
    LocalMux I__3809 (
            .O(N__17648),
            .I(N__17613));
    Span4Mux_h I__3808 (
            .O(N__17645),
            .I(N__17608));
    Span4Mux_v I__3807 (
            .O(N__17640),
            .I(N__17608));
    InMux I__3806 (
            .O(N__17639),
            .I(N__17605));
    LocalMux I__3805 (
            .O(N__17636),
            .I(\b2v_inst.stateZ0Z_17 ));
    LocalMux I__3804 (
            .O(N__17633),
            .I(\b2v_inst.stateZ0Z_17 ));
    LocalMux I__3803 (
            .O(N__17628),
            .I(\b2v_inst.stateZ0Z_17 ));
    LocalMux I__3802 (
            .O(N__17625),
            .I(\b2v_inst.stateZ0Z_17 ));
    Odrv4 I__3801 (
            .O(N__17622),
            .I(\b2v_inst.stateZ0Z_17 ));
    Odrv12 I__3800 (
            .O(N__17613),
            .I(\b2v_inst.stateZ0Z_17 ));
    Odrv4 I__3799 (
            .O(N__17608),
            .I(\b2v_inst.stateZ0Z_17 ));
    LocalMux I__3798 (
            .O(N__17605),
            .I(\b2v_inst.stateZ0Z_17 ));
    CascadeMux I__3797 (
            .O(N__17588),
            .I(\b2v_inst.un2_indice_20_0_cascade_ ));
    InMux I__3796 (
            .O(N__17585),
            .I(N__17582));
    LocalMux I__3795 (
            .O(N__17582),
            .I(N__17579));
    Span4Mux_v I__3794 (
            .O(N__17579),
            .I(N__17576));
    Odrv4 I__3793 (
            .O(N__17576),
            .I(\b2v_inst.N_4_0 ));
    InMux I__3792 (
            .O(N__17573),
            .I(N__17569));
    CascadeMux I__3791 (
            .O(N__17572),
            .I(N__17566));
    LocalMux I__3790 (
            .O(N__17569),
            .I(N__17563));
    InMux I__3789 (
            .O(N__17566),
            .I(N__17560));
    Span4Mux_h I__3788 (
            .O(N__17563),
            .I(N__17557));
    LocalMux I__3787 (
            .O(N__17560),
            .I(\b2v_inst.un2_cuentalto7_3 ));
    Odrv4 I__3786 (
            .O(N__17557),
            .I(\b2v_inst.un2_cuentalto7_3 ));
    CascadeMux I__3785 (
            .O(N__17552),
            .I(\b2v_inst.N_228_cascade_ ));
    InMux I__3784 (
            .O(N__17549),
            .I(N__17546));
    LocalMux I__3783 (
            .O(N__17546),
            .I(N__17543));
    Span4Mux_h I__3782 (
            .O(N__17543),
            .I(N__17540));
    Odrv4 I__3781 (
            .O(N__17540),
            .I(\b2v_inst.cuenta_RNI925FZ0Z_7 ));
    InMux I__3780 (
            .O(N__17537),
            .I(N__17527));
    InMux I__3779 (
            .O(N__17536),
            .I(N__17527));
    InMux I__3778 (
            .O(N__17535),
            .I(N__17527));
    InMux I__3777 (
            .O(N__17534),
            .I(N__17522));
    LocalMux I__3776 (
            .O(N__17527),
            .I(N__17519));
    InMux I__3775 (
            .O(N__17526),
            .I(N__17514));
    InMux I__3774 (
            .O(N__17525),
            .I(N__17514));
    LocalMux I__3773 (
            .O(N__17522),
            .I(\b2v_inst.N_234 ));
    Odrv4 I__3772 (
            .O(N__17519),
            .I(\b2v_inst.N_234 ));
    LocalMux I__3771 (
            .O(N__17514),
            .I(\b2v_inst.N_234 ));
    InMux I__3770 (
            .O(N__17507),
            .I(N__17503));
    InMux I__3769 (
            .O(N__17506),
            .I(N__17500));
    LocalMux I__3768 (
            .O(N__17503),
            .I(\b2v_inst.un2_indice_3_0_iv_0_a2_0_8_2_2 ));
    LocalMux I__3767 (
            .O(N__17500),
            .I(\b2v_inst.un2_indice_3_0_iv_0_a2_0_8_2_2 ));
    InMux I__3766 (
            .O(N__17495),
            .I(N__17492));
    LocalMux I__3765 (
            .O(N__17492),
            .I(\b2v_inst.N_228 ));
    CascadeMux I__3764 (
            .O(N__17489),
            .I(\b2v_inst.N_383_8_cascade_ ));
    InMux I__3763 (
            .O(N__17486),
            .I(N__17483));
    LocalMux I__3762 (
            .O(N__17483),
            .I(N__17479));
    InMux I__3761 (
            .O(N__17482),
            .I(N__17476));
    Odrv4 I__3760 (
            .O(N__17479),
            .I(\b2v_inst.un2_indice_3_0_iv_0_a2_0_8_3_2 ));
    LocalMux I__3759 (
            .O(N__17476),
            .I(\b2v_inst.un2_indice_3_0_iv_0_a2_0_8_3_2 ));
    CascadeMux I__3758 (
            .O(N__17471),
            .I(N__17468));
    InMux I__3757 (
            .O(N__17468),
            .I(N__17464));
    CascadeMux I__3756 (
            .O(N__17467),
            .I(N__17461));
    LocalMux I__3755 (
            .O(N__17464),
            .I(N__17458));
    InMux I__3754 (
            .O(N__17461),
            .I(N__17455));
    Span4Mux_v I__3753 (
            .O(N__17458),
            .I(N__17452));
    LocalMux I__3752 (
            .O(N__17455),
            .I(N__17449));
    Odrv4 I__3751 (
            .O(N__17452),
            .I(\b2v_inst.un2_indice_21_s0_2 ));
    Odrv4 I__3750 (
            .O(N__17449),
            .I(\b2v_inst.un2_indice_21_s0_2 ));
    InMux I__3749 (
            .O(N__17444),
            .I(N__17441));
    LocalMux I__3748 (
            .O(N__17441),
            .I(\b2v_inst.un2_indice_20_2 ));
    InMux I__3747 (
            .O(N__17438),
            .I(N__17435));
    LocalMux I__3746 (
            .O(N__17435),
            .I(\b2v_inst.un2_indice_21_s1_2 ));
    CascadeMux I__3745 (
            .O(N__17432),
            .I(\b2v_inst.un2_indice_3_0_iv_0_1_2_cascade_ ));
    CascadeMux I__3744 (
            .O(N__17429),
            .I(N__17426));
    InMux I__3743 (
            .O(N__17426),
            .I(N__17423));
    LocalMux I__3742 (
            .O(N__17423),
            .I(N__17420));
    Odrv4 I__3741 (
            .O(N__17420),
            .I(\b2v_inst.dir_mem_RNO_3Z0Z_4 ));
    InMux I__3740 (
            .O(N__17417),
            .I(N__17414));
    LocalMux I__3739 (
            .O(N__17414),
            .I(\b2v_inst.un2_indice_0_d1_c2 ));
    InMux I__3738 (
            .O(N__17411),
            .I(N__17404));
    InMux I__3737 (
            .O(N__17410),
            .I(N__17404));
    InMux I__3736 (
            .O(N__17409),
            .I(N__17401));
    LocalMux I__3735 (
            .O(N__17404),
            .I(N__17395));
    LocalMux I__3734 (
            .O(N__17401),
            .I(N__17392));
    InMux I__3733 (
            .O(N__17400),
            .I(N__17387));
    InMux I__3732 (
            .O(N__17399),
            .I(N__17384));
    CascadeMux I__3731 (
            .O(N__17398),
            .I(N__17381));
    Span4Mux_v I__3730 (
            .O(N__17395),
            .I(N__17377));
    Span12Mux_h I__3729 (
            .O(N__17392),
            .I(N__17374));
    InMux I__3728 (
            .O(N__17391),
            .I(N__17371));
    InMux I__3727 (
            .O(N__17390),
            .I(N__17368));
    LocalMux I__3726 (
            .O(N__17387),
            .I(N__17363));
    LocalMux I__3725 (
            .O(N__17384),
            .I(N__17363));
    InMux I__3724 (
            .O(N__17381),
            .I(N__17360));
    InMux I__3723 (
            .O(N__17380),
            .I(N__17357));
    Odrv4 I__3722 (
            .O(N__17377),
            .I(\b2v_inst.N_451 ));
    Odrv12 I__3721 (
            .O(N__17374),
            .I(\b2v_inst.N_451 ));
    LocalMux I__3720 (
            .O(N__17371),
            .I(\b2v_inst.N_451 ));
    LocalMux I__3719 (
            .O(N__17368),
            .I(\b2v_inst.N_451 ));
    Odrv4 I__3718 (
            .O(N__17363),
            .I(\b2v_inst.N_451 ));
    LocalMux I__3717 (
            .O(N__17360),
            .I(\b2v_inst.N_451 ));
    LocalMux I__3716 (
            .O(N__17357),
            .I(\b2v_inst.N_451 ));
    CascadeMux I__3715 (
            .O(N__17342),
            .I(N__17338));
    InMux I__3714 (
            .O(N__17341),
            .I(N__17335));
    InMux I__3713 (
            .O(N__17338),
            .I(N__17332));
    LocalMux I__3712 (
            .O(N__17335),
            .I(\b2v_inst.un2_indice_21_s0_3 ));
    LocalMux I__3711 (
            .O(N__17332),
            .I(\b2v_inst.un2_indice_21_s0_3 ));
    InMux I__3710 (
            .O(N__17327),
            .I(N__17324));
    LocalMux I__3709 (
            .O(N__17324),
            .I(N__17321));
    Odrv4 I__3708 (
            .O(N__17321),
            .I(\b2v_inst.un2_indice_20_3 ));
    InMux I__3707 (
            .O(N__17318),
            .I(N__17315));
    LocalMux I__3706 (
            .O(N__17315),
            .I(\b2v_inst.un2_indice_21_s1_3 ));
    CascadeMux I__3705 (
            .O(N__17312),
            .I(\b2v_inst.un2_indice_3_0_iv_0_0_3_cascade_ ));
    InMux I__3704 (
            .O(N__17309),
            .I(N__17306));
    LocalMux I__3703 (
            .O(N__17306),
            .I(\b2v_inst.dir_mem_RNO_5Z0Z_4 ));
    InMux I__3702 (
            .O(N__17303),
            .I(N__17300));
    LocalMux I__3701 (
            .O(N__17300),
            .I(\b2v_inst.un2_indice_3_iv_0_1_0_5 ));
    CascadeMux I__3700 (
            .O(N__17297),
            .I(\b2v_inst1.g0_0_i_a6_2_2_cascade_ ));
    InMux I__3699 (
            .O(N__17294),
            .I(N__17291));
    LocalMux I__3698 (
            .O(N__17291),
            .I(\b2v_inst1.g0_0_i_a6_2_1 ));
    InMux I__3697 (
            .O(N__17288),
            .I(N__17285));
    LocalMux I__3696 (
            .O(N__17285),
            .I(\b2v_inst1.N_18 ));
    InMux I__3695 (
            .O(N__17282),
            .I(N__17279));
    LocalMux I__3694 (
            .O(N__17279),
            .I(N__17276));
    Span4Mux_v I__3693 (
            .O(N__17276),
            .I(N__17273));
    Odrv4 I__3692 (
            .O(N__17273),
            .I(\b2v_inst.dir_mem_RNO_2Z0Z_4 ));
    CascadeMux I__3691 (
            .O(N__17270),
            .I(\b2v_inst.un2_indice_3_0_i_1_4_cascade_ ));
    InMux I__3690 (
            .O(N__17267),
            .I(N__17264));
    LocalMux I__3689 (
            .O(N__17264),
            .I(N__17261));
    Odrv4 I__3688 (
            .O(N__17261),
            .I(\b2v_inst.un2_indice_20_4 ));
    CascadeMux I__3687 (
            .O(N__17258),
            .I(N__17255));
    InMux I__3686 (
            .O(N__17255),
            .I(N__17252));
    LocalMux I__3685 (
            .O(N__17252),
            .I(N__17249));
    Odrv4 I__3684 (
            .O(N__17249),
            .I(\b2v_inst.dir_mem_RNO_2Z0Z_7 ));
    InMux I__3683 (
            .O(N__17246),
            .I(N__17243));
    LocalMux I__3682 (
            .O(N__17243),
            .I(\b2v_inst.un2_indice_20_7 ));
    CascadeMux I__3681 (
            .O(N__17240),
            .I(\b2v_inst.un2_indice_3_0_iv_0_0_7_cascade_ ));
    CascadeMux I__3680 (
            .O(N__17237),
            .I(\b2v_inst1.N_7_cascade_ ));
    InMux I__3679 (
            .O(N__17234),
            .I(N__17231));
    LocalMux I__3678 (
            .O(N__17231),
            .I(\b2v_inst1.g0_0_i_a6_1_2 ));
    CascadeMux I__3677 (
            .O(N__17228),
            .I(\b2v_inst1.N_9_cascade_ ));
    InMux I__3676 (
            .O(N__17225),
            .I(N__17222));
    LocalMux I__3675 (
            .O(N__17222),
            .I(N__17219));
    Odrv12 I__3674 (
            .O(N__17219),
            .I(\b2v_inst1.g0_0_i_a6_3_5 ));
    CascadeMux I__3673 (
            .O(N__17216),
            .I(\b2v_inst1.N_19_cascade_ ));
    InMux I__3672 (
            .O(N__17213),
            .I(N__17210));
    LocalMux I__3671 (
            .O(N__17210),
            .I(N__17207));
    Odrv4 I__3670 (
            .O(N__17207),
            .I(\b2v_inst1.N_6 ));
    InMux I__3669 (
            .O(N__17204),
            .I(N__17201));
    LocalMux I__3668 (
            .O(N__17201),
            .I(\b2v_inst1.r_SM_Main_1_sqmuxa_1_0 ));
    CascadeMux I__3667 (
            .O(N__17198),
            .I(N__17195));
    InMux I__3666 (
            .O(N__17195),
            .I(N__17192));
    LocalMux I__3665 (
            .O(N__17192),
            .I(\b2v_inst1.g0_3_4 ));
    InMux I__3664 (
            .O(N__17189),
            .I(N__17186));
    LocalMux I__3663 (
            .O(N__17186),
            .I(N__17183));
    Span4Mux_h I__3662 (
            .O(N__17183),
            .I(N__17180));
    Odrv4 I__3661 (
            .O(N__17180),
            .I(\b2v_inst1.r_RX_Bytece_0_2 ));
    InMux I__3660 (
            .O(N__17177),
            .I(N__17167));
    InMux I__3659 (
            .O(N__17176),
            .I(N__17154));
    InMux I__3658 (
            .O(N__17175),
            .I(N__17154));
    InMux I__3657 (
            .O(N__17174),
            .I(N__17154));
    InMux I__3656 (
            .O(N__17173),
            .I(N__17154));
    InMux I__3655 (
            .O(N__17172),
            .I(N__17154));
    InMux I__3654 (
            .O(N__17171),
            .I(N__17154));
    InMux I__3653 (
            .O(N__17170),
            .I(N__17151));
    LocalMux I__3652 (
            .O(N__17167),
            .I(N__17148));
    LocalMux I__3651 (
            .O(N__17154),
            .I(N__17145));
    LocalMux I__3650 (
            .O(N__17151),
            .I(N__17142));
    Span4Mux_h I__3649 (
            .O(N__17148),
            .I(N__17139));
    Span4Mux_h I__3648 (
            .O(N__17145),
            .I(N__17136));
    Span4Mux_v I__3647 (
            .O(N__17142),
            .I(N__17133));
    Odrv4 I__3646 (
            .O(N__17139),
            .I(\b2v_inst1.r_RX_Byte_1_sqmuxa ));
    Odrv4 I__3645 (
            .O(N__17136),
            .I(\b2v_inst1.r_RX_Byte_1_sqmuxa ));
    Odrv4 I__3644 (
            .O(N__17133),
            .I(\b2v_inst1.r_RX_Byte_1_sqmuxa ));
    InMux I__3643 (
            .O(N__17126),
            .I(N__17123));
    LocalMux I__3642 (
            .O(N__17123),
            .I(N__17120));
    Odrv12 I__3641 (
            .O(N__17120),
            .I(\b2v_inst1.r_RX_Bytece_0_0_0 ));
    CascadeMux I__3640 (
            .O(N__17117),
            .I(N__17109));
    InMux I__3639 (
            .O(N__17116),
            .I(N__17105));
    InMux I__3638 (
            .O(N__17115),
            .I(N__17102));
    InMux I__3637 (
            .O(N__17114),
            .I(N__17099));
    InMux I__3636 (
            .O(N__17113),
            .I(N__17094));
    InMux I__3635 (
            .O(N__17112),
            .I(N__17094));
    InMux I__3634 (
            .O(N__17109),
            .I(N__17089));
    InMux I__3633 (
            .O(N__17108),
            .I(N__17089));
    LocalMux I__3632 (
            .O(N__17105),
            .I(N__17084));
    LocalMux I__3631 (
            .O(N__17102),
            .I(N__17081));
    LocalMux I__3630 (
            .O(N__17099),
            .I(N__17074));
    LocalMux I__3629 (
            .O(N__17094),
            .I(N__17074));
    LocalMux I__3628 (
            .O(N__17089),
            .I(N__17074));
    InMux I__3627 (
            .O(N__17088),
            .I(N__17069));
    InMux I__3626 (
            .O(N__17087),
            .I(N__17069));
    Odrv4 I__3625 (
            .O(N__17084),
            .I(\b2v_inst.indice_3_repZ0Z1 ));
    Odrv4 I__3624 (
            .O(N__17081),
            .I(\b2v_inst.indice_3_repZ0Z1 ));
    Odrv12 I__3623 (
            .O(N__17074),
            .I(\b2v_inst.indice_3_repZ0Z1 ));
    LocalMux I__3622 (
            .O(N__17069),
            .I(\b2v_inst.indice_3_repZ0Z1 ));
    CascadeMux I__3621 (
            .O(N__17060),
            .I(N__17057));
    InMux I__3620 (
            .O(N__17057),
            .I(N__17054));
    LocalMux I__3619 (
            .O(N__17054),
            .I(N__17051));
    Odrv4 I__3618 (
            .O(N__17051),
            .I(\b2v_inst.un2_dir_mem_2_c4_d ));
    CascadeMux I__3617 (
            .O(N__17048),
            .I(\b2v_inst.dir_mem_RNO_4Z0Z_4_cascade_ ));
    InMux I__3616 (
            .O(N__17045),
            .I(N__17042));
    LocalMux I__3615 (
            .O(N__17042),
            .I(N__17039));
    Span4Mux_h I__3614 (
            .O(N__17039),
            .I(N__17036));
    Odrv4 I__3613 (
            .O(N__17036),
            .I(\b2v_inst.indice_RNIA33NZ0Z_1 ));
    InMux I__3612 (
            .O(N__17033),
            .I(N__17021));
    InMux I__3611 (
            .O(N__17032),
            .I(N__17021));
    InMux I__3610 (
            .O(N__17031),
            .I(N__17021));
    InMux I__3609 (
            .O(N__17030),
            .I(N__17021));
    LocalMux I__3608 (
            .O(N__17021),
            .I(N__17014));
    InMux I__3607 (
            .O(N__17020),
            .I(N__17004));
    InMux I__3606 (
            .O(N__17019),
            .I(N__17004));
    InMux I__3605 (
            .O(N__17018),
            .I(N__17004));
    InMux I__3604 (
            .O(N__17017),
            .I(N__17001));
    Span4Mux_v I__3603 (
            .O(N__17014),
            .I(N__16997));
    InMux I__3602 (
            .O(N__17013),
            .I(N__16994));
    InMux I__3601 (
            .O(N__17012),
            .I(N__16991));
    InMux I__3600 (
            .O(N__17011),
            .I(N__16988));
    LocalMux I__3599 (
            .O(N__17004),
            .I(N__16985));
    LocalMux I__3598 (
            .O(N__17001),
            .I(N__16982));
    InMux I__3597 (
            .O(N__17000),
            .I(N__16979));
    Span4Mux_h I__3596 (
            .O(N__16997),
            .I(N__16976));
    LocalMux I__3595 (
            .O(N__16994),
            .I(N__16969));
    LocalMux I__3594 (
            .O(N__16991),
            .I(N__16969));
    LocalMux I__3593 (
            .O(N__16988),
            .I(N__16969));
    Odrv4 I__3592 (
            .O(N__16985),
            .I(\b2v_inst.N_238 ));
    Odrv4 I__3591 (
            .O(N__16982),
            .I(\b2v_inst.N_238 ));
    LocalMux I__3590 (
            .O(N__16979),
            .I(\b2v_inst.N_238 ));
    Odrv4 I__3589 (
            .O(N__16976),
            .I(\b2v_inst.N_238 ));
    Odrv12 I__3588 (
            .O(N__16969),
            .I(\b2v_inst.N_238 ));
    InMux I__3587 (
            .O(N__16958),
            .I(N__16954));
    InMux I__3586 (
            .O(N__16957),
            .I(N__16947));
    LocalMux I__3585 (
            .O(N__16954),
            .I(N__16943));
    InMux I__3584 (
            .O(N__16953),
            .I(N__16940));
    InMux I__3583 (
            .O(N__16952),
            .I(N__16937));
    InMux I__3582 (
            .O(N__16951),
            .I(N__16930));
    InMux I__3581 (
            .O(N__16950),
            .I(N__16930));
    LocalMux I__3580 (
            .O(N__16947),
            .I(N__16927));
    InMux I__3579 (
            .O(N__16946),
            .I(N__16924));
    Span4Mux_v I__3578 (
            .O(N__16943),
            .I(N__16921));
    LocalMux I__3577 (
            .O(N__16940),
            .I(N__16916));
    LocalMux I__3576 (
            .O(N__16937),
            .I(N__16916));
    InMux I__3575 (
            .O(N__16936),
            .I(N__16911));
    InMux I__3574 (
            .O(N__16935),
            .I(N__16911));
    LocalMux I__3573 (
            .O(N__16930),
            .I(N__16906));
    Span4Mux_h I__3572 (
            .O(N__16927),
            .I(N__16906));
    LocalMux I__3571 (
            .O(N__16924),
            .I(\b2v_inst.N_236 ));
    Odrv4 I__3570 (
            .O(N__16921),
            .I(\b2v_inst.N_236 ));
    Odrv4 I__3569 (
            .O(N__16916),
            .I(\b2v_inst.N_236 ));
    LocalMux I__3568 (
            .O(N__16911),
            .I(\b2v_inst.N_236 ));
    Odrv4 I__3567 (
            .O(N__16906),
            .I(\b2v_inst.N_236 ));
    CascadeMux I__3566 (
            .O(N__16895),
            .I(N__16892));
    InMux I__3565 (
            .O(N__16892),
            .I(N__16889));
    LocalMux I__3564 (
            .O(N__16889),
            .I(N__16886));
    Span4Mux_h I__3563 (
            .O(N__16886),
            .I(N__16883));
    Odrv4 I__3562 (
            .O(N__16883),
            .I(\b2v_inst.dir_mem_3Z0Z_2 ));
    InMux I__3561 (
            .O(N__16880),
            .I(N__16877));
    LocalMux I__3560 (
            .O(N__16877),
            .I(N__16874));
    Odrv12 I__3559 (
            .O(N__16874),
            .I(\b2v_inst.addr_ram_1_0_iv_i_1_2 ));
    CascadeMux I__3558 (
            .O(N__16871),
            .I(\b2v_inst.un10_indice_cascade_ ));
    InMux I__3557 (
            .O(N__16868),
            .I(N__16865));
    LocalMux I__3556 (
            .O(N__16865),
            .I(\b2v_inst.un2_indice_3_iv_0_a2_2_sx_5 ));
    CascadeMux I__3555 (
            .O(N__16862),
            .I(N__16859));
    InMux I__3554 (
            .O(N__16859),
            .I(N__16856));
    LocalMux I__3553 (
            .O(N__16856),
            .I(N__16852));
    InMux I__3552 (
            .O(N__16855),
            .I(N__16849));
    Odrv4 I__3551 (
            .O(N__16852),
            .I(\b2v_inst.un2_indice_0_d0_c4_d ));
    LocalMux I__3550 (
            .O(N__16849),
            .I(\b2v_inst.un2_indice_0_d0_c4_d ));
    CascadeMux I__3549 (
            .O(N__16844),
            .I(\b2v_inst.un2_m1_e_0_cascade_ ));
    CascadeMux I__3548 (
            .O(N__16841),
            .I(N__16838));
    InMux I__3547 (
            .O(N__16838),
            .I(N__16835));
    LocalMux I__3546 (
            .O(N__16835),
            .I(N__16832));
    Odrv4 I__3545 (
            .O(N__16832),
            .I(\b2v_inst.dir_mem_RNIR93H1Z0Z_5 ));
    CascadeMux I__3544 (
            .O(N__16829),
            .I(N__16826));
    InMux I__3543 (
            .O(N__16826),
            .I(N__16823));
    LocalMux I__3542 (
            .O(N__16823),
            .I(N__16820));
    Span4Mux_h I__3541 (
            .O(N__16820),
            .I(N__16817));
    Odrv4 I__3540 (
            .O(N__16817),
            .I(\b2v_inst.g1_0_3 ));
    InMux I__3539 (
            .O(N__16814),
            .I(N__16811));
    LocalMux I__3538 (
            .O(N__16811),
            .I(\b2v_inst.g0_2_7 ));
    InMux I__3537 (
            .O(N__16808),
            .I(N__16805));
    LocalMux I__3536 (
            .O(N__16805),
            .I(N__16800));
    InMux I__3535 (
            .O(N__16804),
            .I(N__16797));
    InMux I__3534 (
            .O(N__16803),
            .I(N__16794));
    Odrv4 I__3533 (
            .O(N__16800),
            .I(\b2v_inst.N_467 ));
    LocalMux I__3532 (
            .O(N__16797),
            .I(\b2v_inst.N_467 ));
    LocalMux I__3531 (
            .O(N__16794),
            .I(\b2v_inst.N_467 ));
    CascadeMux I__3530 (
            .O(N__16787),
            .I(\b2v_inst.N_411_cascade_ ));
    InMux I__3529 (
            .O(N__16784),
            .I(N__16781));
    LocalMux I__3528 (
            .O(N__16781),
            .I(N__16778));
    Odrv4 I__3527 (
            .O(N__16778),
            .I(\b2v_inst.un2_indice_20_5 ));
    InMux I__3526 (
            .O(N__16775),
            .I(\b2v_inst.un2_indice_cry_6 ));
    CascadeMux I__3525 (
            .O(N__16772),
            .I(\b2v_inst.un2_indice_21_s0_1_cascade_ ));
    CascadeMux I__3524 (
            .O(N__16769),
            .I(N__16766));
    InMux I__3523 (
            .O(N__16766),
            .I(N__16763));
    LocalMux I__3522 (
            .O(N__16763),
            .I(\b2v_inst.un2_indice_21_s0_1 ));
    InMux I__3521 (
            .O(N__16760),
            .I(N__16757));
    LocalMux I__3520 (
            .O(N__16757),
            .I(\b2v_inst.un2_indice_20_1 ));
    InMux I__3519 (
            .O(N__16754),
            .I(N__16751));
    LocalMux I__3518 (
            .O(N__16751),
            .I(\b2v_inst.dir_mem_RNO_2Z0Z_1 ));
    CascadeMux I__3517 (
            .O(N__16748),
            .I(\b2v_inst.dir_mem_RNO_3Z0Z_1_cascade_ ));
    CascadeMux I__3516 (
            .O(N__16745),
            .I(N__16742));
    InMux I__3515 (
            .O(N__16742),
            .I(N__16739));
    LocalMux I__3514 (
            .O(N__16739),
            .I(N__16736));
    Odrv4 I__3513 (
            .O(N__16736),
            .I(\b2v_inst.dir_mem_RNIP73H1Z0Z_4 ));
    InMux I__3512 (
            .O(N__16733),
            .I(N__16729));
    InMux I__3511 (
            .O(N__16732),
            .I(N__16726));
    LocalMux I__3510 (
            .O(N__16729),
            .I(N__16719));
    LocalMux I__3509 (
            .O(N__16726),
            .I(N__16716));
    InMux I__3508 (
            .O(N__16725),
            .I(N__16713));
    InMux I__3507 (
            .O(N__16724),
            .I(N__16706));
    InMux I__3506 (
            .O(N__16723),
            .I(N__16706));
    InMux I__3505 (
            .O(N__16722),
            .I(N__16706));
    Odrv4 I__3504 (
            .O(N__16719),
            .I(\b2v_inst.dir_mem_215_0 ));
    Odrv4 I__3503 (
            .O(N__16716),
            .I(\b2v_inst.dir_mem_215_0 ));
    LocalMux I__3502 (
            .O(N__16713),
            .I(\b2v_inst.dir_mem_215_0 ));
    LocalMux I__3501 (
            .O(N__16706),
            .I(\b2v_inst.dir_mem_215_0 ));
    CascadeMux I__3500 (
            .O(N__16697),
            .I(N__16694));
    InMux I__3499 (
            .O(N__16694),
            .I(N__16691));
    LocalMux I__3498 (
            .O(N__16691),
            .I(N__16688));
    Span4Mux_v I__3497 (
            .O(N__16688),
            .I(N__16685));
    Odrv4 I__3496 (
            .O(N__16685),
            .I(\b2v_inst.dir_mem_2Z0Z_5 ));
    CEMux I__3495 (
            .O(N__16682),
            .I(N__16679));
    LocalMux I__3494 (
            .O(N__16679),
            .I(N__16674));
    CEMux I__3493 (
            .O(N__16678),
            .I(N__16670));
    CEMux I__3492 (
            .O(N__16677),
            .I(N__16667));
    Span4Mux_v I__3491 (
            .O(N__16674),
            .I(N__16664));
    CEMux I__3490 (
            .O(N__16673),
            .I(N__16661));
    LocalMux I__3489 (
            .O(N__16670),
            .I(N__16656));
    LocalMux I__3488 (
            .O(N__16667),
            .I(N__16656));
    Span4Mux_h I__3487 (
            .O(N__16664),
            .I(N__16651));
    LocalMux I__3486 (
            .O(N__16661),
            .I(N__16651));
    Span4Mux_v I__3485 (
            .O(N__16656),
            .I(N__16648));
    Span4Mux_h I__3484 (
            .O(N__16651),
            .I(N__16645));
    Span4Mux_h I__3483 (
            .O(N__16648),
            .I(N__16642));
    Span4Mux_h I__3482 (
            .O(N__16645),
            .I(N__16639));
    Odrv4 I__3481 (
            .O(N__16642),
            .I(\b2v_inst.N_136_i ));
    Odrv4 I__3480 (
            .O(N__16639),
            .I(\b2v_inst.N_136_i ));
    InMux I__3479 (
            .O(N__16634),
            .I(N__16628));
    InMux I__3478 (
            .O(N__16633),
            .I(N__16628));
    LocalMux I__3477 (
            .O(N__16628),
            .I(\b2v_inst1.N_14 ));
    CascadeMux I__3476 (
            .O(N__16625),
            .I(N__16622));
    InMux I__3475 (
            .O(N__16622),
            .I(N__16619));
    LocalMux I__3474 (
            .O(N__16619),
            .I(\b2v_inst.dir_mem_RNIGVEE1Z0Z_0 ));
    InMux I__3473 (
            .O(N__16616),
            .I(N__16613));
    LocalMux I__3472 (
            .O(N__16613),
            .I(\b2v_inst.dir_mem_RNII5PO1Z0Z_1 ));
    InMux I__3471 (
            .O(N__16610),
            .I(\b2v_inst.un2_indice_cry_0 ));
    InMux I__3470 (
            .O(N__16607),
            .I(N__16604));
    LocalMux I__3469 (
            .O(N__16604),
            .I(\b2v_inst.dir_mem_RNIL33H1Z0Z_2 ));
    InMux I__3468 (
            .O(N__16601),
            .I(\b2v_inst.un2_indice_cry_1 ));
    InMux I__3467 (
            .O(N__16598),
            .I(N__16595));
    LocalMux I__3466 (
            .O(N__16595),
            .I(\b2v_inst.dir_mem_RNIN53H1Z0Z_3 ));
    InMux I__3465 (
            .O(N__16592),
            .I(\b2v_inst.un2_indice_cry_2 ));
    InMux I__3464 (
            .O(N__16589),
            .I(\b2v_inst.un2_indice_cry_3 ));
    InMux I__3463 (
            .O(N__16586),
            .I(\b2v_inst.un2_indice_cry_4 ));
    CascadeMux I__3462 (
            .O(N__16583),
            .I(N__16580));
    InMux I__3461 (
            .O(N__16580),
            .I(N__16577));
    LocalMux I__3460 (
            .O(N__16577),
            .I(\b2v_inst.dir_mem_RNITB3H1Z0Z_6 ));
    InMux I__3459 (
            .O(N__16574),
            .I(N__16571));
    LocalMux I__3458 (
            .O(N__16571),
            .I(\b2v_inst.un2_indice_20_6 ));
    InMux I__3457 (
            .O(N__16568),
            .I(\b2v_inst.un2_indice_cry_5 ));
    CascadeMux I__3456 (
            .O(N__16565),
            .I(N__16562));
    InMux I__3455 (
            .O(N__16562),
            .I(N__16559));
    LocalMux I__3454 (
            .O(N__16559),
            .I(\b2v_inst.m7_1 ));
    CascadeMux I__3453 (
            .O(N__16556),
            .I(\b2v_inst.un8_dir_mem_3_c4_cascade_ ));
    InMux I__3452 (
            .O(N__16553),
            .I(N__16550));
    LocalMux I__3451 (
            .O(N__16550),
            .I(N__16547));
    Odrv4 I__3450 (
            .O(N__16547),
            .I(\b2v_inst.un8_dir_mem_3_c6 ));
    CascadeMux I__3449 (
            .O(N__16544),
            .I(\b2v_inst.un2_indice_1_1_4_cascade_ ));
    CascadeMux I__3448 (
            .O(N__16541),
            .I(N__16538));
    InMux I__3447 (
            .O(N__16538),
            .I(N__16535));
    LocalMux I__3446 (
            .O(N__16535),
            .I(N__16532));
    Span4Mux_h I__3445 (
            .O(N__16532),
            .I(N__16529));
    Odrv4 I__3444 (
            .O(N__16529),
            .I(\b2v_inst.dir_mem_2Z0Z_4 ));
    CascadeMux I__3443 (
            .O(N__16526),
            .I(N__16523));
    InMux I__3442 (
            .O(N__16523),
            .I(N__16520));
    LocalMux I__3441 (
            .O(N__16520),
            .I(N__16517));
    Span4Mux_h I__3440 (
            .O(N__16517),
            .I(N__16514));
    Sp12to4 I__3439 (
            .O(N__16514),
            .I(N__16511));
    Odrv12 I__3438 (
            .O(N__16511),
            .I(\b2v_inst.dir_mem_2Z0Z_1 ));
    InMux I__3437 (
            .O(N__16508),
            .I(N__16505));
    LocalMux I__3436 (
            .O(N__16505),
            .I(N__16502));
    Span4Mux_v I__3435 (
            .O(N__16502),
            .I(N__16499));
    Odrv4 I__3434 (
            .O(N__16499),
            .I(\b2v_inst.dir_mem_2Z0Z_2 ));
    CascadeMux I__3433 (
            .O(N__16496),
            .I(\b2v_inst.dir_mem_215_0_cascade_ ));
    InMux I__3432 (
            .O(N__16493),
            .I(N__16490));
    LocalMux I__3431 (
            .O(N__16490),
            .I(N__16487));
    Span4Mux_v I__3430 (
            .O(N__16487),
            .I(N__16484));
    Odrv4 I__3429 (
            .O(N__16484),
            .I(\b2v_inst.dir_mem_2Z0Z_0 ));
    InMux I__3428 (
            .O(N__16481),
            .I(N__16475));
    CascadeMux I__3427 (
            .O(N__16480),
            .I(N__16470));
    CascadeMux I__3426 (
            .O(N__16479),
            .I(N__16467));
    InMux I__3425 (
            .O(N__16478),
            .I(N__16462));
    LocalMux I__3424 (
            .O(N__16475),
            .I(N__16459));
    InMux I__3423 (
            .O(N__16474),
            .I(N__16455));
    InMux I__3422 (
            .O(N__16473),
            .I(N__16452));
    InMux I__3421 (
            .O(N__16470),
            .I(N__16445));
    InMux I__3420 (
            .O(N__16467),
            .I(N__16445));
    InMux I__3419 (
            .O(N__16466),
            .I(N__16445));
    InMux I__3418 (
            .O(N__16465),
            .I(N__16442));
    LocalMux I__3417 (
            .O(N__16462),
            .I(N__16437));
    Span4Mux_v I__3416 (
            .O(N__16459),
            .I(N__16437));
    InMux I__3415 (
            .O(N__16458),
            .I(N__16434));
    LocalMux I__3414 (
            .O(N__16455),
            .I(N__16431));
    LocalMux I__3413 (
            .O(N__16452),
            .I(\b2v_inst.N_237 ));
    LocalMux I__3412 (
            .O(N__16445),
            .I(\b2v_inst.N_237 ));
    LocalMux I__3411 (
            .O(N__16442),
            .I(\b2v_inst.N_237 ));
    Odrv4 I__3410 (
            .O(N__16437),
            .I(\b2v_inst.N_237 ));
    LocalMux I__3409 (
            .O(N__16434),
            .I(\b2v_inst.N_237 ));
    Odrv4 I__3408 (
            .O(N__16431),
            .I(\b2v_inst.N_237 ));
    CascadeMux I__3407 (
            .O(N__16418),
            .I(N__16415));
    InMux I__3406 (
            .O(N__16415),
            .I(N__16412));
    LocalMux I__3405 (
            .O(N__16412),
            .I(\b2v_inst.dir_mem_2Z0Z_7 ));
    InMux I__3404 (
            .O(N__16409),
            .I(N__16406));
    LocalMux I__3403 (
            .O(N__16406),
            .I(N__16402));
    CascadeMux I__3402 (
            .O(N__16405),
            .I(N__16397));
    Span4Mux_h I__3401 (
            .O(N__16402),
            .I(N__16391));
    InMux I__3400 (
            .O(N__16401),
            .I(N__16388));
    InMux I__3399 (
            .O(N__16400),
            .I(N__16381));
    InMux I__3398 (
            .O(N__16397),
            .I(N__16381));
    InMux I__3397 (
            .O(N__16396),
            .I(N__16381));
    InMux I__3396 (
            .O(N__16395),
            .I(N__16378));
    InMux I__3395 (
            .O(N__16394),
            .I(N__16375));
    Span4Mux_v I__3394 (
            .O(N__16391),
            .I(N__16371));
    LocalMux I__3393 (
            .O(N__16388),
            .I(N__16368));
    LocalMux I__3392 (
            .O(N__16381),
            .I(N__16361));
    LocalMux I__3391 (
            .O(N__16378),
            .I(N__16361));
    LocalMux I__3390 (
            .O(N__16375),
            .I(N__16361));
    InMux I__3389 (
            .O(N__16374),
            .I(N__16358));
    Odrv4 I__3388 (
            .O(N__16371),
            .I(\b2v_inst.N_239 ));
    Odrv4 I__3387 (
            .O(N__16368),
            .I(\b2v_inst.N_239 ));
    Odrv4 I__3386 (
            .O(N__16361),
            .I(\b2v_inst.N_239 ));
    LocalMux I__3385 (
            .O(N__16358),
            .I(\b2v_inst.N_239 ));
    CascadeMux I__3384 (
            .O(N__16349),
            .I(\b2v_inst.addr_ram_1_0_iv_i_1_7_cascade_ ));
    InMux I__3383 (
            .O(N__16346),
            .I(N__16343));
    LocalMux I__3382 (
            .O(N__16343),
            .I(N__16340));
    Span4Mux_h I__3381 (
            .O(N__16340),
            .I(N__16337));
    Odrv4 I__3380 (
            .O(N__16337),
            .I(\b2v_inst.addr_ram_1_0_iv_i_0_7 ));
    CascadeMux I__3379 (
            .O(N__16334),
            .I(N__16331));
    InMux I__3378 (
            .O(N__16331),
            .I(N__16327));
    CascadeMux I__3377 (
            .O(N__16330),
            .I(N__16324));
    LocalMux I__3376 (
            .O(N__16327),
            .I(N__16321));
    InMux I__3375 (
            .O(N__16324),
            .I(N__16318));
    Span4Mux_h I__3374 (
            .O(N__16321),
            .I(N__16315));
    LocalMux I__3373 (
            .O(N__16318),
            .I(N__16312));
    Span4Mux_h I__3372 (
            .O(N__16315),
            .I(N__16309));
    Odrv12 I__3371 (
            .O(N__16312),
            .I(N_50));
    Odrv4 I__3370 (
            .O(N__16309),
            .I(N_50));
    CascadeMux I__3369 (
            .O(N__16304),
            .I(\b2v_inst.g0_2_6_cascade_ ));
    InMux I__3368 (
            .O(N__16301),
            .I(N__16298));
    LocalMux I__3367 (
            .O(N__16298),
            .I(N__16295));
    Span4Mux_h I__3366 (
            .O(N__16295),
            .I(N__16292));
    Odrv4 I__3365 (
            .O(N__16292),
            .I(\b2v_inst.g0_2_8 ));
    CascadeMux I__3364 (
            .O(N__16289),
            .I(\b2v_inst.i4_mux_cascade_ ));
    InMux I__3363 (
            .O(N__16286),
            .I(N__16283));
    LocalMux I__3362 (
            .O(N__16283),
            .I(N__16280));
    Span4Mux_h I__3361 (
            .O(N__16280),
            .I(N__16277));
    Odrv4 I__3360 (
            .O(N__16277),
            .I(\b2v_inst.dir_mem_1Z0Z_6 ));
    InMux I__3359 (
            .O(N__16274),
            .I(N__16271));
    LocalMux I__3358 (
            .O(N__16271),
            .I(N__16267));
    InMux I__3357 (
            .O(N__16270),
            .I(N__16264));
    Odrv4 I__3356 (
            .O(N__16267),
            .I(\b2v_inst.un2_dir_mem_3_c5 ));
    LocalMux I__3355 (
            .O(N__16264),
            .I(\b2v_inst.un2_dir_mem_3_c5 ));
    CascadeMux I__3354 (
            .O(N__16259),
            .I(N__16256));
    InMux I__3353 (
            .O(N__16256),
            .I(N__16253));
    LocalMux I__3352 (
            .O(N__16253),
            .I(\b2v_inst.un2_dir_mem_3_ac0_3 ));
    CascadeMux I__3351 (
            .O(N__16250),
            .I(\b2v_inst.un2_dir_mem_3_ac0_3_cascade_ ));
    InMux I__3350 (
            .O(N__16247),
            .I(N__16244));
    LocalMux I__3349 (
            .O(N__16244),
            .I(N__16241));
    Odrv4 I__3348 (
            .O(N__16241),
            .I(\b2v_inst.un1_dir_mem_3_ns_1_5 ));
    CascadeMux I__3347 (
            .O(N__16238),
            .I(\b2v_inst.g4_0_cascade_ ));
    InMux I__3346 (
            .O(N__16235),
            .I(N__16232));
    LocalMux I__3345 (
            .O(N__16232),
            .I(\b2v_inst.g0_0 ));
    CascadeMux I__3344 (
            .O(N__16229),
            .I(N__16225));
    InMux I__3343 (
            .O(N__16228),
            .I(N__16218));
    InMux I__3342 (
            .O(N__16225),
            .I(N__16214));
    InMux I__3341 (
            .O(N__16224),
            .I(N__16211));
    InMux I__3340 (
            .O(N__16223),
            .I(N__16206));
    InMux I__3339 (
            .O(N__16222),
            .I(N__16206));
    InMux I__3338 (
            .O(N__16221),
            .I(N__16203));
    LocalMux I__3337 (
            .O(N__16218),
            .I(N__16199));
    InMux I__3336 (
            .O(N__16217),
            .I(N__16196));
    LocalMux I__3335 (
            .O(N__16214),
            .I(N__16187));
    LocalMux I__3334 (
            .O(N__16211),
            .I(N__16187));
    LocalMux I__3333 (
            .O(N__16206),
            .I(N__16187));
    LocalMux I__3332 (
            .O(N__16203),
            .I(N__16187));
    InMux I__3331 (
            .O(N__16202),
            .I(N__16184));
    Odrv4 I__3330 (
            .O(N__16199),
            .I(\b2v_inst.state_ns_a2_0_o2_1_0_2 ));
    LocalMux I__3329 (
            .O(N__16196),
            .I(\b2v_inst.state_ns_a2_0_o2_1_0_2 ));
    Odrv4 I__3328 (
            .O(N__16187),
            .I(\b2v_inst.state_ns_a2_0_o2_1_0_2 ));
    LocalMux I__3327 (
            .O(N__16184),
            .I(\b2v_inst.state_ns_a2_0_o2_1_0_2 ));
    InMux I__3326 (
            .O(N__16175),
            .I(N__16165));
    InMux I__3325 (
            .O(N__16174),
            .I(N__16162));
    InMux I__3324 (
            .O(N__16173),
            .I(N__16159));
    InMux I__3323 (
            .O(N__16172),
            .I(N__16152));
    InMux I__3322 (
            .O(N__16171),
            .I(N__16152));
    InMux I__3321 (
            .O(N__16170),
            .I(N__16152));
    InMux I__3320 (
            .O(N__16169),
            .I(N__16147));
    InMux I__3319 (
            .O(N__16168),
            .I(N__16144));
    LocalMux I__3318 (
            .O(N__16165),
            .I(N__16141));
    LocalMux I__3317 (
            .O(N__16162),
            .I(N__16138));
    LocalMux I__3316 (
            .O(N__16159),
            .I(N__16133));
    LocalMux I__3315 (
            .O(N__16152),
            .I(N__16133));
    InMux I__3314 (
            .O(N__16151),
            .I(N__16128));
    InMux I__3313 (
            .O(N__16150),
            .I(N__16128));
    LocalMux I__3312 (
            .O(N__16147),
            .I(\b2v_inst.cuenta_RNI4SC81Z0Z_7 ));
    LocalMux I__3311 (
            .O(N__16144),
            .I(\b2v_inst.cuenta_RNI4SC81Z0Z_7 ));
    Odrv4 I__3310 (
            .O(N__16141),
            .I(\b2v_inst.cuenta_RNI4SC81Z0Z_7 ));
    Odrv12 I__3309 (
            .O(N__16138),
            .I(\b2v_inst.cuenta_RNI4SC81Z0Z_7 ));
    Odrv4 I__3308 (
            .O(N__16133),
            .I(\b2v_inst.cuenta_RNI4SC81Z0Z_7 ));
    LocalMux I__3307 (
            .O(N__16128),
            .I(\b2v_inst.cuenta_RNI4SC81Z0Z_7 ));
    CascadeMux I__3306 (
            .O(N__16115),
            .I(N__16108));
    CascadeMux I__3305 (
            .O(N__16114),
            .I(N__16105));
    CascadeMux I__3304 (
            .O(N__16113),
            .I(N__16102));
    CascadeMux I__3303 (
            .O(N__16112),
            .I(N__16097));
    InMux I__3302 (
            .O(N__16111),
            .I(N__16094));
    InMux I__3301 (
            .O(N__16108),
            .I(N__16091));
    InMux I__3300 (
            .O(N__16105),
            .I(N__16088));
    InMux I__3299 (
            .O(N__16102),
            .I(N__16085));
    InMux I__3298 (
            .O(N__16101),
            .I(N__16078));
    InMux I__3297 (
            .O(N__16100),
            .I(N__16078));
    InMux I__3296 (
            .O(N__16097),
            .I(N__16078));
    LocalMux I__3295 (
            .O(N__16094),
            .I(N__16069));
    LocalMux I__3294 (
            .O(N__16091),
            .I(N__16069));
    LocalMux I__3293 (
            .O(N__16088),
            .I(N__16069));
    LocalMux I__3292 (
            .O(N__16085),
            .I(N__16064));
    LocalMux I__3291 (
            .O(N__16078),
            .I(N__16064));
    InMux I__3290 (
            .O(N__16077),
            .I(N__16059));
    InMux I__3289 (
            .O(N__16076),
            .I(N__16059));
    Span4Mux_v I__3288 (
            .O(N__16069),
            .I(N__16056));
    Span4Mux_h I__3287 (
            .O(N__16064),
            .I(N__16051));
    LocalMux I__3286 (
            .O(N__16059),
            .I(N__16051));
    Odrv4 I__3285 (
            .O(N__16056),
            .I(\b2v_inst.state_ns_a2_0_o2_0_2 ));
    Odrv4 I__3284 (
            .O(N__16051),
            .I(\b2v_inst.state_ns_a2_0_o2_0_2 ));
    CEMux I__3283 (
            .O(N__16046),
            .I(N__16041));
    CEMux I__3282 (
            .O(N__16045),
            .I(N__16038));
    CascadeMux I__3281 (
            .O(N__16044),
            .I(N__16034));
    LocalMux I__3280 (
            .O(N__16041),
            .I(N__16031));
    LocalMux I__3279 (
            .O(N__16038),
            .I(N__16028));
    InMux I__3278 (
            .O(N__16037),
            .I(N__16025));
    InMux I__3277 (
            .O(N__16034),
            .I(N__16020));
    Span4Mux_h I__3276 (
            .O(N__16031),
            .I(N__16017));
    Span4Mux_h I__3275 (
            .O(N__16028),
            .I(N__16014));
    LocalMux I__3274 (
            .O(N__16025),
            .I(N__16011));
    InMux I__3273 (
            .O(N__16024),
            .I(N__16008));
    InMux I__3272 (
            .O(N__16023),
            .I(N__16005));
    LocalMux I__3271 (
            .O(N__16020),
            .I(\b2v_inst.stateZ0Z_8 ));
    Odrv4 I__3270 (
            .O(N__16017),
            .I(\b2v_inst.stateZ0Z_8 ));
    Odrv4 I__3269 (
            .O(N__16014),
            .I(\b2v_inst.stateZ0Z_8 ));
    Odrv4 I__3268 (
            .O(N__16011),
            .I(\b2v_inst.stateZ0Z_8 ));
    LocalMux I__3267 (
            .O(N__16008),
            .I(\b2v_inst.stateZ0Z_8 ));
    LocalMux I__3266 (
            .O(N__16005),
            .I(\b2v_inst.stateZ0Z_8 ));
    CascadeMux I__3265 (
            .O(N__15992),
            .I(\b2v_inst.dir_mem_2_RNO_0Z0Z_3_cascade_ ));
    InMux I__3264 (
            .O(N__15989),
            .I(N__15986));
    LocalMux I__3263 (
            .O(N__15986),
            .I(N__15983));
    Odrv4 I__3262 (
            .O(N__15983),
            .I(\b2v_inst.dir_mem_2Z0Z_3 ));
    CascadeMux I__3261 (
            .O(N__15980),
            .I(N__15977));
    InMux I__3260 (
            .O(N__15977),
            .I(N__15974));
    LocalMux I__3259 (
            .O(N__15974),
            .I(N__15971));
    Span4Mux_h I__3258 (
            .O(N__15971),
            .I(N__15968));
    Odrv4 I__3257 (
            .O(N__15968),
            .I(\b2v_inst.un1_dir_mem_3_ns_1_4 ));
    InMux I__3256 (
            .O(N__15965),
            .I(N__15962));
    LocalMux I__3255 (
            .O(N__15962),
            .I(\b2v_inst.dir_mem_2_RNO_0Z0Z_7 ));
    InMux I__3254 (
            .O(N__15959),
            .I(N__15956));
    LocalMux I__3253 (
            .O(N__15956),
            .I(\b2v_inst.un2_indice_3_0_iv_0_a2_5_sx_2 ));
    CascadeMux I__3252 (
            .O(N__15953),
            .I(\b2v_inst.N_452_cascade_ ));
    InMux I__3251 (
            .O(N__15950),
            .I(N__15947));
    LocalMux I__3250 (
            .O(N__15947),
            .I(N__15942));
    InMux I__3249 (
            .O(N__15946),
            .I(N__15937));
    InMux I__3248 (
            .O(N__15945),
            .I(N__15937));
    Span4Mux_h I__3247 (
            .O(N__15942),
            .I(N__15934));
    LocalMux I__3246 (
            .O(N__15937),
            .I(N__15931));
    Odrv4 I__3245 (
            .O(N__15934),
            .I(\b2v_inst.stateZ0Z_13 ));
    Odrv4 I__3244 (
            .O(N__15931),
            .I(\b2v_inst.stateZ0Z_13 ));
    InMux I__3243 (
            .O(N__15926),
            .I(N__15923));
    LocalMux I__3242 (
            .O(N__15923),
            .I(N__15920));
    Span4Mux_h I__3241 (
            .O(N__15920),
            .I(N__15917));
    Odrv4 I__3240 (
            .O(N__15917),
            .I(\b2v_inst.g2_3 ));
    InMux I__3239 (
            .O(N__15914),
            .I(N__15911));
    LocalMux I__3238 (
            .O(N__15911),
            .I(N__15907));
    InMux I__3237 (
            .O(N__15910),
            .I(N__15904));
    Span4Mux_h I__3236 (
            .O(N__15907),
            .I(N__15896));
    LocalMux I__3235 (
            .O(N__15904),
            .I(N__15896));
    InMux I__3234 (
            .O(N__15903),
            .I(N__15893));
    InMux I__3233 (
            .O(N__15902),
            .I(N__15890));
    InMux I__3232 (
            .O(N__15901),
            .I(N__15887));
    Span4Mux_h I__3231 (
            .O(N__15896),
            .I(N__15884));
    LocalMux I__3230 (
            .O(N__15893),
            .I(N__15879));
    LocalMux I__3229 (
            .O(N__15890),
            .I(N__15879));
    LocalMux I__3228 (
            .O(N__15887),
            .I(\b2v_inst.borradoZ0 ));
    Odrv4 I__3227 (
            .O(N__15884),
            .I(\b2v_inst.borradoZ0 ));
    Odrv12 I__3226 (
            .O(N__15879),
            .I(\b2v_inst.borradoZ0 ));
    InMux I__3225 (
            .O(N__15872),
            .I(N__15868));
    InMux I__3224 (
            .O(N__15871),
            .I(N__15862));
    LocalMux I__3223 (
            .O(N__15868),
            .I(N__15859));
    InMux I__3222 (
            .O(N__15867),
            .I(N__15854));
    InMux I__3221 (
            .O(N__15866),
            .I(N__15854));
    InMux I__3220 (
            .O(N__15865),
            .I(N__15851));
    LocalMux I__3219 (
            .O(N__15862),
            .I(N__15848));
    Span4Mux_h I__3218 (
            .O(N__15859),
            .I(N__15841));
    LocalMux I__3217 (
            .O(N__15854),
            .I(N__15838));
    LocalMux I__3216 (
            .O(N__15851),
            .I(N__15835));
    Span4Mux_h I__3215 (
            .O(N__15848),
            .I(N__15832));
    InMux I__3214 (
            .O(N__15847),
            .I(N__15829));
    InMux I__3213 (
            .O(N__15846),
            .I(N__15822));
    InMux I__3212 (
            .O(N__15845),
            .I(N__15822));
    InMux I__3211 (
            .O(N__15844),
            .I(N__15822));
    Odrv4 I__3210 (
            .O(N__15841),
            .I(\b2v_inst.stateZ0Z_5 ));
    Odrv12 I__3209 (
            .O(N__15838),
            .I(\b2v_inst.stateZ0Z_5 ));
    Odrv4 I__3208 (
            .O(N__15835),
            .I(\b2v_inst.stateZ0Z_5 ));
    Odrv4 I__3207 (
            .O(N__15832),
            .I(\b2v_inst.stateZ0Z_5 ));
    LocalMux I__3206 (
            .O(N__15829),
            .I(\b2v_inst.stateZ0Z_5 ));
    LocalMux I__3205 (
            .O(N__15822),
            .I(\b2v_inst.stateZ0Z_5 ));
    CascadeMux I__3204 (
            .O(N__15809),
            .I(\b2v_inst.N_7_1_cascade_ ));
    CascadeMux I__3203 (
            .O(N__15806),
            .I(\b2v_inst.g2_2_cascade_ ));
    InMux I__3202 (
            .O(N__15803),
            .I(N__15800));
    LocalMux I__3201 (
            .O(N__15800),
            .I(\b2v_inst.g1 ));
    InMux I__3200 (
            .O(N__15797),
            .I(N__15794));
    LocalMux I__3199 (
            .O(N__15794),
            .I(\b2v_inst.un2_indice_21_s0_0_6 ));
    CascadeMux I__3198 (
            .O(N__15791),
            .I(\b2v_inst.N_253_cascade_ ));
    InMux I__3197 (
            .O(N__15788),
            .I(N__15782));
    InMux I__3196 (
            .O(N__15787),
            .I(N__15782));
    LocalMux I__3195 (
            .O(N__15782),
            .I(N__15779));
    Odrv4 I__3194 (
            .O(N__15779),
            .I(\b2v_inst.state_fastZ0Z_17 ));
    InMux I__3193 (
            .O(N__15776),
            .I(N__15770));
    InMux I__3192 (
            .O(N__15775),
            .I(N__15770));
    LocalMux I__3191 (
            .O(N__15770),
            .I(N__15767));
    Odrv4 I__3190 (
            .O(N__15767),
            .I(\b2v_inst.state_fastZ0Z_15 ));
    CascadeMux I__3189 (
            .O(N__15764),
            .I(\b2v_inst.N_253_i_cascade_ ));
    InMux I__3188 (
            .O(N__15761),
            .I(N__15758));
    LocalMux I__3187 (
            .O(N__15758),
            .I(N__15755));
    Odrv4 I__3186 (
            .O(N__15755),
            .I(\b2v_inst.dir_mem_3_RNO_0Z0Z_3 ));
    CascadeMux I__3185 (
            .O(N__15752),
            .I(\b2v_inst1.r_RX_Bytece_0_0_1_cascade_ ));
    InMux I__3184 (
            .O(N__15749),
            .I(N__15746));
    LocalMux I__3183 (
            .O(N__15746),
            .I(N__15743));
    Span4Mux_h I__3182 (
            .O(N__15743),
            .I(N__15739));
    InMux I__3181 (
            .O(N__15742),
            .I(N__15736));
    Odrv4 I__3180 (
            .O(N__15739),
            .I(SYNTHESIZED_WIRE_10_1));
    LocalMux I__3179 (
            .O(N__15736),
            .I(SYNTHESIZED_WIRE_10_1));
    InMux I__3178 (
            .O(N__15731),
            .I(N__15728));
    LocalMux I__3177 (
            .O(N__15728),
            .I(\b2v_inst.dir_mem_2_RNO_0Z0Z_6 ));
    InMux I__3176 (
            .O(N__15725),
            .I(N__15722));
    LocalMux I__3175 (
            .O(N__15722),
            .I(N__15716));
    InMux I__3174 (
            .O(N__15721),
            .I(N__15711));
    InMux I__3173 (
            .O(N__15720),
            .I(N__15711));
    CascadeMux I__3172 (
            .O(N__15719),
            .I(N__15708));
    Span4Mux_h I__3171 (
            .O(N__15716),
            .I(N__15705));
    LocalMux I__3170 (
            .O(N__15711),
            .I(N__15702));
    InMux I__3169 (
            .O(N__15708),
            .I(N__15699));
    Span4Mux_v I__3168 (
            .O(N__15705),
            .I(N__15696));
    Span12Mux_v I__3167 (
            .O(N__15702),
            .I(N__15693));
    LocalMux I__3166 (
            .O(N__15699),
            .I(SYNTHESIZED_WIRE_9));
    Odrv4 I__3165 (
            .O(N__15696),
            .I(SYNTHESIZED_WIRE_9));
    Odrv12 I__3164 (
            .O(N__15693),
            .I(SYNTHESIZED_WIRE_9));
    CascadeMux I__3163 (
            .O(N__15686),
            .I(N__15674));
    CascadeMux I__3162 (
            .O(N__15685),
            .I(N__15671));
    InMux I__3161 (
            .O(N__15684),
            .I(N__15668));
    InMux I__3160 (
            .O(N__15683),
            .I(N__15665));
    InMux I__3159 (
            .O(N__15682),
            .I(N__15660));
    InMux I__3158 (
            .O(N__15681),
            .I(N__15660));
    InMux I__3157 (
            .O(N__15680),
            .I(N__15655));
    InMux I__3156 (
            .O(N__15679),
            .I(N__15655));
    InMux I__3155 (
            .O(N__15678),
            .I(N__15652));
    InMux I__3154 (
            .O(N__15677),
            .I(N__15645));
    InMux I__3153 (
            .O(N__15674),
            .I(N__15645));
    InMux I__3152 (
            .O(N__15671),
            .I(N__15645));
    LocalMux I__3151 (
            .O(N__15668),
            .I(N__15642));
    LocalMux I__3150 (
            .O(N__15665),
            .I(N__15639));
    LocalMux I__3149 (
            .O(N__15660),
            .I(N__15634));
    LocalMux I__3148 (
            .O(N__15655),
            .I(N__15634));
    LocalMux I__3147 (
            .O(N__15652),
            .I(N__15629));
    LocalMux I__3146 (
            .O(N__15645),
            .I(N__15626));
    Span12Mux_h I__3145 (
            .O(N__15642),
            .I(N__15621));
    Span12Mux_s8_h I__3144 (
            .O(N__15639),
            .I(N__15621));
    Span4Mux_h I__3143 (
            .O(N__15634),
            .I(N__15618));
    InMux I__3142 (
            .O(N__15633),
            .I(N__15613));
    InMux I__3141 (
            .O(N__15632),
            .I(N__15613));
    Span4Mux_v I__3140 (
            .O(N__15629),
            .I(N__15608));
    Span4Mux_v I__3139 (
            .O(N__15626),
            .I(N__15608));
    Odrv12 I__3138 (
            .O(N__15621),
            .I(\b2v_inst.stateZ0Z_16 ));
    Odrv4 I__3137 (
            .O(N__15618),
            .I(\b2v_inst.stateZ0Z_16 ));
    LocalMux I__3136 (
            .O(N__15613),
            .I(\b2v_inst.stateZ0Z_16 ));
    Odrv4 I__3135 (
            .O(N__15608),
            .I(\b2v_inst.stateZ0Z_16 ));
    InMux I__3134 (
            .O(N__15599),
            .I(N__15581));
    InMux I__3133 (
            .O(N__15598),
            .I(N__15581));
    InMux I__3132 (
            .O(N__15597),
            .I(N__15581));
    InMux I__3131 (
            .O(N__15596),
            .I(N__15581));
    InMux I__3130 (
            .O(N__15595),
            .I(N__15581));
    InMux I__3129 (
            .O(N__15594),
            .I(N__15581));
    LocalMux I__3128 (
            .O(N__15581),
            .I(N__15578));
    Span4Mux_v I__3127 (
            .O(N__15578),
            .I(N__15572));
    InMux I__3126 (
            .O(N__15577),
            .I(N__15567));
    InMux I__3125 (
            .O(N__15576),
            .I(N__15567));
    CascadeMux I__3124 (
            .O(N__15575),
            .I(N__15560));
    Span4Mux_v I__3123 (
            .O(N__15572),
            .I(N__15554));
    LocalMux I__3122 (
            .O(N__15567),
            .I(N__15554));
    InMux I__3121 (
            .O(N__15566),
            .I(N__15541));
    InMux I__3120 (
            .O(N__15565),
            .I(N__15541));
    InMux I__3119 (
            .O(N__15564),
            .I(N__15541));
    InMux I__3118 (
            .O(N__15563),
            .I(N__15541));
    InMux I__3117 (
            .O(N__15560),
            .I(N__15541));
    InMux I__3116 (
            .O(N__15559),
            .I(N__15541));
    Span4Mux_h I__3115 (
            .O(N__15554),
            .I(N__15536));
    LocalMux I__3114 (
            .O(N__15541),
            .I(N__15536));
    Span4Mux_v I__3113 (
            .O(N__15536),
            .I(N__15531));
    InMux I__3112 (
            .O(N__15535),
            .I(N__15526));
    InMux I__3111 (
            .O(N__15534),
            .I(N__15526));
    Odrv4 I__3110 (
            .O(N__15531),
            .I(\b2v_inst.ignorar_anteriorZ0 ));
    LocalMux I__3109 (
            .O(N__15526),
            .I(\b2v_inst.ignorar_anteriorZ0 ));
    CEMux I__3108 (
            .O(N__15521),
            .I(N__15518));
    LocalMux I__3107 (
            .O(N__15518),
            .I(N__15515));
    Span4Mux_h I__3106 (
            .O(N__15515),
            .I(N__15512));
    Span4Mux_h I__3105 (
            .O(N__15512),
            .I(N__15509));
    Odrv4 I__3104 (
            .O(N__15509),
            .I(\b2v_inst.un1_state_19_0 ));
    CascadeMux I__3103 (
            .O(N__15506),
            .I(N__15503));
    InMux I__3102 (
            .O(N__15503),
            .I(N__15500));
    LocalMux I__3101 (
            .O(N__15500),
            .I(N__15497));
    Span4Mux_v I__3100 (
            .O(N__15497),
            .I(N__15494));
    Odrv4 I__3099 (
            .O(N__15494),
            .I(\b2v_inst.N_5 ));
    CEMux I__3098 (
            .O(N__15491),
            .I(N__15487));
    CEMux I__3097 (
            .O(N__15490),
            .I(N__15484));
    LocalMux I__3096 (
            .O(N__15487),
            .I(N__15481));
    LocalMux I__3095 (
            .O(N__15484),
            .I(N__15478));
    Span4Mux_h I__3094 (
            .O(N__15481),
            .I(N__15474));
    Span4Mux_h I__3093 (
            .O(N__15478),
            .I(N__15471));
    InMux I__3092 (
            .O(N__15477),
            .I(N__15466));
    Span4Mux_v I__3091 (
            .O(N__15474),
            .I(N__15463));
    Span4Mux_h I__3090 (
            .O(N__15471),
            .I(N__15460));
    InMux I__3089 (
            .O(N__15470),
            .I(N__15457));
    InMux I__3088 (
            .O(N__15469),
            .I(N__15454));
    LocalMux I__3087 (
            .O(N__15466),
            .I(N__15451));
    Odrv4 I__3086 (
            .O(N__15463),
            .I(\b2v_inst.stateZ0Z_10 ));
    Odrv4 I__3085 (
            .O(N__15460),
            .I(\b2v_inst.stateZ0Z_10 ));
    LocalMux I__3084 (
            .O(N__15457),
            .I(\b2v_inst.stateZ0Z_10 ));
    LocalMux I__3083 (
            .O(N__15454),
            .I(\b2v_inst.stateZ0Z_10 ));
    Odrv4 I__3082 (
            .O(N__15451),
            .I(\b2v_inst.stateZ0Z_10 ));
    InMux I__3081 (
            .O(N__15440),
            .I(N__15434));
    InMux I__3080 (
            .O(N__15439),
            .I(N__15434));
    LocalMux I__3079 (
            .O(N__15434),
            .I(\b2v_inst.stateZ0Z_1 ));
    CascadeMux I__3078 (
            .O(N__15431),
            .I(N__15428));
    InMux I__3077 (
            .O(N__15428),
            .I(N__15425));
    LocalMux I__3076 (
            .O(N__15425),
            .I(N__15422));
    Odrv4 I__3075 (
            .O(N__15422),
            .I(\b2v_inst.dir_mem_3Z0Z_4 ));
    CascadeMux I__3074 (
            .O(N__15419),
            .I(\b2v_inst.addr_ram_1_0_iv_i_1_4_cascade_ ));
    CascadeMux I__3073 (
            .O(N__15416),
            .I(N__15413));
    InMux I__3072 (
            .O(N__15413),
            .I(N__15409));
    CascadeMux I__3071 (
            .O(N__15412),
            .I(N__15406));
    LocalMux I__3070 (
            .O(N__15409),
            .I(N__15403));
    InMux I__3069 (
            .O(N__15406),
            .I(N__15400));
    Span4Mux_v I__3068 (
            .O(N__15403),
            .I(N__15395));
    LocalMux I__3067 (
            .O(N__15400),
            .I(N__15395));
    Span4Mux_h I__3066 (
            .O(N__15395),
            .I(N__15392));
    Odrv4 I__3065 (
            .O(N__15392),
            .I(N_163));
    CascadeMux I__3064 (
            .O(N__15389),
            .I(\b2v_inst.g0_11_1_cascade_ ));
    InMux I__3063 (
            .O(N__15386),
            .I(N__15383));
    LocalMux I__3062 (
            .O(N__15383),
            .I(\b2v_inst.dir_mem_1Z0Z_4 ));
    InMux I__3061 (
            .O(N__15380),
            .I(N__15377));
    LocalMux I__3060 (
            .O(N__15377),
            .I(N__15366));
    InMux I__3059 (
            .O(N__15376),
            .I(N__15363));
    InMux I__3058 (
            .O(N__15375),
            .I(N__15360));
    InMux I__3057 (
            .O(N__15374),
            .I(N__15357));
    InMux I__3056 (
            .O(N__15373),
            .I(N__15350));
    InMux I__3055 (
            .O(N__15372),
            .I(N__15350));
    InMux I__3054 (
            .O(N__15371),
            .I(N__15350));
    InMux I__3053 (
            .O(N__15370),
            .I(N__15345));
    InMux I__3052 (
            .O(N__15369),
            .I(N__15345));
    Odrv4 I__3051 (
            .O(N__15366),
            .I(\b2v_inst.N_235 ));
    LocalMux I__3050 (
            .O(N__15363),
            .I(\b2v_inst.N_235 ));
    LocalMux I__3049 (
            .O(N__15360),
            .I(\b2v_inst.N_235 ));
    LocalMux I__3048 (
            .O(N__15357),
            .I(\b2v_inst.N_235 ));
    LocalMux I__3047 (
            .O(N__15350),
            .I(\b2v_inst.N_235 ));
    LocalMux I__3046 (
            .O(N__15345),
            .I(\b2v_inst.N_235 ));
    InMux I__3045 (
            .O(N__15332),
            .I(N__15329));
    LocalMux I__3044 (
            .O(N__15329),
            .I(\b2v_inst.addr_ram_1_0_iv_i_0_4 ));
    CascadeMux I__3043 (
            .O(N__15326),
            .I(N__15321));
    CascadeMux I__3042 (
            .O(N__15325),
            .I(N__15318));
    InMux I__3041 (
            .O(N__15324),
            .I(N__15312));
    InMux I__3040 (
            .O(N__15321),
            .I(N__15301));
    InMux I__3039 (
            .O(N__15318),
            .I(N__15301));
    InMux I__3038 (
            .O(N__15317),
            .I(N__15301));
    InMux I__3037 (
            .O(N__15316),
            .I(N__15301));
    InMux I__3036 (
            .O(N__15315),
            .I(N__15301));
    LocalMux I__3035 (
            .O(N__15312),
            .I(\b2v_inst.dir_mem_315_0 ));
    LocalMux I__3034 (
            .O(N__15301),
            .I(\b2v_inst.dir_mem_315_0 ));
    InMux I__3033 (
            .O(N__15296),
            .I(N__15293));
    LocalMux I__3032 (
            .O(N__15293),
            .I(N__15290));
    Odrv4 I__3031 (
            .O(N__15290),
            .I(\b2v_inst.dir_mem_3Z0Z_3 ));
    InMux I__3030 (
            .O(N__15287),
            .I(N__15284));
    LocalMux I__3029 (
            .O(N__15284),
            .I(N__15281));
    Span4Mux_h I__3028 (
            .O(N__15281),
            .I(N__15278));
    Odrv4 I__3027 (
            .O(N__15278),
            .I(\b2v_inst.dir_mem_3Z0Z_7 ));
    CEMux I__3026 (
            .O(N__15275),
            .I(N__15271));
    CEMux I__3025 (
            .O(N__15274),
            .I(N__15268));
    LocalMux I__3024 (
            .O(N__15271),
            .I(N__15263));
    LocalMux I__3023 (
            .O(N__15268),
            .I(N__15263));
    Span4Mux_v I__3022 (
            .O(N__15263),
            .I(N__15260));
    Span4Mux_v I__3021 (
            .O(N__15260),
            .I(N__15257));
    Sp12to4 I__3020 (
            .O(N__15257),
            .I(N__15254));
    Odrv12 I__3019 (
            .O(N__15254),
            .I(\b2v_inst.N_138_i ));
    InMux I__3018 (
            .O(N__15251),
            .I(N__15248));
    LocalMux I__3017 (
            .O(N__15248),
            .I(N__15245));
    Span4Mux_v I__3016 (
            .O(N__15245),
            .I(N__15242));
    Odrv4 I__3015 (
            .O(N__15242),
            .I(\b2v_inst1.r_RX_Bytece_0_5 ));
    CEMux I__3014 (
            .O(N__15239),
            .I(N__15236));
    LocalMux I__3013 (
            .O(N__15236),
            .I(N__15231));
    CEMux I__3012 (
            .O(N__15235),
            .I(N__15228));
    InMux I__3011 (
            .O(N__15234),
            .I(N__15225));
    Span4Mux_h I__3010 (
            .O(N__15231),
            .I(N__15219));
    LocalMux I__3009 (
            .O(N__15228),
            .I(N__15219));
    LocalMux I__3008 (
            .O(N__15225),
            .I(N__15216));
    CascadeMux I__3007 (
            .O(N__15224),
            .I(N__15210));
    Span4Mux_v I__3006 (
            .O(N__15219),
            .I(N__15207));
    Span4Mux_h I__3005 (
            .O(N__15216),
            .I(N__15204));
    InMux I__3004 (
            .O(N__15215),
            .I(N__15197));
    InMux I__3003 (
            .O(N__15214),
            .I(N__15197));
    InMux I__3002 (
            .O(N__15213),
            .I(N__15197));
    InMux I__3001 (
            .O(N__15210),
            .I(N__15194));
    Odrv4 I__3000 (
            .O(N__15207),
            .I(\b2v_inst.stateZ0Z_14 ));
    Odrv4 I__2999 (
            .O(N__15204),
            .I(\b2v_inst.stateZ0Z_14 ));
    LocalMux I__2998 (
            .O(N__15197),
            .I(\b2v_inst.stateZ0Z_14 ));
    LocalMux I__2997 (
            .O(N__15194),
            .I(\b2v_inst.stateZ0Z_14 ));
    InMux I__2996 (
            .O(N__15185),
            .I(N__15177));
    InMux I__2995 (
            .O(N__15184),
            .I(N__15174));
    InMux I__2994 (
            .O(N__15183),
            .I(N__15165));
    InMux I__2993 (
            .O(N__15182),
            .I(N__15165));
    InMux I__2992 (
            .O(N__15181),
            .I(N__15165));
    InMux I__2991 (
            .O(N__15180),
            .I(N__15165));
    LocalMux I__2990 (
            .O(N__15177),
            .I(N__15162));
    LocalMux I__2989 (
            .O(N__15174),
            .I(N__15157));
    LocalMux I__2988 (
            .O(N__15165),
            .I(N__15157));
    Span12Mux_h I__2987 (
            .O(N__15162),
            .I(N__15154));
    Span4Mux_v I__2986 (
            .O(N__15157),
            .I(N__15151));
    Odrv12 I__2985 (
            .O(N__15154),
            .I(\b2v_inst.stateZ0Z_6 ));
    Odrv4 I__2984 (
            .O(N__15151),
            .I(\b2v_inst.stateZ0Z_6 ));
    InMux I__2983 (
            .O(N__15146),
            .I(N__15140));
    InMux I__2982 (
            .O(N__15145),
            .I(N__15140));
    LocalMux I__2981 (
            .O(N__15140),
            .I(N__15135));
    InMux I__2980 (
            .O(N__15139),
            .I(N__15132));
    InMux I__2979 (
            .O(N__15138),
            .I(N__15129));
    Span4Mux_v I__2978 (
            .O(N__15135),
            .I(N__15126));
    LocalMux I__2977 (
            .O(N__15132),
            .I(\b2v_inst.state_RNITETBZ0Z_0 ));
    LocalMux I__2976 (
            .O(N__15129),
            .I(\b2v_inst.state_RNITETBZ0Z_0 ));
    Odrv4 I__2975 (
            .O(N__15126),
            .I(\b2v_inst.state_RNITETBZ0Z_0 ));
    CascadeMux I__2974 (
            .O(N__15119),
            .I(\b2v_inst.N_351_cascade_ ));
    InMux I__2973 (
            .O(N__15116),
            .I(N__15113));
    LocalMux I__2972 (
            .O(N__15113),
            .I(\b2v_inst.addr_ram_1_iv_i_1_3 ));
    CascadeMux I__2971 (
            .O(N__15110),
            .I(\b2v_inst.addr_ram_1_iv_i_2_3_cascade_ ));
    CascadeMux I__2970 (
            .O(N__15107),
            .I(N__15104));
    InMux I__2969 (
            .O(N__15104),
            .I(N__15100));
    CascadeMux I__2968 (
            .O(N__15103),
            .I(N__15097));
    LocalMux I__2967 (
            .O(N__15100),
            .I(N__15094));
    InMux I__2966 (
            .O(N__15097),
            .I(N__15091));
    Span4Mux_v I__2965 (
            .O(N__15094),
            .I(N__15086));
    LocalMux I__2964 (
            .O(N__15091),
            .I(N__15086));
    Span4Mux_h I__2963 (
            .O(N__15086),
            .I(N__15083));
    Odrv4 I__2962 (
            .O(N__15083),
            .I(N_58));
    InMux I__2961 (
            .O(N__15080),
            .I(N__15077));
    LocalMux I__2960 (
            .O(N__15077),
            .I(N__15074));
    Span4Mux_v I__2959 (
            .O(N__15074),
            .I(N__15070));
    InMux I__2958 (
            .O(N__15073),
            .I(N__15067));
    Odrv4 I__2957 (
            .O(N__15070),
            .I(\b2v_inst.stateZ0Z_0 ));
    LocalMux I__2956 (
            .O(N__15067),
            .I(\b2v_inst.stateZ0Z_0 ));
    CascadeMux I__2955 (
            .O(N__15062),
            .I(N__15055));
    InMux I__2954 (
            .O(N__15061),
            .I(N__15046));
    InMux I__2953 (
            .O(N__15060),
            .I(N__15046));
    InMux I__2952 (
            .O(N__15059),
            .I(N__15046));
    InMux I__2951 (
            .O(N__15058),
            .I(N__15043));
    InMux I__2950 (
            .O(N__15055),
            .I(N__15036));
    InMux I__2949 (
            .O(N__15054),
            .I(N__15036));
    InMux I__2948 (
            .O(N__15053),
            .I(N__15036));
    LocalMux I__2947 (
            .O(N__15046),
            .I(\b2v_inst.cuentaZ0Z_5 ));
    LocalMux I__2946 (
            .O(N__15043),
            .I(\b2v_inst.cuentaZ0Z_5 ));
    LocalMux I__2945 (
            .O(N__15036),
            .I(\b2v_inst.cuentaZ0Z_5 ));
    CascadeMux I__2944 (
            .O(N__15029),
            .I(N__15023));
    InMux I__2943 (
            .O(N__15028),
            .I(N__15017));
    InMux I__2942 (
            .O(N__15027),
            .I(N__15008));
    InMux I__2941 (
            .O(N__15026),
            .I(N__15008));
    InMux I__2940 (
            .O(N__15023),
            .I(N__15008));
    InMux I__2939 (
            .O(N__15022),
            .I(N__15008));
    InMux I__2938 (
            .O(N__15021),
            .I(N__15003));
    InMux I__2937 (
            .O(N__15020),
            .I(N__15003));
    LocalMux I__2936 (
            .O(N__15017),
            .I(N__14998));
    LocalMux I__2935 (
            .O(N__15008),
            .I(N__14998));
    LocalMux I__2934 (
            .O(N__15003),
            .I(\b2v_inst.cuentaZ0Z_4 ));
    Odrv4 I__2933 (
            .O(N__14998),
            .I(\b2v_inst.cuentaZ0Z_4 ));
    CascadeMux I__2932 (
            .O(N__14993),
            .I(\b2v_inst.un4_cuenta_ac0_9_0_cascade_ ));
    InMux I__2931 (
            .O(N__14990),
            .I(N__14981));
    InMux I__2930 (
            .O(N__14989),
            .I(N__14978));
    InMux I__2929 (
            .O(N__14988),
            .I(N__14975));
    InMux I__2928 (
            .O(N__14987),
            .I(N__14966));
    InMux I__2927 (
            .O(N__14986),
            .I(N__14966));
    InMux I__2926 (
            .O(N__14985),
            .I(N__14966));
    InMux I__2925 (
            .O(N__14984),
            .I(N__14966));
    LocalMux I__2924 (
            .O(N__14981),
            .I(\b2v_inst.un4_cuenta_c4 ));
    LocalMux I__2923 (
            .O(N__14978),
            .I(\b2v_inst.un4_cuenta_c4 ));
    LocalMux I__2922 (
            .O(N__14975),
            .I(\b2v_inst.un4_cuenta_c4 ));
    LocalMux I__2921 (
            .O(N__14966),
            .I(\b2v_inst.un4_cuenta_c4 ));
    InMux I__2920 (
            .O(N__14957),
            .I(N__14949));
    InMux I__2919 (
            .O(N__14956),
            .I(N__14942));
    InMux I__2918 (
            .O(N__14955),
            .I(N__14942));
    InMux I__2917 (
            .O(N__14954),
            .I(N__14942));
    InMux I__2916 (
            .O(N__14953),
            .I(N__14939));
    InMux I__2915 (
            .O(N__14952),
            .I(N__14936));
    LocalMux I__2914 (
            .O(N__14949),
            .I(\b2v_inst.cuentaZ0Z_6 ));
    LocalMux I__2913 (
            .O(N__14942),
            .I(\b2v_inst.cuentaZ0Z_6 ));
    LocalMux I__2912 (
            .O(N__14939),
            .I(\b2v_inst.cuentaZ0Z_6 ));
    LocalMux I__2911 (
            .O(N__14936),
            .I(\b2v_inst.cuentaZ0Z_6 ));
    InMux I__2910 (
            .O(N__14927),
            .I(N__14919));
    InMux I__2909 (
            .O(N__14926),
            .I(N__14919));
    InMux I__2908 (
            .O(N__14925),
            .I(N__14916));
    InMux I__2907 (
            .O(N__14924),
            .I(N__14913));
    LocalMux I__2906 (
            .O(N__14919),
            .I(\b2v_inst.cuentaZ0Z_7 ));
    LocalMux I__2905 (
            .O(N__14916),
            .I(\b2v_inst.cuentaZ0Z_7 ));
    LocalMux I__2904 (
            .O(N__14913),
            .I(\b2v_inst.cuentaZ0Z_7 ));
    CEMux I__2903 (
            .O(N__14906),
            .I(N__14902));
    CEMux I__2902 (
            .O(N__14905),
            .I(N__14899));
    LocalMux I__2901 (
            .O(N__14902),
            .I(N__14892));
    LocalMux I__2900 (
            .O(N__14899),
            .I(N__14892));
    CEMux I__2899 (
            .O(N__14898),
            .I(N__14889));
    CEMux I__2898 (
            .O(N__14897),
            .I(N__14886));
    Span4Mux_v I__2897 (
            .O(N__14892),
            .I(N__14883));
    LocalMux I__2896 (
            .O(N__14889),
            .I(N__14880));
    LocalMux I__2895 (
            .O(N__14886),
            .I(\b2v_inst.N_399_i ));
    Odrv4 I__2894 (
            .O(N__14883),
            .I(\b2v_inst.N_399_i ));
    Odrv4 I__2893 (
            .O(N__14880),
            .I(\b2v_inst.N_399_i ));
    InMux I__2892 (
            .O(N__14873),
            .I(N__14869));
    InMux I__2891 (
            .O(N__14872),
            .I(N__14866));
    LocalMux I__2890 (
            .O(N__14869),
            .I(N__14863));
    LocalMux I__2889 (
            .O(N__14866),
            .I(N__14860));
    Span4Mux_h I__2888 (
            .O(N__14863),
            .I(N__14853));
    Span4Mux_v I__2887 (
            .O(N__14860),
            .I(N__14850));
    InMux I__2886 (
            .O(N__14859),
            .I(N__14847));
    InMux I__2885 (
            .O(N__14858),
            .I(N__14844));
    InMux I__2884 (
            .O(N__14857),
            .I(N__14839));
    InMux I__2883 (
            .O(N__14856),
            .I(N__14839));
    Span4Mux_h I__2882 (
            .O(N__14853),
            .I(N__14834));
    Span4Mux_h I__2881 (
            .O(N__14850),
            .I(N__14834));
    LocalMux I__2880 (
            .O(N__14847),
            .I(\b2v_inst.N_227 ));
    LocalMux I__2879 (
            .O(N__14844),
            .I(\b2v_inst.N_227 ));
    LocalMux I__2878 (
            .O(N__14839),
            .I(\b2v_inst.N_227 ));
    Odrv4 I__2877 (
            .O(N__14834),
            .I(\b2v_inst.N_227 ));
    InMux I__2876 (
            .O(N__14825),
            .I(N__14821));
    InMux I__2875 (
            .O(N__14824),
            .I(N__14817));
    LocalMux I__2874 (
            .O(N__14821),
            .I(N__14814));
    InMux I__2873 (
            .O(N__14820),
            .I(N__14811));
    LocalMux I__2872 (
            .O(N__14817),
            .I(N__14808));
    Odrv4 I__2871 (
            .O(N__14814),
            .I(\b2v_inst.N_232 ));
    LocalMux I__2870 (
            .O(N__14811),
            .I(\b2v_inst.N_232 ));
    Odrv12 I__2869 (
            .O(N__14808),
            .I(\b2v_inst.N_232 ));
    CascadeMux I__2868 (
            .O(N__14801),
            .I(\b2v_inst.N_232_cascade_ ));
    InMux I__2867 (
            .O(N__14798),
            .I(N__14788));
    InMux I__2866 (
            .O(N__14797),
            .I(N__14782));
    CascadeMux I__2865 (
            .O(N__14796),
            .I(N__14778));
    InMux I__2864 (
            .O(N__14795),
            .I(N__14769));
    InMux I__2863 (
            .O(N__14794),
            .I(N__14769));
    InMux I__2862 (
            .O(N__14793),
            .I(N__14769));
    InMux I__2861 (
            .O(N__14792),
            .I(N__14769));
    InMux I__2860 (
            .O(N__14791),
            .I(N__14766));
    LocalMux I__2859 (
            .O(N__14788),
            .I(N__14763));
    InMux I__2858 (
            .O(N__14787),
            .I(N__14756));
    InMux I__2857 (
            .O(N__14786),
            .I(N__14756));
    InMux I__2856 (
            .O(N__14785),
            .I(N__14756));
    LocalMux I__2855 (
            .O(N__14782),
            .I(N__14753));
    InMux I__2854 (
            .O(N__14781),
            .I(N__14750));
    InMux I__2853 (
            .O(N__14778),
            .I(N__14747));
    LocalMux I__2852 (
            .O(N__14769),
            .I(N__14744));
    LocalMux I__2851 (
            .O(N__14766),
            .I(N__14741));
    Span4Mux_v I__2850 (
            .O(N__14763),
            .I(N__14736));
    LocalMux I__2849 (
            .O(N__14756),
            .I(N__14736));
    Span4Mux_v I__2848 (
            .O(N__14753),
            .I(N__14731));
    LocalMux I__2847 (
            .O(N__14750),
            .I(N__14731));
    LocalMux I__2846 (
            .O(N__14747),
            .I(N__14728));
    Span4Mux_v I__2845 (
            .O(N__14744),
            .I(N__14725));
    Span4Mux_v I__2844 (
            .O(N__14741),
            .I(N__14718));
    Span4Mux_v I__2843 (
            .O(N__14736),
            .I(N__14718));
    Span4Mux_v I__2842 (
            .O(N__14731),
            .I(N__14718));
    Span4Mux_v I__2841 (
            .O(N__14728),
            .I(N__14713));
    Span4Mux_h I__2840 (
            .O(N__14725),
            .I(N__14713));
    Span4Mux_h I__2839 (
            .O(N__14718),
            .I(N__14710));
    Odrv4 I__2838 (
            .O(N__14713),
            .I(\b2v_inst.stateZ0Z_7 ));
    Odrv4 I__2837 (
            .O(N__14710),
            .I(\b2v_inst.stateZ0Z_7 ));
    InMux I__2836 (
            .O(N__14705),
            .I(N__14701));
    InMux I__2835 (
            .O(N__14704),
            .I(N__14698));
    LocalMux I__2834 (
            .O(N__14701),
            .I(N__14695));
    LocalMux I__2833 (
            .O(N__14698),
            .I(N__14690));
    Span4Mux_v I__2832 (
            .O(N__14695),
            .I(N__14687));
    InMux I__2831 (
            .O(N__14694),
            .I(N__14684));
    InMux I__2830 (
            .O(N__14693),
            .I(N__14681));
    Span4Mux_h I__2829 (
            .O(N__14690),
            .I(N__14678));
    Span4Mux_h I__2828 (
            .O(N__14687),
            .I(N__14675));
    LocalMux I__2827 (
            .O(N__14684),
            .I(N__14670));
    LocalMux I__2826 (
            .O(N__14681),
            .I(N__14670));
    Odrv4 I__2825 (
            .O(N__14678),
            .I(SYNTHESIZED_WIRE_1_5));
    Odrv4 I__2824 (
            .O(N__14675),
            .I(SYNTHESIZED_WIRE_1_5));
    Odrv12 I__2823 (
            .O(N__14670),
            .I(SYNTHESIZED_WIRE_1_5));
    InMux I__2822 (
            .O(N__14663),
            .I(N__14660));
    LocalMux I__2821 (
            .O(N__14660),
            .I(N__14655));
    InMux I__2820 (
            .O(N__14659),
            .I(N__14652));
    InMux I__2819 (
            .O(N__14658),
            .I(N__14649));
    Span4Mux_v I__2818 (
            .O(N__14655),
            .I(N__14643));
    LocalMux I__2817 (
            .O(N__14652),
            .I(N__14643));
    LocalMux I__2816 (
            .O(N__14649),
            .I(N__14640));
    InMux I__2815 (
            .O(N__14648),
            .I(N__14637));
    Span4Mux_h I__2814 (
            .O(N__14643),
            .I(N__14634));
    Span4Mux_h I__2813 (
            .O(N__14640),
            .I(N__14631));
    LocalMux I__2812 (
            .O(N__14637),
            .I(\b2v_inst.reg_anteriorZ0Z_5 ));
    Odrv4 I__2811 (
            .O(N__14634),
            .I(\b2v_inst.reg_anteriorZ0Z_5 ));
    Odrv4 I__2810 (
            .O(N__14631),
            .I(\b2v_inst.reg_anteriorZ0Z_5 ));
    CascadeMux I__2809 (
            .O(N__14624),
            .I(\b2v_inst.un4_cuenta_ac0_11_0_cascade_ ));
    InMux I__2808 (
            .O(N__14621),
            .I(N__14618));
    LocalMux I__2807 (
            .O(N__14618),
            .I(N__14615));
    Odrv4 I__2806 (
            .O(N__14615),
            .I(\b2v_inst.N_491 ));
    CascadeMux I__2805 (
            .O(N__14612),
            .I(\b2v_inst.cuenta_5_i_o2_0_0_1_cascade_ ));
    CascadeMux I__2804 (
            .O(N__14609),
            .I(\b2v_inst.state_ns_a2_0_o2_1_0_2_cascade_ ));
    InMux I__2803 (
            .O(N__14606),
            .I(N__14602));
    InMux I__2802 (
            .O(N__14605),
            .I(N__14599));
    LocalMux I__2801 (
            .O(N__14602),
            .I(\b2v_inst.cuenta_5_i_o2_0_0_1 ));
    LocalMux I__2800 (
            .O(N__14599),
            .I(\b2v_inst.cuenta_5_i_o2_0_0_1 ));
    CascadeMux I__2799 (
            .O(N__14594),
            .I(\b2v_inst.state_17_rep1_RNICDKZ0Z34_cascade_ ));
    InMux I__2798 (
            .O(N__14591),
            .I(N__14588));
    LocalMux I__2797 (
            .O(N__14588),
            .I(\b2v_inst.cuenta_RNIO2VO3Z0Z_4 ));
    InMux I__2796 (
            .O(N__14585),
            .I(N__14576));
    InMux I__2795 (
            .O(N__14584),
            .I(N__14576));
    InMux I__2794 (
            .O(N__14583),
            .I(N__14576));
    LocalMux I__2793 (
            .O(N__14576),
            .I(\b2v_inst.N_374 ));
    InMux I__2792 (
            .O(N__14573),
            .I(N__14570));
    LocalMux I__2791 (
            .O(N__14570),
            .I(N__14567));
    Span4Mux_h I__2790 (
            .O(N__14567),
            .I(N__14564));
    Odrv4 I__2789 (
            .O(N__14564),
            .I(\b2v_inst1.r_RX_Bytece_0_3 ));
    InMux I__2788 (
            .O(N__14561),
            .I(N__14558));
    LocalMux I__2787 (
            .O(N__14558),
            .I(N__14555));
    Span4Mux_h I__2786 (
            .O(N__14555),
            .I(N__14552));
    Odrv4 I__2785 (
            .O(N__14552),
            .I(\b2v_inst1.r_RX_Bytece_0_0_4 ));
    InMux I__2784 (
            .O(N__14549),
            .I(N__14546));
    LocalMux I__2783 (
            .O(N__14546),
            .I(N__14542));
    InMux I__2782 (
            .O(N__14545),
            .I(N__14539));
    Span4Mux_v I__2781 (
            .O(N__14542),
            .I(N__14536));
    LocalMux I__2780 (
            .O(N__14539),
            .I(N__14533));
    Span4Mux_h I__2779 (
            .O(N__14536),
            .I(N__14530));
    Odrv12 I__2778 (
            .O(N__14533),
            .I(b2v_inst_data_a_escribir_3));
    Odrv4 I__2777 (
            .O(N__14530),
            .I(b2v_inst_data_a_escribir_3));
    InMux I__2776 (
            .O(N__14525),
            .I(N__14522));
    LocalMux I__2775 (
            .O(N__14522),
            .I(N__14519));
    Odrv4 I__2774 (
            .O(N__14519),
            .I(\b2v_inst3.data_to_sendZ0Z_3 ));
    InMux I__2773 (
            .O(N__14516),
            .I(N__14513));
    LocalMux I__2772 (
            .O(N__14513),
            .I(N__14510));
    Span12Mux_v I__2771 (
            .O(N__14510),
            .I(N__14506));
    InMux I__2770 (
            .O(N__14509),
            .I(N__14503));
    Odrv12 I__2769 (
            .O(N__14506),
            .I(b2v_inst_data_a_escribir_4));
    LocalMux I__2768 (
            .O(N__14503),
            .I(b2v_inst_data_a_escribir_4));
    CascadeMux I__2767 (
            .O(N__14498),
            .I(N__14495));
    InMux I__2766 (
            .O(N__14495),
            .I(N__14492));
    LocalMux I__2765 (
            .O(N__14492),
            .I(\b2v_inst3.data_to_sendZ0Z_4 ));
    InMux I__2764 (
            .O(N__14489),
            .I(N__14486));
    LocalMux I__2763 (
            .O(N__14486),
            .I(N__14482));
    InMux I__2762 (
            .O(N__14485),
            .I(N__14479));
    Span4Mux_h I__2761 (
            .O(N__14482),
            .I(N__14476));
    LocalMux I__2760 (
            .O(N__14479),
            .I(N__14473));
    Span4Mux_v I__2759 (
            .O(N__14476),
            .I(N__14470));
    Odrv12 I__2758 (
            .O(N__14473),
            .I(b2v_inst_data_a_escribir_5));
    Odrv4 I__2757 (
            .O(N__14470),
            .I(b2v_inst_data_a_escribir_5));
    CascadeMux I__2756 (
            .O(N__14465),
            .I(N__14462));
    InMux I__2755 (
            .O(N__14462),
            .I(N__14459));
    LocalMux I__2754 (
            .O(N__14459),
            .I(\b2v_inst3.data_to_sendZ0Z_5 ));
    InMux I__2753 (
            .O(N__14456),
            .I(N__14452));
    InMux I__2752 (
            .O(N__14455),
            .I(N__14449));
    LocalMux I__2751 (
            .O(N__14452),
            .I(N__14446));
    LocalMux I__2750 (
            .O(N__14449),
            .I(N__14443));
    Span4Mux_h I__2749 (
            .O(N__14446),
            .I(N__14440));
    Span4Mux_v I__2748 (
            .O(N__14443),
            .I(N__14437));
    Span4Mux_h I__2747 (
            .O(N__14440),
            .I(N__14434));
    Odrv4 I__2746 (
            .O(N__14437),
            .I(b2v_inst_data_a_escribir_6));
    Odrv4 I__2745 (
            .O(N__14434),
            .I(b2v_inst_data_a_escribir_6));
    CascadeMux I__2744 (
            .O(N__14429),
            .I(N__14426));
    InMux I__2743 (
            .O(N__14426),
            .I(N__14423));
    LocalMux I__2742 (
            .O(N__14423),
            .I(\b2v_inst3.data_to_sendZ0Z_6 ));
    InMux I__2741 (
            .O(N__14420),
            .I(N__14410));
    InMux I__2740 (
            .O(N__14419),
            .I(N__14405));
    InMux I__2739 (
            .O(N__14418),
            .I(N__14405));
    InMux I__2738 (
            .O(N__14417),
            .I(N__14394));
    InMux I__2737 (
            .O(N__14416),
            .I(N__14394));
    InMux I__2736 (
            .O(N__14415),
            .I(N__14394));
    InMux I__2735 (
            .O(N__14414),
            .I(N__14394));
    InMux I__2734 (
            .O(N__14413),
            .I(N__14394));
    LocalMux I__2733 (
            .O(N__14410),
            .I(N__14389));
    LocalMux I__2732 (
            .O(N__14405),
            .I(N__14389));
    LocalMux I__2731 (
            .O(N__14394),
            .I(N__14386));
    Span4Mux_v I__2730 (
            .O(N__14389),
            .I(N__14383));
    Span4Mux_v I__2729 (
            .O(N__14386),
            .I(N__14380));
    Odrv4 I__2728 (
            .O(N__14383),
            .I(N_458));
    Odrv4 I__2727 (
            .O(N__14380),
            .I(N_458));
    CascadeMux I__2726 (
            .O(N__14375),
            .I(N__14372));
    InMux I__2725 (
            .O(N__14372),
            .I(N__14368));
    InMux I__2724 (
            .O(N__14371),
            .I(N__14365));
    LocalMux I__2723 (
            .O(N__14368),
            .I(N__14362));
    LocalMux I__2722 (
            .O(N__14365),
            .I(N__14359));
    Span4Mux_h I__2721 (
            .O(N__14362),
            .I(N__14356));
    Span4Mux_h I__2720 (
            .O(N__14359),
            .I(N__14353));
    Odrv4 I__2719 (
            .O(N__14356),
            .I(b2v_inst_data_a_escribir_7));
    Odrv4 I__2718 (
            .O(N__14353),
            .I(b2v_inst_data_a_escribir_7));
    InMux I__2717 (
            .O(N__14348),
            .I(N__14328));
    InMux I__2716 (
            .O(N__14347),
            .I(N__14328));
    InMux I__2715 (
            .O(N__14346),
            .I(N__14328));
    InMux I__2714 (
            .O(N__14345),
            .I(N__14328));
    InMux I__2713 (
            .O(N__14344),
            .I(N__14328));
    InMux I__2712 (
            .O(N__14343),
            .I(N__14323));
    InMux I__2711 (
            .O(N__14342),
            .I(N__14323));
    InMux I__2710 (
            .O(N__14341),
            .I(N__14314));
    InMux I__2709 (
            .O(N__14340),
            .I(N__14314));
    InMux I__2708 (
            .O(N__14339),
            .I(N__14314));
    LocalMux I__2707 (
            .O(N__14328),
            .I(N__14311));
    LocalMux I__2706 (
            .O(N__14323),
            .I(N__14308));
    InMux I__2705 (
            .O(N__14322),
            .I(N__14303));
    InMux I__2704 (
            .O(N__14321),
            .I(N__14303));
    LocalMux I__2703 (
            .O(N__14314),
            .I(N__14300));
    Span4Mux_v I__2702 (
            .O(N__14311),
            .I(N__14295));
    Span4Mux_h I__2701 (
            .O(N__14308),
            .I(N__14292));
    LocalMux I__2700 (
            .O(N__14303),
            .I(N__14287));
    Span12Mux_h I__2699 (
            .O(N__14300),
            .I(N__14287));
    InMux I__2698 (
            .O(N__14299),
            .I(N__14282));
    InMux I__2697 (
            .O(N__14298),
            .I(N__14282));
    Span4Mux_v I__2696 (
            .O(N__14295),
            .I(N__14279));
    Odrv4 I__2695 (
            .O(N__14292),
            .I(N_230));
    Odrv12 I__2694 (
            .O(N__14287),
            .I(N_230));
    LocalMux I__2693 (
            .O(N__14282),
            .I(N_230));
    Odrv4 I__2692 (
            .O(N__14279),
            .I(N_230));
    CascadeMux I__2691 (
            .O(N__14270),
            .I(N__14266));
    InMux I__2690 (
            .O(N__14269),
            .I(N__14261));
    InMux I__2689 (
            .O(N__14266),
            .I(N__14261));
    LocalMux I__2688 (
            .O(N__14261),
            .I(\b2v_inst3.data_to_sendZ0Z_7 ));
    CEMux I__2687 (
            .O(N__14258),
            .I(N__14255));
    LocalMux I__2686 (
            .O(N__14255),
            .I(N__14251));
    CEMux I__2685 (
            .O(N__14254),
            .I(N__14248));
    Odrv12 I__2684 (
            .O(N__14251),
            .I(\b2v_inst3.un2_n_fsm_state_0_sqmuxa_2_0_i_0 ));
    LocalMux I__2683 (
            .O(N__14248),
            .I(\b2v_inst3.un2_n_fsm_state_0_sqmuxa_2_0_i_0 ));
    InMux I__2682 (
            .O(N__14243),
            .I(N__14238));
    InMux I__2681 (
            .O(N__14242),
            .I(N__14235));
    InMux I__2680 (
            .O(N__14241),
            .I(N__14232));
    LocalMux I__2679 (
            .O(N__14238),
            .I(N__14228));
    LocalMux I__2678 (
            .O(N__14235),
            .I(N__14225));
    LocalMux I__2677 (
            .O(N__14232),
            .I(N__14222));
    InMux I__2676 (
            .O(N__14231),
            .I(N__14219));
    Span4Mux_h I__2675 (
            .O(N__14228),
            .I(N__14216));
    Span4Mux_v I__2674 (
            .O(N__14225),
            .I(N__14209));
    Span4Mux_h I__2673 (
            .O(N__14222),
            .I(N__14209));
    LocalMux I__2672 (
            .O(N__14219),
            .I(N__14209));
    Odrv4 I__2671 (
            .O(N__14216),
            .I(SYNTHESIZED_WIRE_1_6));
    Odrv4 I__2670 (
            .O(N__14209),
            .I(SYNTHESIZED_WIRE_1_6));
    InMux I__2669 (
            .O(N__14204),
            .I(N__14201));
    LocalMux I__2668 (
            .O(N__14201),
            .I(N__14195));
    InMux I__2667 (
            .O(N__14200),
            .I(N__14192));
    InMux I__2666 (
            .O(N__14199),
            .I(N__14189));
    InMux I__2665 (
            .O(N__14198),
            .I(N__14186));
    Span4Mux_h I__2664 (
            .O(N__14195),
            .I(N__14181));
    LocalMux I__2663 (
            .O(N__14192),
            .I(N__14181));
    LocalMux I__2662 (
            .O(N__14189),
            .I(N__14178));
    LocalMux I__2661 (
            .O(N__14186),
            .I(\b2v_inst.reg_anteriorZ0Z_6 ));
    Odrv4 I__2660 (
            .O(N__14181),
            .I(\b2v_inst.reg_anteriorZ0Z_6 ));
    Odrv12 I__2659 (
            .O(N__14178),
            .I(\b2v_inst.reg_anteriorZ0Z_6 ));
    CascadeMux I__2658 (
            .O(N__14171),
            .I(\b2v_inst.dir_mem_315_0_cascade_ ));
    InMux I__2657 (
            .O(N__14168),
            .I(N__14165));
    LocalMux I__2656 (
            .O(N__14165),
            .I(\b2v_inst.dir_mem_3Z0Z_1 ));
    InMux I__2655 (
            .O(N__14162),
            .I(N__14159));
    LocalMux I__2654 (
            .O(N__14159),
            .I(\b2v_inst.addr_ram_1_0_iv_i_1_1 ));
    InMux I__2653 (
            .O(N__14156),
            .I(N__14153));
    LocalMux I__2652 (
            .O(N__14153),
            .I(\b2v_inst.dir_mem_3Z0Z_0 ));
    CascadeMux I__2651 (
            .O(N__14150),
            .I(N__14147));
    InMux I__2650 (
            .O(N__14147),
            .I(N__14144));
    LocalMux I__2649 (
            .O(N__14144),
            .I(N__14141));
    Span4Mux_v I__2648 (
            .O(N__14141),
            .I(N__14138));
    Odrv4 I__2647 (
            .O(N__14138),
            .I(\b2v_inst.dir_mem_3Z0Z_5 ));
    InMux I__2646 (
            .O(N__14135),
            .I(N__14132));
    LocalMux I__2645 (
            .O(N__14132),
            .I(N__14129));
    Odrv4 I__2644 (
            .O(N__14129),
            .I(\b2v_inst.dir_mem_3Z0Z_6 ));
    InMux I__2643 (
            .O(N__14126),
            .I(N__14123));
    LocalMux I__2642 (
            .O(N__14123),
            .I(N__14120));
    Span4Mux_v I__2641 (
            .O(N__14120),
            .I(N__14117));
    Span4Mux_h I__2640 (
            .O(N__14117),
            .I(N__14114));
    Odrv4 I__2639 (
            .O(N__14114),
            .I(N_205_i));
    CascadeMux I__2638 (
            .O(N__14111),
            .I(N__14108));
    InMux I__2637 (
            .O(N__14108),
            .I(N__14105));
    LocalMux I__2636 (
            .O(N__14105),
            .I(N__14102));
    Odrv4 I__2635 (
            .O(N__14102),
            .I(\b2v_inst.dir_mem_2Z0Z_6 ));
    CascadeMux I__2634 (
            .O(N__14099),
            .I(\b2v_inst.N_235_cascade_ ));
    InMux I__2633 (
            .O(N__14096),
            .I(N__14089));
    InMux I__2632 (
            .O(N__14095),
            .I(N__14089));
    InMux I__2631 (
            .O(N__14094),
            .I(N__14086));
    LocalMux I__2630 (
            .O(N__14089),
            .I(N__14083));
    LocalMux I__2629 (
            .O(N__14086),
            .I(N__14078));
    Span4Mux_h I__2628 (
            .O(N__14083),
            .I(N__14078));
    Span4Mux_v I__2627 (
            .O(N__14078),
            .I(N__14075));
    Odrv4 I__2626 (
            .O(N__14075),
            .I(\b2v_inst.stateZ0Z_11 ));
    CascadeMux I__2625 (
            .O(N__14072),
            .I(\b2v_inst.N_237_cascade_ ));
    InMux I__2624 (
            .O(N__14069),
            .I(N__14066));
    LocalMux I__2623 (
            .O(N__14066),
            .I(\b2v_inst.addr_ram_1_iv_i_2_0 ));
    CascadeMux I__2622 (
            .O(N__14063),
            .I(\b2v_inst.addr_ram_1_iv_i_1_0_cascade_ ));
    CascadeMux I__2621 (
            .O(N__14060),
            .I(N__14056));
    CascadeMux I__2620 (
            .O(N__14059),
            .I(N__14053));
    InMux I__2619 (
            .O(N__14056),
            .I(N__14050));
    InMux I__2618 (
            .O(N__14053),
            .I(N__14047));
    LocalMux I__2617 (
            .O(N__14050),
            .I(N__14044));
    LocalMux I__2616 (
            .O(N__14047),
            .I(N__14041));
    Span4Mux_v I__2615 (
            .O(N__14044),
            .I(N__14038));
    Odrv4 I__2614 (
            .O(N__14041),
            .I(N_167));
    Odrv4 I__2613 (
            .O(N__14038),
            .I(N_167));
    InMux I__2612 (
            .O(N__14033),
            .I(N__14030));
    LocalMux I__2611 (
            .O(N__14030),
            .I(\b2v_inst.addr_ram_1_0_iv_i_0_1 ));
    CascadeMux I__2610 (
            .O(N__14027),
            .I(N__14023));
    CascadeMux I__2609 (
            .O(N__14026),
            .I(N__14020));
    InMux I__2608 (
            .O(N__14023),
            .I(N__14017));
    InMux I__2607 (
            .O(N__14020),
            .I(N__14014));
    LocalMux I__2606 (
            .O(N__14017),
            .I(N__14011));
    LocalMux I__2605 (
            .O(N__14014),
            .I(N__14006));
    Span4Mux_v I__2604 (
            .O(N__14011),
            .I(N__14006));
    Odrv4 I__2603 (
            .O(N__14006),
            .I(N_60));
    CascadeMux I__2602 (
            .O(N__14003),
            .I(\b2v_inst.addr_ram_1_0_iv_i_0_2_cascade_ ));
    CascadeMux I__2601 (
            .O(N__14000),
            .I(N__13996));
    CascadeMux I__2600 (
            .O(N__13999),
            .I(N__13993));
    InMux I__2599 (
            .O(N__13996),
            .I(N__13990));
    InMux I__2598 (
            .O(N__13993),
            .I(N__13987));
    LocalMux I__2597 (
            .O(N__13990),
            .I(N__13984));
    LocalMux I__2596 (
            .O(N__13987),
            .I(N__13981));
    Span4Mux_h I__2595 (
            .O(N__13984),
            .I(N__13978));
    Odrv4 I__2594 (
            .O(N__13981),
            .I(N_56));
    Odrv4 I__2593 (
            .O(N__13978),
            .I(N_56));
    CascadeMux I__2592 (
            .O(N__13973),
            .I(\b2v_inst.N_236_cascade_ ));
    InMux I__2591 (
            .O(N__13970),
            .I(N__13967));
    LocalMux I__2590 (
            .O(N__13967),
            .I(N__13964));
    Span4Mux_h I__2589 (
            .O(N__13964),
            .I(N__13959));
    InMux I__2588 (
            .O(N__13963),
            .I(N__13954));
    InMux I__2587 (
            .O(N__13962),
            .I(N__13954));
    Odrv4 I__2586 (
            .O(N__13959),
            .I(\b2v_inst.stateZ0Z_9 ));
    LocalMux I__2585 (
            .O(N__13954),
            .I(\b2v_inst.stateZ0Z_9 ));
    CascadeMux I__2584 (
            .O(N__13949),
            .I(\b2v_inst.N_399_cascade_ ));
    InMux I__2583 (
            .O(N__13946),
            .I(N__13943));
    LocalMux I__2582 (
            .O(N__13943),
            .I(\b2v_inst.addr_ram_1_iv_i_1_6 ));
    CascadeMux I__2581 (
            .O(N__13940),
            .I(\b2v_inst.addr_ram_1_iv_i_2_6_cascade_ ));
    CascadeMux I__2580 (
            .O(N__13937),
            .I(N__13933));
    CascadeMux I__2579 (
            .O(N__13936),
            .I(N__13930));
    InMux I__2578 (
            .O(N__13933),
            .I(N__13927));
    InMux I__2577 (
            .O(N__13930),
            .I(N__13924));
    LocalMux I__2576 (
            .O(N__13927),
            .I(N__13919));
    LocalMux I__2575 (
            .O(N__13924),
            .I(N__13919));
    Span4Mux_v I__2574 (
            .O(N__13919),
            .I(N__13916));
    Odrv4 I__2573 (
            .O(N__13916),
            .I(N_165));
    CEMux I__2572 (
            .O(N__13913),
            .I(N__13909));
    CEMux I__2571 (
            .O(N__13912),
            .I(N__13906));
    LocalMux I__2570 (
            .O(N__13909),
            .I(N__13903));
    LocalMux I__2569 (
            .O(N__13906),
            .I(N__13900));
    Span4Mux_h I__2568 (
            .O(N__13903),
            .I(N__13895));
    Span4Mux_h I__2567 (
            .O(N__13900),
            .I(N__13895));
    Span4Mux_h I__2566 (
            .O(N__13895),
            .I(N__13889));
    InMux I__2565 (
            .O(N__13894),
            .I(N__13886));
    InMux I__2564 (
            .O(N__13893),
            .I(N__13881));
    InMux I__2563 (
            .O(N__13892),
            .I(N__13881));
    Odrv4 I__2562 (
            .O(N__13889),
            .I(\b2v_inst.stateZ0Z_12 ));
    LocalMux I__2561 (
            .O(N__13886),
            .I(\b2v_inst.stateZ0Z_12 ));
    LocalMux I__2560 (
            .O(N__13881),
            .I(\b2v_inst.stateZ0Z_12 ));
    CascadeMux I__2559 (
            .O(N__13874),
            .I(\b2v_inst.un2_cuentalto7_3_cascade_ ));
    CascadeMux I__2558 (
            .O(N__13871),
            .I(\b2v_inst.N_351_0_cascade_ ));
    CascadeMux I__2557 (
            .O(N__13868),
            .I(N__13864));
    InMux I__2556 (
            .O(N__13867),
            .I(N__13861));
    InMux I__2555 (
            .O(N__13864),
            .I(N__13858));
    LocalMux I__2554 (
            .O(N__13861),
            .I(\b2v_inst.cuenta_fastZ0Z_4 ));
    LocalMux I__2553 (
            .O(N__13858),
            .I(\b2v_inst.cuenta_fastZ0Z_4 ));
    InMux I__2552 (
            .O(N__13853),
            .I(N__13848));
    InMux I__2551 (
            .O(N__13852),
            .I(N__13845));
    InMux I__2550 (
            .O(N__13851),
            .I(N__13842));
    LocalMux I__2549 (
            .O(N__13848),
            .I(\b2v_inst.cuenta_RNIQ56K_0Z0Z_3 ));
    LocalMux I__2548 (
            .O(N__13845),
            .I(\b2v_inst.cuenta_RNIQ56K_0Z0Z_3 ));
    LocalMux I__2547 (
            .O(N__13842),
            .I(\b2v_inst.cuenta_RNIQ56K_0Z0Z_3 ));
    InMux I__2546 (
            .O(N__13835),
            .I(N__13832));
    LocalMux I__2545 (
            .O(N__13832),
            .I(\b2v_inst.N_376_1 ));
    InMux I__2544 (
            .O(N__13829),
            .I(N__13823));
    InMux I__2543 (
            .O(N__13828),
            .I(N__13823));
    LocalMux I__2542 (
            .O(N__13823),
            .I(\b2v_inst.cuenta_RNIQI4FZ0Z_2 ));
    CascadeMux I__2541 (
            .O(N__13820),
            .I(N__13817));
    InMux I__2540 (
            .O(N__13817),
            .I(N__13811));
    InMux I__2539 (
            .O(N__13816),
            .I(N__13811));
    LocalMux I__2538 (
            .O(N__13811),
            .I(\b2v_inst.cuenta_RNIR03AZ0Z_1 ));
    CascadeMux I__2537 (
            .O(N__13808),
            .I(\b2v_inst.N_376_1_cascade_ ));
    CascadeMux I__2536 (
            .O(N__13805),
            .I(N__13797));
    InMux I__2535 (
            .O(N__13804),
            .I(N__13793));
    InMux I__2534 (
            .O(N__13803),
            .I(N__13790));
    InMux I__2533 (
            .O(N__13802),
            .I(N__13787));
    InMux I__2532 (
            .O(N__13801),
            .I(N__13778));
    InMux I__2531 (
            .O(N__13800),
            .I(N__13778));
    InMux I__2530 (
            .O(N__13797),
            .I(N__13778));
    InMux I__2529 (
            .O(N__13796),
            .I(N__13778));
    LocalMux I__2528 (
            .O(N__13793),
            .I(\b2v_inst.cuentaZ0Z_1 ));
    LocalMux I__2527 (
            .O(N__13790),
            .I(\b2v_inst.cuentaZ0Z_1 ));
    LocalMux I__2526 (
            .O(N__13787),
            .I(\b2v_inst.cuentaZ0Z_1 ));
    LocalMux I__2525 (
            .O(N__13778),
            .I(\b2v_inst.cuentaZ0Z_1 ));
    InMux I__2524 (
            .O(N__13769),
            .I(N__13766));
    LocalMux I__2523 (
            .O(N__13766),
            .I(N__13763));
    Odrv4 I__2522 (
            .O(N__13763),
            .I(\b2v_inst.cuenta_5_i_a2_0_3 ));
    InMux I__2521 (
            .O(N__13760),
            .I(N__13754));
    InMux I__2520 (
            .O(N__13759),
            .I(N__13751));
    InMux I__2519 (
            .O(N__13758),
            .I(N__13746));
    InMux I__2518 (
            .O(N__13757),
            .I(N__13746));
    LocalMux I__2517 (
            .O(N__13754),
            .I(N__13734));
    LocalMux I__2516 (
            .O(N__13751),
            .I(N__13734));
    LocalMux I__2515 (
            .O(N__13746),
            .I(N__13734));
    InMux I__2514 (
            .O(N__13745),
            .I(N__13723));
    InMux I__2513 (
            .O(N__13744),
            .I(N__13723));
    InMux I__2512 (
            .O(N__13743),
            .I(N__13723));
    InMux I__2511 (
            .O(N__13742),
            .I(N__13723));
    InMux I__2510 (
            .O(N__13741),
            .I(N__13723));
    Odrv4 I__2509 (
            .O(N__13734),
            .I(\b2v_inst.cuentaZ0Z_0 ));
    LocalMux I__2508 (
            .O(N__13723),
            .I(\b2v_inst.cuentaZ0Z_0 ));
    InMux I__2507 (
            .O(N__13718),
            .I(N__13715));
    LocalMux I__2506 (
            .O(N__13715),
            .I(\b2v_inst.N_377 ));
    CascadeMux I__2505 (
            .O(N__13712),
            .I(\b2v_inst.N_491_cascade_ ));
    InMux I__2504 (
            .O(N__13709),
            .I(N__13706));
    LocalMux I__2503 (
            .O(N__13706),
            .I(N__13703));
    Span4Mux_h I__2502 (
            .O(N__13703),
            .I(N__13700));
    Odrv4 I__2501 (
            .O(N__13700),
            .I(\b2v_inst.state_RNIFQKOZ0Z_17 ));
    CascadeMux I__2500 (
            .O(N__13697),
            .I(\b2v_inst.state_RNIFQKOZ0Z_17_cascade_ ));
    CascadeMux I__2499 (
            .O(N__13694),
            .I(\b2v_inst.cuenta_5_i_a2_2_0_1_cascade_ ));
    CascadeMux I__2498 (
            .O(N__13691),
            .I(\b2v_inst.un4_cuenta_c4_cascade_ ));
    CascadeMux I__2497 (
            .O(N__13688),
            .I(N__13683));
    InMux I__2496 (
            .O(N__13687),
            .I(N__13680));
    InMux I__2495 (
            .O(N__13686),
            .I(N__13675));
    InMux I__2494 (
            .O(N__13683),
            .I(N__13675));
    LocalMux I__2493 (
            .O(N__13680),
            .I(\b2v_inst.cuentaZ0Z_3 ));
    LocalMux I__2492 (
            .O(N__13675),
            .I(\b2v_inst.cuentaZ0Z_3 ));
    InMux I__2491 (
            .O(N__13670),
            .I(N__13662));
    InMux I__2490 (
            .O(N__13669),
            .I(N__13659));
    InMux I__2489 (
            .O(N__13668),
            .I(N__13650));
    InMux I__2488 (
            .O(N__13667),
            .I(N__13650));
    InMux I__2487 (
            .O(N__13666),
            .I(N__13650));
    InMux I__2486 (
            .O(N__13665),
            .I(N__13650));
    LocalMux I__2485 (
            .O(N__13662),
            .I(\b2v_inst.cuentaZ0Z_2 ));
    LocalMux I__2484 (
            .O(N__13659),
            .I(\b2v_inst.cuentaZ0Z_2 ));
    LocalMux I__2483 (
            .O(N__13650),
            .I(\b2v_inst.cuentaZ0Z_2 ));
    InMux I__2482 (
            .O(N__13643),
            .I(N__13639));
    InMux I__2481 (
            .O(N__13642),
            .I(N__13635));
    LocalMux I__2480 (
            .O(N__13639),
            .I(N__13632));
    InMux I__2479 (
            .O(N__13638),
            .I(N__13629));
    LocalMux I__2478 (
            .O(N__13635),
            .I(N__13626));
    Span4Mux_v I__2477 (
            .O(N__13632),
            .I(N__13623));
    LocalMux I__2476 (
            .O(N__13629),
            .I(N__13620));
    Span4Mux_v I__2475 (
            .O(N__13626),
            .I(N__13612));
    Span4Mux_h I__2474 (
            .O(N__13623),
            .I(N__13612));
    Span4Mux_h I__2473 (
            .O(N__13620),
            .I(N__13612));
    InMux I__2472 (
            .O(N__13619),
            .I(N__13609));
    Odrv4 I__2471 (
            .O(N__13612),
            .I(SYNTHESIZED_WIRE_1_7));
    LocalMux I__2470 (
            .O(N__13609),
            .I(SYNTHESIZED_WIRE_1_7));
    InMux I__2469 (
            .O(N__13604),
            .I(N__13598));
    CascadeMux I__2468 (
            .O(N__13603),
            .I(N__13595));
    InMux I__2467 (
            .O(N__13602),
            .I(N__13592));
    InMux I__2466 (
            .O(N__13601),
            .I(N__13589));
    LocalMux I__2465 (
            .O(N__13598),
            .I(N__13586));
    InMux I__2464 (
            .O(N__13595),
            .I(N__13583));
    LocalMux I__2463 (
            .O(N__13592),
            .I(N__13578));
    LocalMux I__2462 (
            .O(N__13589),
            .I(N__13578));
    Span4Mux_h I__2461 (
            .O(N__13586),
            .I(N__13575));
    LocalMux I__2460 (
            .O(N__13583),
            .I(\b2v_inst.reg_anteriorZ0Z_7 ));
    Odrv4 I__2459 (
            .O(N__13578),
            .I(\b2v_inst.reg_anteriorZ0Z_7 ));
    Odrv4 I__2458 (
            .O(N__13575),
            .I(\b2v_inst.reg_anteriorZ0Z_7 ));
    InMux I__2457 (
            .O(N__13568),
            .I(N__13565));
    LocalMux I__2456 (
            .O(N__13565),
            .I(N__13562));
    Span4Mux_h I__2455 (
            .O(N__13562),
            .I(N__13559));
    Span4Mux_v I__2454 (
            .O(N__13559),
            .I(N__13556));
    Odrv4 I__2453 (
            .O(N__13556),
            .I(\b2v_inst.data_a_escribir9_7_and ));
    InMux I__2452 (
            .O(N__13553),
            .I(N__13549));
    InMux I__2451 (
            .O(N__13552),
            .I(N__13546));
    LocalMux I__2450 (
            .O(N__13549),
            .I(N__13542));
    LocalMux I__2449 (
            .O(N__13546),
            .I(N__13539));
    InMux I__2448 (
            .O(N__13545),
            .I(N__13536));
    Span4Mux_h I__2447 (
            .O(N__13542),
            .I(N__13532));
    Span12Mux_h I__2446 (
            .O(N__13539),
            .I(N__13529));
    LocalMux I__2445 (
            .O(N__13536),
            .I(N__13526));
    InMux I__2444 (
            .O(N__13535),
            .I(N__13523));
    Odrv4 I__2443 (
            .O(N__13532),
            .I(SYNTHESIZED_WIRE_1_4));
    Odrv12 I__2442 (
            .O(N__13529),
            .I(SYNTHESIZED_WIRE_1_4));
    Odrv12 I__2441 (
            .O(N__13526),
            .I(SYNTHESIZED_WIRE_1_4));
    LocalMux I__2440 (
            .O(N__13523),
            .I(SYNTHESIZED_WIRE_1_4));
    InMux I__2439 (
            .O(N__13514),
            .I(N__13510));
    InMux I__2438 (
            .O(N__13513),
            .I(N__13505));
    LocalMux I__2437 (
            .O(N__13510),
            .I(N__13502));
    InMux I__2436 (
            .O(N__13509),
            .I(N__13499));
    InMux I__2435 (
            .O(N__13508),
            .I(N__13496));
    LocalMux I__2434 (
            .O(N__13505),
            .I(N__13493));
    Span4Mux_v I__2433 (
            .O(N__13502),
            .I(N__13488));
    LocalMux I__2432 (
            .O(N__13499),
            .I(N__13488));
    LocalMux I__2431 (
            .O(N__13496),
            .I(\b2v_inst.reg_anteriorZ0Z_4 ));
    Odrv4 I__2430 (
            .O(N__13493),
            .I(\b2v_inst.reg_anteriorZ0Z_4 ));
    Odrv4 I__2429 (
            .O(N__13488),
            .I(\b2v_inst.reg_anteriorZ0Z_4 ));
    InMux I__2428 (
            .O(N__13481),
            .I(N__13477));
    CascadeMux I__2427 (
            .O(N__13480),
            .I(N__13474));
    LocalMux I__2426 (
            .O(N__13477),
            .I(N__13471));
    InMux I__2425 (
            .O(N__13474),
            .I(N__13468));
    Span4Mux_h I__2424 (
            .O(N__13471),
            .I(N__13463));
    LocalMux I__2423 (
            .O(N__13468),
            .I(N__13463));
    Odrv4 I__2422 (
            .O(N__13463),
            .I(b2v_inst_data_a_escribir_1));
    InMux I__2421 (
            .O(N__13460),
            .I(N__13456));
    CascadeMux I__2420 (
            .O(N__13459),
            .I(N__13453));
    LocalMux I__2419 (
            .O(N__13456),
            .I(N__13450));
    InMux I__2418 (
            .O(N__13453),
            .I(N__13447));
    Span4Mux_v I__2417 (
            .O(N__13450),
            .I(N__13444));
    LocalMux I__2416 (
            .O(N__13447),
            .I(N__13441));
    Odrv4 I__2415 (
            .O(N__13444),
            .I(b2v_inst_data_a_escribir_0));
    Odrv4 I__2414 (
            .O(N__13441),
            .I(b2v_inst_data_a_escribir_0));
    CascadeMux I__2413 (
            .O(N__13436),
            .I(N__13433));
    InMux I__2412 (
            .O(N__13433),
            .I(N__13430));
    LocalMux I__2411 (
            .O(N__13430),
            .I(\b2v_inst3.data_to_sendZ0Z_1 ));
    InMux I__2410 (
            .O(N__13427),
            .I(N__13424));
    LocalMux I__2409 (
            .O(N__13424),
            .I(N__13421));
    Span12Mux_v I__2408 (
            .O(N__13421),
            .I(N__13418));
    Odrv12 I__2407 (
            .O(N__13418),
            .I(\b2v_inst3.data_to_sendZ0Z_0 ));
    CascadeMux I__2406 (
            .O(N__13415),
            .I(N__13412));
    InMux I__2405 (
            .O(N__13412),
            .I(N__13408));
    InMux I__2404 (
            .O(N__13411),
            .I(N__13405));
    LocalMux I__2403 (
            .O(N__13408),
            .I(N__13402));
    LocalMux I__2402 (
            .O(N__13405),
            .I(N__13399));
    Span4Mux_h I__2401 (
            .O(N__13402),
            .I(N__13394));
    Span4Mux_h I__2400 (
            .O(N__13399),
            .I(N__13394));
    Odrv4 I__2399 (
            .O(N__13394),
            .I(b2v_inst_data_a_escribir_2));
    CascadeMux I__2398 (
            .O(N__13391),
            .I(N__13388));
    InMux I__2397 (
            .O(N__13388),
            .I(N__13385));
    LocalMux I__2396 (
            .O(N__13385),
            .I(\b2v_inst3.data_to_sendZ0Z_2 ));
    CascadeMux I__2395 (
            .O(N__13382),
            .I(N__13376));
    InMux I__2394 (
            .O(N__13381),
            .I(N__13373));
    InMux I__2393 (
            .O(N__13380),
            .I(N__13370));
    InMux I__2392 (
            .O(N__13379),
            .I(N__13365));
    InMux I__2391 (
            .O(N__13376),
            .I(N__13365));
    LocalMux I__2390 (
            .O(N__13373),
            .I(\b2v_inst3.fsm_state_RNIEPSN1Z0Z_0 ));
    LocalMux I__2389 (
            .O(N__13370),
            .I(\b2v_inst3.fsm_state_RNIEPSN1Z0Z_0 ));
    LocalMux I__2388 (
            .O(N__13365),
            .I(\b2v_inst3.fsm_state_RNIEPSN1Z0Z_0 ));
    InMux I__2387 (
            .O(N__13358),
            .I(N__13352));
    InMux I__2386 (
            .O(N__13357),
            .I(N__13344));
    InMux I__2385 (
            .O(N__13356),
            .I(N__13339));
    InMux I__2384 (
            .O(N__13355),
            .I(N__13339));
    LocalMux I__2383 (
            .O(N__13352),
            .I(N__13336));
    InMux I__2382 (
            .O(N__13351),
            .I(N__13333));
    InMux I__2381 (
            .O(N__13350),
            .I(N__13330));
    InMux I__2380 (
            .O(N__13349),
            .I(N__13325));
    InMux I__2379 (
            .O(N__13348),
            .I(N__13325));
    InMux I__2378 (
            .O(N__13347),
            .I(N__13322));
    LocalMux I__2377 (
            .O(N__13344),
            .I(N__13317));
    LocalMux I__2376 (
            .O(N__13339),
            .I(N__13317));
    Odrv4 I__2375 (
            .O(N__13336),
            .I(\b2v_inst3.N_105_7 ));
    LocalMux I__2374 (
            .O(N__13333),
            .I(\b2v_inst3.N_105_7 ));
    LocalMux I__2373 (
            .O(N__13330),
            .I(\b2v_inst3.N_105_7 ));
    LocalMux I__2372 (
            .O(N__13325),
            .I(\b2v_inst3.N_105_7 ));
    LocalMux I__2371 (
            .O(N__13322),
            .I(\b2v_inst3.N_105_7 ));
    Odrv4 I__2370 (
            .O(N__13317),
            .I(\b2v_inst3.N_105_7 ));
    InMux I__2369 (
            .O(N__13304),
            .I(N__13297));
    InMux I__2368 (
            .O(N__13303),
            .I(N__13294));
    InMux I__2367 (
            .O(N__13302),
            .I(N__13287));
    InMux I__2366 (
            .O(N__13301),
            .I(N__13287));
    InMux I__2365 (
            .O(N__13300),
            .I(N__13287));
    LocalMux I__2364 (
            .O(N__13297),
            .I(\b2v_inst3.bit_counterZ0Z_0 ));
    LocalMux I__2363 (
            .O(N__13294),
            .I(\b2v_inst3.bit_counterZ0Z_0 ));
    LocalMux I__2362 (
            .O(N__13287),
            .I(\b2v_inst3.bit_counterZ0Z_0 ));
    CascadeMux I__2361 (
            .O(N__13280),
            .I(N__13277));
    InMux I__2360 (
            .O(N__13277),
            .I(N__13274));
    LocalMux I__2359 (
            .O(N__13274),
            .I(\b2v_inst.state_ns_a2_0_a2_0_1_2 ));
    CascadeMux I__2358 (
            .O(N__13271),
            .I(N__13268));
    InMux I__2357 (
            .O(N__13268),
            .I(N__13263));
    CascadeMux I__2356 (
            .O(N__13267),
            .I(N__13260));
    CascadeMux I__2355 (
            .O(N__13266),
            .I(N__13257));
    LocalMux I__2354 (
            .O(N__13263),
            .I(N__13254));
    InMux I__2353 (
            .O(N__13260),
            .I(N__13251));
    InMux I__2352 (
            .O(N__13257),
            .I(N__13248));
    Odrv4 I__2351 (
            .O(N__13254),
            .I(\b2v_inst.reg_ancho_3_i_7 ));
    LocalMux I__2350 (
            .O(N__13251),
            .I(\b2v_inst.reg_ancho_3_i_7 ));
    LocalMux I__2349 (
            .O(N__13248),
            .I(\b2v_inst.reg_ancho_3_i_7 ));
    InMux I__2348 (
            .O(N__13241),
            .I(bfn_6_18_0_));
    CascadeMux I__2347 (
            .O(N__13238),
            .I(N__13234));
    InMux I__2346 (
            .O(N__13237),
            .I(N__13224));
    InMux I__2345 (
            .O(N__13234),
            .I(N__13220));
    InMux I__2344 (
            .O(N__13233),
            .I(N__13215));
    InMux I__2343 (
            .O(N__13232),
            .I(N__13210));
    InMux I__2342 (
            .O(N__13231),
            .I(N__13210));
    InMux I__2341 (
            .O(N__13230),
            .I(N__13207));
    InMux I__2340 (
            .O(N__13229),
            .I(N__13204));
    InMux I__2339 (
            .O(N__13228),
            .I(N__13199));
    InMux I__2338 (
            .O(N__13227),
            .I(N__13199));
    LocalMux I__2337 (
            .O(N__13224),
            .I(N__13196));
    InMux I__2336 (
            .O(N__13223),
            .I(N__13193));
    LocalMux I__2335 (
            .O(N__13220),
            .I(N__13190));
    InMux I__2334 (
            .O(N__13219),
            .I(N__13185));
    InMux I__2333 (
            .O(N__13218),
            .I(N__13185));
    LocalMux I__2332 (
            .O(N__13215),
            .I(N__13180));
    LocalMux I__2331 (
            .O(N__13210),
            .I(N__13180));
    LocalMux I__2330 (
            .O(N__13207),
            .I(N__13173));
    LocalMux I__2329 (
            .O(N__13204),
            .I(N__13173));
    LocalMux I__2328 (
            .O(N__13199),
            .I(N__13173));
    Span4Mux_v I__2327 (
            .O(N__13196),
            .I(N__13170));
    LocalMux I__2326 (
            .O(N__13193),
            .I(N__13163));
    Span12Mux_s8_v I__2325 (
            .O(N__13190),
            .I(N__13163));
    LocalMux I__2324 (
            .O(N__13185),
            .I(N__13163));
    Span4Mux_h I__2323 (
            .O(N__13180),
            .I(N__13158));
    Span4Mux_h I__2322 (
            .O(N__13173),
            .I(N__13158));
    Odrv4 I__2321 (
            .O(N__13170),
            .I(\b2v_inst.un3_valor_max2_THRU_CO ));
    Odrv12 I__2320 (
            .O(N__13163),
            .I(\b2v_inst.un3_valor_max2_THRU_CO ));
    Odrv4 I__2319 (
            .O(N__13158),
            .I(\b2v_inst.un3_valor_max2_THRU_CO ));
    IoInMux I__2318 (
            .O(N__13151),
            .I(N__13148));
    LocalMux I__2317 (
            .O(N__13148),
            .I(N__13145));
    Span4Mux_s2_h I__2316 (
            .O(N__13145),
            .I(N__13142));
    Sp12to4 I__2315 (
            .O(N__13142),
            .I(N__13138));
    InMux I__2314 (
            .O(N__13141),
            .I(N__13135));
    Span12Mux_v I__2313 (
            .O(N__13138),
            .I(N__13130));
    LocalMux I__2312 (
            .O(N__13135),
            .I(N__13130));
    Odrv12 I__2311 (
            .O(N__13130),
            .I(reset_i));
    InMux I__2310 (
            .O(N__13127),
            .I(N__13124));
    LocalMux I__2309 (
            .O(N__13124),
            .I(N__13121));
    Span4Mux_v I__2308 (
            .O(N__13121),
            .I(N__13118));
    Odrv4 I__2307 (
            .O(N__13118),
            .I(\b2v_inst3.un2_n_fsm_state_0_sqmuxa_2_0_i ));
    InMux I__2306 (
            .O(N__13115),
            .I(N__13112));
    LocalMux I__2305 (
            .O(N__13112),
            .I(N__13109));
    Span4Mux_h I__2304 (
            .O(N__13109),
            .I(N__13106));
    Odrv4 I__2303 (
            .O(N__13106),
            .I(\b2v_inst1.r_RX_Bytece_0_6 ));
    InMux I__2302 (
            .O(N__13103),
            .I(N__13099));
    InMux I__2301 (
            .O(N__13102),
            .I(N__13096));
    LocalMux I__2300 (
            .O(N__13099),
            .I(N__13092));
    LocalMux I__2299 (
            .O(N__13096),
            .I(N__13089));
    InMux I__2298 (
            .O(N__13095),
            .I(N__13086));
    Span4Mux_h I__2297 (
            .O(N__13092),
            .I(N__13080));
    Span4Mux_h I__2296 (
            .O(N__13089),
            .I(N__13080));
    LocalMux I__2295 (
            .O(N__13086),
            .I(N__13077));
    InMux I__2294 (
            .O(N__13085),
            .I(N__13074));
    Odrv4 I__2293 (
            .O(N__13080),
            .I(SYNTHESIZED_WIRE_1_0));
    Odrv4 I__2292 (
            .O(N__13077),
            .I(SYNTHESIZED_WIRE_1_0));
    LocalMux I__2291 (
            .O(N__13074),
            .I(SYNTHESIZED_WIRE_1_0));
    InMux I__2290 (
            .O(N__13067),
            .I(N__13064));
    LocalMux I__2289 (
            .O(N__13064),
            .I(N__13061));
    Span4Mux_v I__2288 (
            .O(N__13061),
            .I(N__13055));
    InMux I__2287 (
            .O(N__13060),
            .I(N__13052));
    InMux I__2286 (
            .O(N__13059),
            .I(N__13049));
    InMux I__2285 (
            .O(N__13058),
            .I(N__13046));
    Span4Mux_h I__2284 (
            .O(N__13055),
            .I(N__13041));
    LocalMux I__2283 (
            .O(N__13052),
            .I(N__13041));
    LocalMux I__2282 (
            .O(N__13049),
            .I(N__13038));
    LocalMux I__2281 (
            .O(N__13046),
            .I(\b2v_inst.reg_anteriorZ0Z_0 ));
    Odrv4 I__2280 (
            .O(N__13041),
            .I(\b2v_inst.reg_anteriorZ0Z_0 ));
    Odrv12 I__2279 (
            .O(N__13038),
            .I(\b2v_inst.reg_anteriorZ0Z_0 ));
    InMux I__2278 (
            .O(N__13031),
            .I(N__13028));
    LocalMux I__2277 (
            .O(N__13028),
            .I(N__13024));
    InMux I__2276 (
            .O(N__13027),
            .I(N__13021));
    Span4Mux_h I__2275 (
            .O(N__13024),
            .I(N__13017));
    LocalMux I__2274 (
            .O(N__13021),
            .I(N__13014));
    InMux I__2273 (
            .O(N__13020),
            .I(N__13011));
    Span4Mux_v I__2272 (
            .O(N__13017),
            .I(N__13005));
    Span4Mux_h I__2271 (
            .O(N__13014),
            .I(N__13005));
    LocalMux I__2270 (
            .O(N__13011),
            .I(N__13002));
    InMux I__2269 (
            .O(N__13010),
            .I(N__12999));
    Odrv4 I__2268 (
            .O(N__13005),
            .I(SYNTHESIZED_WIRE_1_1));
    Odrv4 I__2267 (
            .O(N__13002),
            .I(SYNTHESIZED_WIRE_1_1));
    LocalMux I__2266 (
            .O(N__12999),
            .I(SYNTHESIZED_WIRE_1_1));
    InMux I__2265 (
            .O(N__12992),
            .I(N__12988));
    InMux I__2264 (
            .O(N__12991),
            .I(N__12983));
    LocalMux I__2263 (
            .O(N__12988),
            .I(N__12980));
    InMux I__2262 (
            .O(N__12987),
            .I(N__12977));
    InMux I__2261 (
            .O(N__12986),
            .I(N__12974));
    LocalMux I__2260 (
            .O(N__12983),
            .I(N__12971));
    Span4Mux_v I__2259 (
            .O(N__12980),
            .I(N__12966));
    LocalMux I__2258 (
            .O(N__12977),
            .I(N__12966));
    LocalMux I__2257 (
            .O(N__12974),
            .I(\b2v_inst.reg_anteriorZ0Z_1 ));
    Odrv4 I__2256 (
            .O(N__12971),
            .I(\b2v_inst.reg_anteriorZ0Z_1 ));
    Odrv4 I__2255 (
            .O(N__12966),
            .I(\b2v_inst.reg_anteriorZ0Z_1 ));
    InMux I__2254 (
            .O(N__12959),
            .I(N__12955));
    InMux I__2253 (
            .O(N__12958),
            .I(N__12952));
    LocalMux I__2252 (
            .O(N__12955),
            .I(N__12948));
    LocalMux I__2251 (
            .O(N__12952),
            .I(N__12945));
    InMux I__2250 (
            .O(N__12951),
            .I(N__12942));
    Span4Mux_h I__2249 (
            .O(N__12948),
            .I(N__12936));
    Span4Mux_h I__2248 (
            .O(N__12945),
            .I(N__12936));
    LocalMux I__2247 (
            .O(N__12942),
            .I(N__12933));
    InMux I__2246 (
            .O(N__12941),
            .I(N__12930));
    Odrv4 I__2245 (
            .O(N__12936),
            .I(SYNTHESIZED_WIRE_1_2));
    Odrv12 I__2244 (
            .O(N__12933),
            .I(SYNTHESIZED_WIRE_1_2));
    LocalMux I__2243 (
            .O(N__12930),
            .I(SYNTHESIZED_WIRE_1_2));
    CascadeMux I__2242 (
            .O(N__12923),
            .I(N__12920));
    InMux I__2241 (
            .O(N__12920),
            .I(N__12916));
    InMux I__2240 (
            .O(N__12919),
            .I(N__12911));
    LocalMux I__2239 (
            .O(N__12916),
            .I(N__12908));
    InMux I__2238 (
            .O(N__12915),
            .I(N__12905));
    InMux I__2237 (
            .O(N__12914),
            .I(N__12902));
    LocalMux I__2236 (
            .O(N__12911),
            .I(N__12899));
    Span4Mux_v I__2235 (
            .O(N__12908),
            .I(N__12894));
    LocalMux I__2234 (
            .O(N__12905),
            .I(N__12894));
    LocalMux I__2233 (
            .O(N__12902),
            .I(\b2v_inst.reg_anteriorZ0Z_2 ));
    Odrv4 I__2232 (
            .O(N__12899),
            .I(\b2v_inst.reg_anteriorZ0Z_2 ));
    Odrv4 I__2231 (
            .O(N__12894),
            .I(\b2v_inst.reg_anteriorZ0Z_2 ));
    InMux I__2230 (
            .O(N__12887),
            .I(N__12883));
    InMux I__2229 (
            .O(N__12886),
            .I(N__12880));
    LocalMux I__2228 (
            .O(N__12883),
            .I(N__12876));
    LocalMux I__2227 (
            .O(N__12880),
            .I(N__12873));
    InMux I__2226 (
            .O(N__12879),
            .I(N__12870));
    Span4Mux_h I__2225 (
            .O(N__12876),
            .I(N__12864));
    Span4Mux_h I__2224 (
            .O(N__12873),
            .I(N__12864));
    LocalMux I__2223 (
            .O(N__12870),
            .I(N__12861));
    InMux I__2222 (
            .O(N__12869),
            .I(N__12858));
    Odrv4 I__2221 (
            .O(N__12864),
            .I(SYNTHESIZED_WIRE_1_3));
    Odrv4 I__2220 (
            .O(N__12861),
            .I(SYNTHESIZED_WIRE_1_3));
    LocalMux I__2219 (
            .O(N__12858),
            .I(SYNTHESIZED_WIRE_1_3));
    InMux I__2218 (
            .O(N__12851),
            .I(N__12848));
    LocalMux I__2217 (
            .O(N__12848),
            .I(N__12842));
    CascadeMux I__2216 (
            .O(N__12847),
            .I(N__12839));
    InMux I__2215 (
            .O(N__12846),
            .I(N__12836));
    InMux I__2214 (
            .O(N__12845),
            .I(N__12833));
    Span4Mux_h I__2213 (
            .O(N__12842),
            .I(N__12830));
    InMux I__2212 (
            .O(N__12839),
            .I(N__12827));
    LocalMux I__2211 (
            .O(N__12836),
            .I(N__12824));
    LocalMux I__2210 (
            .O(N__12833),
            .I(N__12821));
    Odrv4 I__2209 (
            .O(N__12830),
            .I(\b2v_inst.reg_anteriorZ0Z_3 ));
    LocalMux I__2208 (
            .O(N__12827),
            .I(\b2v_inst.reg_anteriorZ0Z_3 ));
    Odrv4 I__2207 (
            .O(N__12824),
            .I(\b2v_inst.reg_anteriorZ0Z_3 ));
    Odrv4 I__2206 (
            .O(N__12821),
            .I(\b2v_inst.reg_anteriorZ0Z_3 ));
    InMux I__2205 (
            .O(N__12812),
            .I(N__12809));
    LocalMux I__2204 (
            .O(N__12809),
            .I(N__12804));
    InMux I__2203 (
            .O(N__12808),
            .I(N__12801));
    InMux I__2202 (
            .O(N__12807),
            .I(N__12798));
    Odrv12 I__2201 (
            .O(N__12804),
            .I(\b2v_inst.reg_ancho_3Z0Z_6 ));
    LocalMux I__2200 (
            .O(N__12801),
            .I(\b2v_inst.reg_ancho_3Z0Z_6 ));
    LocalMux I__2199 (
            .O(N__12798),
            .I(\b2v_inst.reg_ancho_3Z0Z_6 ));
    InMux I__2198 (
            .O(N__12791),
            .I(N__12788));
    LocalMux I__2197 (
            .O(N__12788),
            .I(N__12785));
    Span4Mux_h I__2196 (
            .O(N__12785),
            .I(N__12780));
    InMux I__2195 (
            .O(N__12784),
            .I(N__12777));
    InMux I__2194 (
            .O(N__12783),
            .I(N__12774));
    Odrv4 I__2193 (
            .O(N__12780),
            .I(\b2v_inst.reg_ancho_3Z0Z_5 ));
    LocalMux I__2192 (
            .O(N__12777),
            .I(\b2v_inst.reg_ancho_3Z0Z_5 ));
    LocalMux I__2191 (
            .O(N__12774),
            .I(\b2v_inst.reg_ancho_3Z0Z_5 ));
    CascadeMux I__2190 (
            .O(N__12767),
            .I(N__12764));
    InMux I__2189 (
            .O(N__12764),
            .I(N__12759));
    CascadeMux I__2188 (
            .O(N__12763),
            .I(N__12756));
    CascadeMux I__2187 (
            .O(N__12762),
            .I(N__12753));
    LocalMux I__2186 (
            .O(N__12759),
            .I(N__12750));
    InMux I__2185 (
            .O(N__12756),
            .I(N__12747));
    InMux I__2184 (
            .O(N__12753),
            .I(N__12744));
    Odrv4 I__2183 (
            .O(N__12750),
            .I(\b2v_inst.reg_ancho_3_i_0 ));
    LocalMux I__2182 (
            .O(N__12747),
            .I(\b2v_inst.reg_ancho_3_i_0 ));
    LocalMux I__2181 (
            .O(N__12744),
            .I(\b2v_inst.reg_ancho_3_i_0 ));
    CascadeMux I__2180 (
            .O(N__12737),
            .I(N__12732));
    CascadeMux I__2179 (
            .O(N__12736),
            .I(N__12729));
    CascadeMux I__2178 (
            .O(N__12735),
            .I(N__12726));
    InMux I__2177 (
            .O(N__12732),
            .I(N__12723));
    InMux I__2176 (
            .O(N__12729),
            .I(N__12720));
    InMux I__2175 (
            .O(N__12726),
            .I(N__12717));
    LocalMux I__2174 (
            .O(N__12723),
            .I(N__12714));
    LocalMux I__2173 (
            .O(N__12720),
            .I(\b2v_inst.reg_ancho_3_i_1 ));
    LocalMux I__2172 (
            .O(N__12717),
            .I(\b2v_inst.reg_ancho_3_i_1 ));
    Odrv12 I__2171 (
            .O(N__12714),
            .I(\b2v_inst.reg_ancho_3_i_1 ));
    CascadeMux I__2170 (
            .O(N__12707),
            .I(N__12704));
    InMux I__2169 (
            .O(N__12704),
            .I(N__12699));
    CascadeMux I__2168 (
            .O(N__12703),
            .I(N__12696));
    CascadeMux I__2167 (
            .O(N__12702),
            .I(N__12693));
    LocalMux I__2166 (
            .O(N__12699),
            .I(N__12690));
    InMux I__2165 (
            .O(N__12696),
            .I(N__12687));
    InMux I__2164 (
            .O(N__12693),
            .I(N__12684));
    Odrv4 I__2163 (
            .O(N__12690),
            .I(\b2v_inst.reg_ancho_3_i_2 ));
    LocalMux I__2162 (
            .O(N__12687),
            .I(\b2v_inst.reg_ancho_3_i_2 ));
    LocalMux I__2161 (
            .O(N__12684),
            .I(\b2v_inst.reg_ancho_3_i_2 ));
    CascadeMux I__2160 (
            .O(N__12677),
            .I(N__12672));
    CascadeMux I__2159 (
            .O(N__12676),
            .I(N__12669));
    CascadeMux I__2158 (
            .O(N__12675),
            .I(N__12666));
    InMux I__2157 (
            .O(N__12672),
            .I(N__12663));
    InMux I__2156 (
            .O(N__12669),
            .I(N__12660));
    InMux I__2155 (
            .O(N__12666),
            .I(N__12657));
    LocalMux I__2154 (
            .O(N__12663),
            .I(N__12654));
    LocalMux I__2153 (
            .O(N__12660),
            .I(\b2v_inst.reg_ancho_3_i_3 ));
    LocalMux I__2152 (
            .O(N__12657),
            .I(\b2v_inst.reg_ancho_3_i_3 ));
    Odrv12 I__2151 (
            .O(N__12654),
            .I(\b2v_inst.reg_ancho_3_i_3 ));
    CascadeMux I__2150 (
            .O(N__12647),
            .I(N__12644));
    InMux I__2149 (
            .O(N__12644),
            .I(N__12639));
    CascadeMux I__2148 (
            .O(N__12643),
            .I(N__12636));
    CascadeMux I__2147 (
            .O(N__12642),
            .I(N__12633));
    LocalMux I__2146 (
            .O(N__12639),
            .I(N__12630));
    InMux I__2145 (
            .O(N__12636),
            .I(N__12627));
    InMux I__2144 (
            .O(N__12633),
            .I(N__12624));
    Odrv4 I__2143 (
            .O(N__12630),
            .I(\b2v_inst.reg_ancho_3_i_4 ));
    LocalMux I__2142 (
            .O(N__12627),
            .I(\b2v_inst.reg_ancho_3_i_4 ));
    LocalMux I__2141 (
            .O(N__12624),
            .I(\b2v_inst.reg_ancho_3_i_4 ));
    CascadeMux I__2140 (
            .O(N__12617),
            .I(N__12614));
    InMux I__2139 (
            .O(N__12614),
            .I(N__12609));
    CascadeMux I__2138 (
            .O(N__12613),
            .I(N__12606));
    CascadeMux I__2137 (
            .O(N__12612),
            .I(N__12603));
    LocalMux I__2136 (
            .O(N__12609),
            .I(N__12600));
    InMux I__2135 (
            .O(N__12606),
            .I(N__12597));
    InMux I__2134 (
            .O(N__12603),
            .I(N__12594));
    Odrv4 I__2133 (
            .O(N__12600),
            .I(\b2v_inst.reg_ancho_3_i_5 ));
    LocalMux I__2132 (
            .O(N__12597),
            .I(\b2v_inst.reg_ancho_3_i_5 ));
    LocalMux I__2131 (
            .O(N__12594),
            .I(\b2v_inst.reg_ancho_3_i_5 ));
    CascadeMux I__2130 (
            .O(N__12587),
            .I(N__12584));
    InMux I__2129 (
            .O(N__12584),
            .I(N__12579));
    CascadeMux I__2128 (
            .O(N__12583),
            .I(N__12576));
    CascadeMux I__2127 (
            .O(N__12582),
            .I(N__12573));
    LocalMux I__2126 (
            .O(N__12579),
            .I(N__12570));
    InMux I__2125 (
            .O(N__12576),
            .I(N__12567));
    InMux I__2124 (
            .O(N__12573),
            .I(N__12564));
    Odrv4 I__2123 (
            .O(N__12570),
            .I(\b2v_inst.reg_ancho_3_i_6 ));
    LocalMux I__2122 (
            .O(N__12567),
            .I(\b2v_inst.reg_ancho_3_i_6 ));
    LocalMux I__2121 (
            .O(N__12564),
            .I(\b2v_inst.reg_ancho_3_i_6 ));
    InMux I__2120 (
            .O(N__12557),
            .I(N__12553));
    InMux I__2119 (
            .O(N__12556),
            .I(N__12550));
    LocalMux I__2118 (
            .O(N__12553),
            .I(SYNTHESIZED_WIRE_10_7));
    LocalMux I__2117 (
            .O(N__12550),
            .I(SYNTHESIZED_WIRE_10_7));
    CascadeMux I__2116 (
            .O(N__12545),
            .I(\b2v_inst.addr_ram_1_iv_i_2_5_cascade_ ));
    CascadeMux I__2115 (
            .O(N__12542),
            .I(N__12538));
    CascadeMux I__2114 (
            .O(N__12541),
            .I(N__12535));
    InMux I__2113 (
            .O(N__12538),
            .I(N__12532));
    InMux I__2112 (
            .O(N__12535),
            .I(N__12529));
    LocalMux I__2111 (
            .O(N__12532),
            .I(N__12526));
    LocalMux I__2110 (
            .O(N__12529),
            .I(N__12523));
    Span4Mux_h I__2109 (
            .O(N__12526),
            .I(N__12520));
    Odrv4 I__2108 (
            .O(N__12523),
            .I(N_54));
    Odrv4 I__2107 (
            .O(N__12520),
            .I(N_54));
    InMux I__2106 (
            .O(N__12515),
            .I(N__12512));
    LocalMux I__2105 (
            .O(N__12512),
            .I(\b2v_inst.addr_ram_1_iv_i_1_5 ));
    InMux I__2104 (
            .O(N__12509),
            .I(N__12506));
    LocalMux I__2103 (
            .O(N__12506),
            .I(\b2v_inst.N_341 ));
    CascadeMux I__2102 (
            .O(N__12503),
            .I(\b2v_inst.N_404_cascade_ ));
    InMux I__2101 (
            .O(N__12500),
            .I(N__12487));
    InMux I__2100 (
            .O(N__12499),
            .I(N__12487));
    InMux I__2099 (
            .O(N__12498),
            .I(N__12474));
    InMux I__2098 (
            .O(N__12497),
            .I(N__12474));
    InMux I__2097 (
            .O(N__12496),
            .I(N__12474));
    InMux I__2096 (
            .O(N__12495),
            .I(N__12474));
    InMux I__2095 (
            .O(N__12494),
            .I(N__12474));
    InMux I__2094 (
            .O(N__12493),
            .I(N__12474));
    InMux I__2093 (
            .O(N__12492),
            .I(N__12470));
    LocalMux I__2092 (
            .O(N__12487),
            .I(N__12467));
    LocalMux I__2091 (
            .O(N__12474),
            .I(N__12464));
    InMux I__2090 (
            .O(N__12473),
            .I(N__12461));
    LocalMux I__2089 (
            .O(N__12470),
            .I(\b2v_inst.cuenta_pixelZ0Z_0 ));
    Odrv12 I__2088 (
            .O(N__12467),
            .I(\b2v_inst.cuenta_pixelZ0Z_0 ));
    Odrv4 I__2087 (
            .O(N__12464),
            .I(\b2v_inst.cuenta_pixelZ0Z_0 ));
    LocalMux I__2086 (
            .O(N__12461),
            .I(\b2v_inst.cuenta_pixelZ0Z_0 ));
    CascadeMux I__2085 (
            .O(N__12452),
            .I(N__12449));
    InMux I__2084 (
            .O(N__12449),
            .I(N__12443));
    InMux I__2083 (
            .O(N__12448),
            .I(N__12443));
    LocalMux I__2082 (
            .O(N__12443),
            .I(N__12440));
    Span4Mux_h I__2081 (
            .O(N__12440),
            .I(N__12434));
    CascadeMux I__2080 (
            .O(N__12439),
            .I(N__12431));
    CascadeMux I__2079 (
            .O(N__12438),
            .I(N__12428));
    CascadeMux I__2078 (
            .O(N__12437),
            .I(N__12423));
    Span4Mux_h I__2077 (
            .O(N__12434),
            .I(N__12418));
    InMux I__2076 (
            .O(N__12431),
            .I(N__12405));
    InMux I__2075 (
            .O(N__12428),
            .I(N__12405));
    InMux I__2074 (
            .O(N__12427),
            .I(N__12405));
    InMux I__2073 (
            .O(N__12426),
            .I(N__12405));
    InMux I__2072 (
            .O(N__12423),
            .I(N__12405));
    InMux I__2071 (
            .O(N__12422),
            .I(N__12405));
    InMux I__2070 (
            .O(N__12421),
            .I(N__12402));
    Odrv4 I__2069 (
            .O(N__12418),
            .I(\b2v_inst.cuenta_pixelZ0Z_1 ));
    LocalMux I__2068 (
            .O(N__12405),
            .I(\b2v_inst.cuenta_pixelZ0Z_1 ));
    LocalMux I__2067 (
            .O(N__12402),
            .I(\b2v_inst.cuenta_pixelZ0Z_1 ));
    InMux I__2066 (
            .O(N__12395),
            .I(N__12392));
    LocalMux I__2065 (
            .O(N__12392),
            .I(N__12389));
    Odrv12 I__2064 (
            .O(N__12389),
            .I(\b2v_inst.cuenta_pixel_4_i_a2_0_6 ));
    InMux I__2063 (
            .O(N__12386),
            .I(N__12383));
    LocalMux I__2062 (
            .O(N__12383),
            .I(N__12380));
    Span4Mux_h I__2061 (
            .O(N__12380),
            .I(N__12377));
    Odrv4 I__2060 (
            .O(N__12377),
            .I(N_213_i));
    InMux I__2059 (
            .O(N__12374),
            .I(N__12371));
    LocalMux I__2058 (
            .O(N__12371),
            .I(N__12368));
    Span4Mux_h I__2057 (
            .O(N__12368),
            .I(N__12365));
    Odrv4 I__2056 (
            .O(N__12365),
            .I(N_209_i));
    InMux I__2055 (
            .O(N__12362),
            .I(N__12359));
    LocalMux I__2054 (
            .O(N__12359),
            .I(N__12356));
    Span4Mux_h I__2053 (
            .O(N__12356),
            .I(N__12353));
    Odrv4 I__2052 (
            .O(N__12353),
            .I(N_207_i));
    InMux I__2051 (
            .O(N__12350),
            .I(N__12346));
    InMux I__2050 (
            .O(N__12349),
            .I(N__12343));
    LocalMux I__2049 (
            .O(N__12346),
            .I(SYNTHESIZED_WIRE_10_2));
    LocalMux I__2048 (
            .O(N__12343),
            .I(SYNTHESIZED_WIRE_10_2));
    InMux I__2047 (
            .O(N__12338),
            .I(N__12334));
    InMux I__2046 (
            .O(N__12337),
            .I(N__12331));
    LocalMux I__2045 (
            .O(N__12334),
            .I(SYNTHESIZED_WIRE_10_3));
    LocalMux I__2044 (
            .O(N__12331),
            .I(SYNTHESIZED_WIRE_10_3));
    InMux I__2043 (
            .O(N__12326),
            .I(N__12322));
    InMux I__2042 (
            .O(N__12325),
            .I(N__12319));
    LocalMux I__2041 (
            .O(N__12322),
            .I(SYNTHESIZED_WIRE_10_4));
    LocalMux I__2040 (
            .O(N__12319),
            .I(SYNTHESIZED_WIRE_10_4));
    InMux I__2039 (
            .O(N__12314),
            .I(N__12310));
    InMux I__2038 (
            .O(N__12313),
            .I(N__12307));
    LocalMux I__2037 (
            .O(N__12310),
            .I(SYNTHESIZED_WIRE_10_5));
    LocalMux I__2036 (
            .O(N__12307),
            .I(SYNTHESIZED_WIRE_10_5));
    CascadeMux I__2035 (
            .O(N__12302),
            .I(N__12298));
    InMux I__2034 (
            .O(N__12301),
            .I(N__12295));
    InMux I__2033 (
            .O(N__12298),
            .I(N__12292));
    LocalMux I__2032 (
            .O(N__12295),
            .I(SYNTHESIZED_WIRE_10_6));
    LocalMux I__2031 (
            .O(N__12292),
            .I(SYNTHESIZED_WIRE_10_6));
    CascadeMux I__2030 (
            .O(N__12287),
            .I(\b2v_inst3.next_bit_0_a3_4_cascade_ ));
    InMux I__2029 (
            .O(N__12284),
            .I(N__12281));
    LocalMux I__2028 (
            .O(N__12281),
            .I(\b2v_inst3.next_bit_0_a3_3 ));
    CascadeMux I__2027 (
            .O(N__12278),
            .I(N__12273));
    InMux I__2026 (
            .O(N__12277),
            .I(N__12266));
    InMux I__2025 (
            .O(N__12276),
            .I(N__12266));
    InMux I__2024 (
            .O(N__12273),
            .I(N__12266));
    LocalMux I__2023 (
            .O(N__12266),
            .I(N__12261));
    InMux I__2022 (
            .O(N__12265),
            .I(N__12258));
    InMux I__2021 (
            .O(N__12264),
            .I(N__12255));
    Span4Mux_v I__2020 (
            .O(N__12261),
            .I(N__12252));
    LocalMux I__2019 (
            .O(N__12258),
            .I(SYNTHESIZED_WIRE_7));
    LocalMux I__2018 (
            .O(N__12255),
            .I(SYNTHESIZED_WIRE_7));
    Odrv4 I__2017 (
            .O(N__12252),
            .I(SYNTHESIZED_WIRE_7));
    CascadeMux I__2016 (
            .O(N__12245),
            .I(\b2v_inst3.N_105_7_cascade_ ));
    InMux I__2015 (
            .O(N__12242),
            .I(N__12238));
    InMux I__2014 (
            .O(N__12241),
            .I(N__12229));
    LocalMux I__2013 (
            .O(N__12238),
            .I(N__12226));
    InMux I__2012 (
            .O(N__12237),
            .I(N__12221));
    InMux I__2011 (
            .O(N__12236),
            .I(N__12221));
    InMux I__2010 (
            .O(N__12235),
            .I(N__12216));
    InMux I__2009 (
            .O(N__12234),
            .I(N__12216));
    InMux I__2008 (
            .O(N__12233),
            .I(N__12211));
    InMux I__2007 (
            .O(N__12232),
            .I(N__12211));
    LocalMux I__2006 (
            .O(N__12229),
            .I(\b2v_inst3.fsm_stateZ0Z_0 ));
    Odrv4 I__2005 (
            .O(N__12226),
            .I(\b2v_inst3.fsm_stateZ0Z_0 ));
    LocalMux I__2004 (
            .O(N__12221),
            .I(\b2v_inst3.fsm_stateZ0Z_0 ));
    LocalMux I__2003 (
            .O(N__12216),
            .I(\b2v_inst3.fsm_stateZ0Z_0 ));
    LocalMux I__2002 (
            .O(N__12211),
            .I(\b2v_inst3.fsm_stateZ0Z_0 ));
    CascadeMux I__2001 (
            .O(N__12200),
            .I(N__12195));
    InMux I__2000 (
            .O(N__12199),
            .I(N__12188));
    InMux I__1999 (
            .O(N__12198),
            .I(N__12188));
    InMux I__1998 (
            .O(N__12195),
            .I(N__12181));
    InMux I__1997 (
            .O(N__12194),
            .I(N__12181));
    InMux I__1996 (
            .O(N__12193),
            .I(N__12181));
    LocalMux I__1995 (
            .O(N__12188),
            .I(\b2v_inst3.cycle_counterZ0Z_1 ));
    LocalMux I__1994 (
            .O(N__12181),
            .I(\b2v_inst3.cycle_counterZ0Z_1 ));
    CascadeMux I__1993 (
            .O(N__12176),
            .I(N__12173));
    InMux I__1992 (
            .O(N__12173),
            .I(N__12167));
    InMux I__1991 (
            .O(N__12172),
            .I(N__12167));
    LocalMux I__1990 (
            .O(N__12167),
            .I(N__12162));
    CascadeMux I__1989 (
            .O(N__12166),
            .I(N__12154));
    InMux I__1988 (
            .O(N__12165),
            .I(N__12150));
    Span4Mux_h I__1987 (
            .O(N__12162),
            .I(N__12147));
    InMux I__1986 (
            .O(N__12161),
            .I(N__12142));
    InMux I__1985 (
            .O(N__12160),
            .I(N__12142));
    InMux I__1984 (
            .O(N__12159),
            .I(N__12135));
    InMux I__1983 (
            .O(N__12158),
            .I(N__12135));
    InMux I__1982 (
            .O(N__12157),
            .I(N__12135));
    InMux I__1981 (
            .O(N__12154),
            .I(N__12130));
    InMux I__1980 (
            .O(N__12153),
            .I(N__12130));
    LocalMux I__1979 (
            .O(N__12150),
            .I(\b2v_inst3.fsm_stateZ0Z_1 ));
    Odrv4 I__1978 (
            .O(N__12147),
            .I(\b2v_inst3.fsm_stateZ0Z_1 ));
    LocalMux I__1977 (
            .O(N__12142),
            .I(\b2v_inst3.fsm_stateZ0Z_1 ));
    LocalMux I__1976 (
            .O(N__12135),
            .I(\b2v_inst3.fsm_stateZ0Z_1 ));
    LocalMux I__1975 (
            .O(N__12130),
            .I(\b2v_inst3.fsm_stateZ0Z_1 ));
    InMux I__1974 (
            .O(N__12119),
            .I(N__12109));
    InMux I__1973 (
            .O(N__12118),
            .I(N__12109));
    InMux I__1972 (
            .O(N__12117),
            .I(N__12100));
    InMux I__1971 (
            .O(N__12116),
            .I(N__12100));
    InMux I__1970 (
            .O(N__12115),
            .I(N__12100));
    InMux I__1969 (
            .O(N__12114),
            .I(N__12100));
    LocalMux I__1968 (
            .O(N__12109),
            .I(\b2v_inst3.cycle_counterZ0Z_0 ));
    LocalMux I__1967 (
            .O(N__12100),
            .I(\b2v_inst3.cycle_counterZ0Z_0 ));
    InMux I__1966 (
            .O(N__12095),
            .I(N__12092));
    LocalMux I__1965 (
            .O(N__12092),
            .I(\b2v_inst3.un1_cycle_counter_5_c2 ));
    CascadeMux I__1964 (
            .O(N__12089),
            .I(N__12085));
    CascadeMux I__1963 (
            .O(N__12088),
            .I(N__12082));
    InMux I__1962 (
            .O(N__12085),
            .I(N__12076));
    InMux I__1961 (
            .O(N__12082),
            .I(N__12071));
    InMux I__1960 (
            .O(N__12081),
            .I(N__12071));
    InMux I__1959 (
            .O(N__12080),
            .I(N__12066));
    InMux I__1958 (
            .O(N__12079),
            .I(N__12066));
    LocalMux I__1957 (
            .O(N__12076),
            .I(\b2v_inst3.cycle_counterZ0Z_2 ));
    LocalMux I__1956 (
            .O(N__12071),
            .I(\b2v_inst3.cycle_counterZ0Z_2 ));
    LocalMux I__1955 (
            .O(N__12066),
            .I(\b2v_inst3.cycle_counterZ0Z_2 ));
    InMux I__1954 (
            .O(N__12059),
            .I(N__12053));
    InMux I__1953 (
            .O(N__12058),
            .I(N__12050));
    InMux I__1952 (
            .O(N__12057),
            .I(N__12045));
    InMux I__1951 (
            .O(N__12056),
            .I(N__12045));
    LocalMux I__1950 (
            .O(N__12053),
            .I(\b2v_inst3.cycle_counterZ0Z_3 ));
    LocalMux I__1949 (
            .O(N__12050),
            .I(\b2v_inst3.cycle_counterZ0Z_3 ));
    LocalMux I__1948 (
            .O(N__12045),
            .I(\b2v_inst3.cycle_counterZ0Z_3 ));
    CascadeMux I__1947 (
            .O(N__12038),
            .I(\b2v_inst3.un1_cycle_counter_5_c2_cascade_ ));
    InMux I__1946 (
            .O(N__12035),
            .I(N__12030));
    InMux I__1945 (
            .O(N__12034),
            .I(N__12025));
    InMux I__1944 (
            .O(N__12033),
            .I(N__12025));
    LocalMux I__1943 (
            .O(N__12030),
            .I(\b2v_inst3.cycle_counterZ0Z_4 ));
    LocalMux I__1942 (
            .O(N__12025),
            .I(\b2v_inst3.cycle_counterZ0Z_4 ));
    InMux I__1941 (
            .O(N__12020),
            .I(N__12017));
    LocalMux I__1940 (
            .O(N__12017),
            .I(N__12014));
    Span4Mux_h I__1939 (
            .O(N__12014),
            .I(N__12004));
    InMux I__1938 (
            .O(N__12013),
            .I(N__11989));
    InMux I__1937 (
            .O(N__12012),
            .I(N__11989));
    InMux I__1936 (
            .O(N__12011),
            .I(N__11989));
    InMux I__1935 (
            .O(N__12010),
            .I(N__11989));
    InMux I__1934 (
            .O(N__12009),
            .I(N__11989));
    InMux I__1933 (
            .O(N__12008),
            .I(N__11989));
    InMux I__1932 (
            .O(N__12007),
            .I(N__11989));
    Odrv4 I__1931 (
            .O(N__12004),
            .I(\b2v_inst4.un1_pix_count_int_0_sqmuxa_9 ));
    LocalMux I__1930 (
            .O(N__11989),
            .I(\b2v_inst4.un1_pix_count_int_0_sqmuxa_9 ));
    InMux I__1929 (
            .O(N__11984),
            .I(N__11981));
    LocalMux I__1928 (
            .O(N__11981),
            .I(N__11978));
    Span4Mux_v I__1927 (
            .O(N__11978),
            .I(N__11968));
    InMux I__1926 (
            .O(N__11977),
            .I(N__11953));
    InMux I__1925 (
            .O(N__11976),
            .I(N__11953));
    InMux I__1924 (
            .O(N__11975),
            .I(N__11953));
    InMux I__1923 (
            .O(N__11974),
            .I(N__11953));
    InMux I__1922 (
            .O(N__11973),
            .I(N__11953));
    InMux I__1921 (
            .O(N__11972),
            .I(N__11953));
    InMux I__1920 (
            .O(N__11971),
            .I(N__11953));
    Odrv4 I__1919 (
            .O(N__11968),
            .I(\b2v_inst4.un1_pix_count_int_0_sqmuxa_11 ));
    LocalMux I__1918 (
            .O(N__11953),
            .I(\b2v_inst4.un1_pix_count_int_0_sqmuxa_11 ));
    CascadeMux I__1917 (
            .O(N__11948),
            .I(N__11941));
    CascadeMux I__1916 (
            .O(N__11947),
            .I(N__11938));
    CascadeMux I__1915 (
            .O(N__11946),
            .I(N__11935));
    CascadeMux I__1914 (
            .O(N__11945),
            .I(N__11932));
    CascadeMux I__1913 (
            .O(N__11944),
            .I(N__11929));
    InMux I__1912 (
            .O(N__11941),
            .I(N__11926));
    InMux I__1911 (
            .O(N__11938),
            .I(N__11914));
    InMux I__1910 (
            .O(N__11935),
            .I(N__11914));
    InMux I__1909 (
            .O(N__11932),
            .I(N__11914));
    InMux I__1908 (
            .O(N__11929),
            .I(N__11914));
    LocalMux I__1907 (
            .O(N__11926),
            .I(N__11911));
    CascadeMux I__1906 (
            .O(N__11925),
            .I(N__11908));
    CascadeMux I__1905 (
            .O(N__11924),
            .I(N__11905));
    CascadeMux I__1904 (
            .O(N__11923),
            .I(N__11902));
    LocalMux I__1903 (
            .O(N__11914),
            .I(N__11897));
    Span4Mux_h I__1902 (
            .O(N__11911),
            .I(N__11897));
    InMux I__1901 (
            .O(N__11908),
            .I(N__11890));
    InMux I__1900 (
            .O(N__11905),
            .I(N__11890));
    InMux I__1899 (
            .O(N__11902),
            .I(N__11890));
    Span4Mux_h I__1898 (
            .O(N__11897),
            .I(N__11887));
    LocalMux I__1897 (
            .O(N__11890),
            .I(\b2v_inst4.un1_pix_count_int_0_sqmuxa_10 ));
    Odrv4 I__1896 (
            .O(N__11887),
            .I(\b2v_inst4.un1_pix_count_int_0_sqmuxa_10 ));
    InMux I__1895 (
            .O(N__11882),
            .I(N__11879));
    LocalMux I__1894 (
            .O(N__11879),
            .I(N__11876));
    Span4Mux_v I__1893 (
            .O(N__11876),
            .I(N__11873));
    Odrv4 I__1892 (
            .O(N__11873),
            .I(\b2v_inst4.pix_count_int_RNO_0Z0Z_9 ));
    InMux I__1891 (
            .O(N__11870),
            .I(N__11864));
    InMux I__1890 (
            .O(N__11869),
            .I(N__11857));
    InMux I__1889 (
            .O(N__11868),
            .I(N__11857));
    InMux I__1888 (
            .O(N__11867),
            .I(N__11857));
    LocalMux I__1887 (
            .O(N__11864),
            .I(N__11852));
    LocalMux I__1886 (
            .O(N__11857),
            .I(N__11852));
    Span4Mux_h I__1885 (
            .O(N__11852),
            .I(N__11849));
    Odrv4 I__1884 (
            .O(N__11849),
            .I(SYNTHESIZED_WIRE_2_9));
    CascadeMux I__1883 (
            .O(N__11846),
            .I(N__11841));
    CascadeMux I__1882 (
            .O(N__11845),
            .I(N__11838));
    InMux I__1881 (
            .O(N__11844),
            .I(N__11835));
    InMux I__1880 (
            .O(N__11841),
            .I(N__11829));
    InMux I__1879 (
            .O(N__11838),
            .I(N__11826));
    LocalMux I__1878 (
            .O(N__11835),
            .I(N__11823));
    InMux I__1877 (
            .O(N__11834),
            .I(N__11816));
    InMux I__1876 (
            .O(N__11833),
            .I(N__11816));
    InMux I__1875 (
            .O(N__11832),
            .I(N__11816));
    LocalMux I__1874 (
            .O(N__11829),
            .I(N__11813));
    LocalMux I__1873 (
            .O(N__11826),
            .I(N__11810));
    Odrv12 I__1872 (
            .O(N__11823),
            .I(\b2v_inst.cuenta_pixelZ0Z_6 ));
    LocalMux I__1871 (
            .O(N__11816),
            .I(\b2v_inst.cuenta_pixelZ0Z_6 ));
    Odrv4 I__1870 (
            .O(N__11813),
            .I(\b2v_inst.cuenta_pixelZ0Z_6 ));
    Odrv4 I__1869 (
            .O(N__11810),
            .I(\b2v_inst.cuenta_pixelZ0Z_6 ));
    CascadeMux I__1868 (
            .O(N__11801),
            .I(N__11798));
    InMux I__1867 (
            .O(N__11798),
            .I(N__11795));
    LocalMux I__1866 (
            .O(N__11795),
            .I(N__11791));
    CascadeMux I__1865 (
            .O(N__11794),
            .I(N__11788));
    Span4Mux_v I__1864 (
            .O(N__11791),
            .I(N__11784));
    InMux I__1863 (
            .O(N__11788),
            .I(N__11779));
    InMux I__1862 (
            .O(N__11787),
            .I(N__11779));
    Span4Mux_h I__1861 (
            .O(N__11784),
            .I(N__11776));
    LocalMux I__1860 (
            .O(N__11779),
            .I(N__11773));
    Odrv4 I__1859 (
            .O(N__11776),
            .I(\b2v_inst.un11_cuenta_pixel_i_0_o2_0 ));
    Odrv12 I__1858 (
            .O(N__11773),
            .I(\b2v_inst.un11_cuenta_pixel_i_0_o2_0 ));
    InMux I__1857 (
            .O(N__11768),
            .I(N__11765));
    LocalMux I__1856 (
            .O(N__11765),
            .I(N__11761));
    CascadeMux I__1855 (
            .O(N__11764),
            .I(N__11756));
    Span4Mux_h I__1854 (
            .O(N__11761),
            .I(N__11752));
    InMux I__1853 (
            .O(N__11760),
            .I(N__11747));
    InMux I__1852 (
            .O(N__11759),
            .I(N__11747));
    InMux I__1851 (
            .O(N__11756),
            .I(N__11742));
    InMux I__1850 (
            .O(N__11755),
            .I(N__11742));
    Odrv4 I__1849 (
            .O(N__11752),
            .I(\b2v_inst.cuenta_pixelZ0Z_5 ));
    LocalMux I__1848 (
            .O(N__11747),
            .I(\b2v_inst.cuenta_pixelZ0Z_5 ));
    LocalMux I__1847 (
            .O(N__11742),
            .I(\b2v_inst.cuenta_pixelZ0Z_5 ));
    IoInMux I__1846 (
            .O(N__11735),
            .I(N__11732));
    LocalMux I__1845 (
            .O(N__11732),
            .I(N__11729));
    Span4Mux_s3_v I__1844 (
            .O(N__11729),
            .I(N__11726));
    Sp12to4 I__1843 (
            .O(N__11726),
            .I(N__11723));
    Span12Mux_h I__1842 (
            .O(N__11723),
            .I(N__11720));
    Span12Mux_v I__1841 (
            .O(N__11720),
            .I(N__11717));
    Odrv12 I__1840 (
            .O(N__11717),
            .I(uart_tx_o));
    InMux I__1839 (
            .O(N__11714),
            .I(N__11710));
    InMux I__1838 (
            .O(N__11713),
            .I(N__11707));
    LocalMux I__1837 (
            .O(N__11710),
            .I(N__11701));
    LocalMux I__1836 (
            .O(N__11707),
            .I(N__11701));
    InMux I__1835 (
            .O(N__11706),
            .I(N__11698));
    Span4Mux_v I__1834 (
            .O(N__11701),
            .I(N__11695));
    LocalMux I__1833 (
            .O(N__11698),
            .I(\b2v_inst4.stateZ0Z_0 ));
    Odrv4 I__1832 (
            .O(N__11695),
            .I(\b2v_inst4.stateZ0Z_0 ));
    InMux I__1831 (
            .O(N__11690),
            .I(N__11683));
    InMux I__1830 (
            .O(N__11689),
            .I(N__11683));
    InMux I__1829 (
            .O(N__11688),
            .I(N__11680));
    LocalMux I__1828 (
            .O(N__11683),
            .I(N__11675));
    LocalMux I__1827 (
            .O(N__11680),
            .I(N__11675));
    Odrv4 I__1826 (
            .O(N__11675),
            .I(\b2v_inst3.cycle_counterZ0Z_6 ));
    InMux I__1825 (
            .O(N__11672),
            .I(N__11662));
    InMux I__1824 (
            .O(N__11671),
            .I(N__11662));
    InMux I__1823 (
            .O(N__11670),
            .I(N__11662));
    InMux I__1822 (
            .O(N__11669),
            .I(N__11659));
    LocalMux I__1821 (
            .O(N__11662),
            .I(\b2v_inst3.cycle_counterZ0Z_5 ));
    LocalMux I__1820 (
            .O(N__11659),
            .I(\b2v_inst3.cycle_counterZ0Z_5 ));
    CascadeMux I__1819 (
            .O(N__11654),
            .I(N__11650));
    InMux I__1818 (
            .O(N__11653),
            .I(N__11647));
    InMux I__1817 (
            .O(N__11650),
            .I(N__11644));
    LocalMux I__1816 (
            .O(N__11647),
            .I(\b2v_inst3.cycle_counterZ0Z_7 ));
    LocalMux I__1815 (
            .O(N__11644),
            .I(\b2v_inst3.cycle_counterZ0Z_7 ));
    InMux I__1814 (
            .O(N__11639),
            .I(bfn_5_20_0_));
    CascadeMux I__1813 (
            .O(N__11636),
            .I(N__11632));
    InMux I__1812 (
            .O(N__11635),
            .I(N__11629));
    InMux I__1811 (
            .O(N__11632),
            .I(N__11626));
    LocalMux I__1810 (
            .O(N__11629),
            .I(N__11623));
    LocalMux I__1809 (
            .O(N__11626),
            .I(N__11620));
    Span4Mux_v I__1808 (
            .O(N__11623),
            .I(N__11617));
    Span4Mux_h I__1807 (
            .O(N__11620),
            .I(N__11614));
    Odrv4 I__1806 (
            .O(N__11617),
            .I(\b2v_inst.valor_max_final52_THRU_CO ));
    Odrv4 I__1805 (
            .O(N__11614),
            .I(\b2v_inst.valor_max_final52_THRU_CO ));
    InMux I__1804 (
            .O(N__11609),
            .I(N__11606));
    LocalMux I__1803 (
            .O(N__11606),
            .I(\b2v_inst3.un1_bit_counter_3_c2 ));
    CascadeMux I__1802 (
            .O(N__11603),
            .I(\b2v_inst3.un1_bit_counter_3_c2_cascade_ ));
    InMux I__1801 (
            .O(N__11600),
            .I(N__11597));
    LocalMux I__1800 (
            .O(N__11597),
            .I(\b2v_inst3.N_258 ));
    CascadeMux I__1799 (
            .O(N__11594),
            .I(\b2v_inst3.N_258_cascade_ ));
    InMux I__1798 (
            .O(N__11591),
            .I(N__11583));
    InMux I__1797 (
            .O(N__11590),
            .I(N__11583));
    InMux I__1796 (
            .O(N__11589),
            .I(N__11578));
    InMux I__1795 (
            .O(N__11588),
            .I(N__11578));
    LocalMux I__1794 (
            .O(N__11583),
            .I(\b2v_inst3.bit_counterZ0Z_2 ));
    LocalMux I__1793 (
            .O(N__11578),
            .I(\b2v_inst3.bit_counterZ0Z_2 ));
    InMux I__1792 (
            .O(N__11573),
            .I(N__11565));
    InMux I__1791 (
            .O(N__11572),
            .I(N__11565));
    InMux I__1790 (
            .O(N__11571),
            .I(N__11560));
    InMux I__1789 (
            .O(N__11570),
            .I(N__11560));
    LocalMux I__1788 (
            .O(N__11565),
            .I(\b2v_inst3.bit_counterZ1Z_1 ));
    LocalMux I__1787 (
            .O(N__11560),
            .I(\b2v_inst3.bit_counterZ1Z_1 ));
    CascadeMux I__1786 (
            .O(N__11555),
            .I(\b2v_inst3.N_102_2_cascade_ ));
    CascadeMux I__1785 (
            .O(N__11552),
            .I(N__11547));
    InMux I__1784 (
            .O(N__11551),
            .I(N__11540));
    InMux I__1783 (
            .O(N__11550),
            .I(N__11540));
    InMux I__1782 (
            .O(N__11547),
            .I(N__11540));
    LocalMux I__1781 (
            .O(N__11540),
            .I(\b2v_inst3.bit_counterZ0Z_3 ));
    InMux I__1780 (
            .O(N__11537),
            .I(N__11533));
    InMux I__1779 (
            .O(N__11536),
            .I(N__11530));
    LocalMux I__1778 (
            .O(N__11533),
            .I(\b2v_inst3.N_436 ));
    LocalMux I__1777 (
            .O(N__11530),
            .I(\b2v_inst3.N_436 ));
    InMux I__1776 (
            .O(N__11525),
            .I(N__11522));
    LocalMux I__1775 (
            .O(N__11522),
            .I(N__11519));
    Span4Mux_h I__1774 (
            .O(N__11519),
            .I(N__11516));
    Odrv4 I__1773 (
            .O(N__11516),
            .I(\b2v_inst.data_a_escribir9_6_and ));
    CascadeMux I__1772 (
            .O(N__11513),
            .I(N__11507));
    InMux I__1771 (
            .O(N__11512),
            .I(N__11503));
    InMux I__1770 (
            .O(N__11511),
            .I(N__11500));
    InMux I__1769 (
            .O(N__11510),
            .I(N__11497));
    InMux I__1768 (
            .O(N__11507),
            .I(N__11494));
    InMux I__1767 (
            .O(N__11506),
            .I(N__11491));
    LocalMux I__1766 (
            .O(N__11503),
            .I(N__11488));
    LocalMux I__1765 (
            .O(N__11500),
            .I(N__11485));
    LocalMux I__1764 (
            .O(N__11497),
            .I(\b2v_inst.reg_ancho_2Z0Z_0 ));
    LocalMux I__1763 (
            .O(N__11494),
            .I(\b2v_inst.reg_ancho_2Z0Z_0 ));
    LocalMux I__1762 (
            .O(N__11491),
            .I(\b2v_inst.reg_ancho_2Z0Z_0 ));
    Odrv4 I__1761 (
            .O(N__11488),
            .I(\b2v_inst.reg_ancho_2Z0Z_0 ));
    Odrv4 I__1760 (
            .O(N__11485),
            .I(\b2v_inst.reg_ancho_2Z0Z_0 ));
    InMux I__1759 (
            .O(N__11474),
            .I(N__11468));
    InMux I__1758 (
            .O(N__11473),
            .I(N__11465));
    InMux I__1757 (
            .O(N__11472),
            .I(N__11462));
    CascadeMux I__1756 (
            .O(N__11471),
            .I(N__11459));
    LocalMux I__1755 (
            .O(N__11468),
            .I(N__11455));
    LocalMux I__1754 (
            .O(N__11465),
            .I(N__11452));
    LocalMux I__1753 (
            .O(N__11462),
            .I(N__11449));
    InMux I__1752 (
            .O(N__11459),
            .I(N__11446));
    InMux I__1751 (
            .O(N__11458),
            .I(N__11443));
    Span4Mux_h I__1750 (
            .O(N__11455),
            .I(N__11438));
    Span4Mux_v I__1749 (
            .O(N__11452),
            .I(N__11438));
    Odrv4 I__1748 (
            .O(N__11449),
            .I(\b2v_inst.reg_ancho_2Z0Z_1 ));
    LocalMux I__1747 (
            .O(N__11446),
            .I(\b2v_inst.reg_ancho_2Z0Z_1 ));
    LocalMux I__1746 (
            .O(N__11443),
            .I(\b2v_inst.reg_ancho_2Z0Z_1 ));
    Odrv4 I__1745 (
            .O(N__11438),
            .I(\b2v_inst.reg_ancho_2Z0Z_1 ));
    CascadeMux I__1744 (
            .O(N__11429),
            .I(N__11423));
    InMux I__1743 (
            .O(N__11428),
            .I(N__11420));
    InMux I__1742 (
            .O(N__11427),
            .I(N__11416));
    InMux I__1741 (
            .O(N__11426),
            .I(N__11413));
    InMux I__1740 (
            .O(N__11423),
            .I(N__11410));
    LocalMux I__1739 (
            .O(N__11420),
            .I(N__11407));
    InMux I__1738 (
            .O(N__11419),
            .I(N__11404));
    LocalMux I__1737 (
            .O(N__11416),
            .I(N__11401));
    LocalMux I__1736 (
            .O(N__11413),
            .I(\b2v_inst.reg_ancho_2Z0Z_2 ));
    LocalMux I__1735 (
            .O(N__11410),
            .I(\b2v_inst.reg_ancho_2Z0Z_2 ));
    Odrv4 I__1734 (
            .O(N__11407),
            .I(\b2v_inst.reg_ancho_2Z0Z_2 ));
    LocalMux I__1733 (
            .O(N__11404),
            .I(\b2v_inst.reg_ancho_2Z0Z_2 ));
    Odrv4 I__1732 (
            .O(N__11401),
            .I(\b2v_inst.reg_ancho_2Z0Z_2 ));
    CascadeMux I__1731 (
            .O(N__11390),
            .I(N__11383));
    CascadeMux I__1730 (
            .O(N__11389),
            .I(N__11380));
    InMux I__1729 (
            .O(N__11388),
            .I(N__11377));
    CascadeMux I__1728 (
            .O(N__11387),
            .I(N__11374));
    InMux I__1727 (
            .O(N__11386),
            .I(N__11371));
    InMux I__1726 (
            .O(N__11383),
            .I(N__11368));
    InMux I__1725 (
            .O(N__11380),
            .I(N__11365));
    LocalMux I__1724 (
            .O(N__11377),
            .I(N__11362));
    InMux I__1723 (
            .O(N__11374),
            .I(N__11359));
    LocalMux I__1722 (
            .O(N__11371),
            .I(N__11356));
    LocalMux I__1721 (
            .O(N__11368),
            .I(\b2v_inst.reg_ancho_2Z0Z_3 ));
    LocalMux I__1720 (
            .O(N__11365),
            .I(\b2v_inst.reg_ancho_2Z0Z_3 ));
    Odrv4 I__1719 (
            .O(N__11362),
            .I(\b2v_inst.reg_ancho_2Z0Z_3 ));
    LocalMux I__1718 (
            .O(N__11359),
            .I(\b2v_inst.reg_ancho_2Z0Z_3 ));
    Odrv4 I__1717 (
            .O(N__11356),
            .I(\b2v_inst.reg_ancho_2Z0Z_3 ));
    InMux I__1716 (
            .O(N__11345),
            .I(N__11341));
    InMux I__1715 (
            .O(N__11344),
            .I(N__11338));
    LocalMux I__1714 (
            .O(N__11341),
            .I(N__11334));
    LocalMux I__1713 (
            .O(N__11338),
            .I(N__11331));
    InMux I__1712 (
            .O(N__11337),
            .I(N__11328));
    Span4Mux_v I__1711 (
            .O(N__11334),
            .I(N__11319));
    Span4Mux_v I__1710 (
            .O(N__11331),
            .I(N__11319));
    LocalMux I__1709 (
            .O(N__11328),
            .I(N__11319));
    InMux I__1708 (
            .O(N__11327),
            .I(N__11314));
    InMux I__1707 (
            .O(N__11326),
            .I(N__11314));
    Odrv4 I__1706 (
            .O(N__11319),
            .I(\b2v_inst.reg_ancho_2Z0Z_4 ));
    LocalMux I__1705 (
            .O(N__11314),
            .I(\b2v_inst.reg_ancho_2Z0Z_4 ));
    InMux I__1704 (
            .O(N__11309),
            .I(N__11305));
    InMux I__1703 (
            .O(N__11308),
            .I(N__11300));
    LocalMux I__1702 (
            .O(N__11305),
            .I(N__11297));
    InMux I__1701 (
            .O(N__11304),
            .I(N__11294));
    InMux I__1700 (
            .O(N__11303),
            .I(N__11290));
    LocalMux I__1699 (
            .O(N__11300),
            .I(N__11287));
    Span4Mux_v I__1698 (
            .O(N__11297),
            .I(N__11284));
    LocalMux I__1697 (
            .O(N__11294),
            .I(N__11281));
    InMux I__1696 (
            .O(N__11293),
            .I(N__11278));
    LocalMux I__1695 (
            .O(N__11290),
            .I(\b2v_inst.reg_ancho_2Z0Z_5 ));
    Odrv4 I__1694 (
            .O(N__11287),
            .I(\b2v_inst.reg_ancho_2Z0Z_5 ));
    Odrv4 I__1693 (
            .O(N__11284),
            .I(\b2v_inst.reg_ancho_2Z0Z_5 ));
    Odrv12 I__1692 (
            .O(N__11281),
            .I(\b2v_inst.reg_ancho_2Z0Z_5 ));
    LocalMux I__1691 (
            .O(N__11278),
            .I(\b2v_inst.reg_ancho_2Z0Z_5 ));
    CascadeMux I__1690 (
            .O(N__11267),
            .I(N__11264));
    InMux I__1689 (
            .O(N__11264),
            .I(N__11259));
    InMux I__1688 (
            .O(N__11263),
            .I(N__11256));
    InMux I__1687 (
            .O(N__11262),
            .I(N__11253));
    LocalMux I__1686 (
            .O(N__11259),
            .I(N__11250));
    LocalMux I__1685 (
            .O(N__11256),
            .I(N__11247));
    LocalMux I__1684 (
            .O(N__11253),
            .I(N__11244));
    Span4Mux_v I__1683 (
            .O(N__11250),
            .I(N__11235));
    Span4Mux_v I__1682 (
            .O(N__11247),
            .I(N__11235));
    Span4Mux_v I__1681 (
            .O(N__11244),
            .I(N__11235));
    InMux I__1680 (
            .O(N__11243),
            .I(N__11232));
    InMux I__1679 (
            .O(N__11242),
            .I(N__11229));
    Odrv4 I__1678 (
            .O(N__11235),
            .I(\b2v_inst.reg_ancho_2Z0Z_6 ));
    LocalMux I__1677 (
            .O(N__11232),
            .I(\b2v_inst.reg_ancho_2Z0Z_6 ));
    LocalMux I__1676 (
            .O(N__11229),
            .I(\b2v_inst.reg_ancho_2Z0Z_6 ));
    CascadeMux I__1675 (
            .O(N__11222),
            .I(N__11218));
    InMux I__1674 (
            .O(N__11221),
            .I(N__11214));
    InMux I__1673 (
            .O(N__11218),
            .I(N__11210));
    CascadeMux I__1672 (
            .O(N__11217),
            .I(N__11207));
    LocalMux I__1671 (
            .O(N__11214),
            .I(N__11204));
    InMux I__1670 (
            .O(N__11213),
            .I(N__11200));
    LocalMux I__1669 (
            .O(N__11210),
            .I(N__11197));
    InMux I__1668 (
            .O(N__11207),
            .I(N__11194));
    Span4Mux_v I__1667 (
            .O(N__11204),
            .I(N__11191));
    CascadeMux I__1666 (
            .O(N__11203),
            .I(N__11188));
    LocalMux I__1665 (
            .O(N__11200),
            .I(N__11185));
    Span4Mux_h I__1664 (
            .O(N__11197),
            .I(N__11178));
    LocalMux I__1663 (
            .O(N__11194),
            .I(N__11178));
    Span4Mux_h I__1662 (
            .O(N__11191),
            .I(N__11178));
    InMux I__1661 (
            .O(N__11188),
            .I(N__11175));
    Odrv4 I__1660 (
            .O(N__11185),
            .I(\b2v_inst.reg_ancho_2Z0Z_7 ));
    Odrv4 I__1659 (
            .O(N__11178),
            .I(\b2v_inst.reg_ancho_2Z0Z_7 ));
    LocalMux I__1658 (
            .O(N__11175),
            .I(\b2v_inst.reg_ancho_2Z0Z_7 ));
    InMux I__1657 (
            .O(N__11168),
            .I(N__11164));
    InMux I__1656 (
            .O(N__11167),
            .I(N__11160));
    LocalMux I__1655 (
            .O(N__11164),
            .I(N__11157));
    InMux I__1654 (
            .O(N__11163),
            .I(N__11152));
    LocalMux I__1653 (
            .O(N__11160),
            .I(N__11149));
    Span4Mux_h I__1652 (
            .O(N__11157),
            .I(N__11146));
    InMux I__1651 (
            .O(N__11156),
            .I(N__11143));
    InMux I__1650 (
            .O(N__11155),
            .I(N__11140));
    LocalMux I__1649 (
            .O(N__11152),
            .I(\b2v_inst.reg_ancho_1Z0Z_1 ));
    Odrv4 I__1648 (
            .O(N__11149),
            .I(\b2v_inst.reg_ancho_1Z0Z_1 ));
    Odrv4 I__1647 (
            .O(N__11146),
            .I(\b2v_inst.reg_ancho_1Z0Z_1 ));
    LocalMux I__1646 (
            .O(N__11143),
            .I(\b2v_inst.reg_ancho_1Z0Z_1 ));
    LocalMux I__1645 (
            .O(N__11140),
            .I(\b2v_inst.reg_ancho_1Z0Z_1 ));
    InMux I__1644 (
            .O(N__11129),
            .I(N__11126));
    LocalMux I__1643 (
            .O(N__11126),
            .I(N__11122));
    InMux I__1642 (
            .O(N__11125),
            .I(N__11118));
    Span4Mux_v I__1641 (
            .O(N__11122),
            .I(N__11115));
    InMux I__1640 (
            .O(N__11121),
            .I(N__11112));
    LocalMux I__1639 (
            .O(N__11118),
            .I(N__11109));
    Odrv4 I__1638 (
            .O(N__11115),
            .I(\b2v_inst.reg_ancho_3Z0Z_1 ));
    LocalMux I__1637 (
            .O(N__11112),
            .I(\b2v_inst.reg_ancho_3Z0Z_1 ));
    Odrv4 I__1636 (
            .O(N__11109),
            .I(\b2v_inst.reg_ancho_3Z0Z_1 ));
    InMux I__1635 (
            .O(N__11102),
            .I(N__11099));
    LocalMux I__1634 (
            .O(N__11099),
            .I(N__11095));
    InMux I__1633 (
            .O(N__11098),
            .I(N__11091));
    Span4Mux_h I__1632 (
            .O(N__11095),
            .I(N__11088));
    InMux I__1631 (
            .O(N__11094),
            .I(N__11085));
    LocalMux I__1630 (
            .O(N__11091),
            .I(N__11082));
    Odrv4 I__1629 (
            .O(N__11088),
            .I(\b2v_inst.reg_ancho_3Z0Z_2 ));
    LocalMux I__1628 (
            .O(N__11085),
            .I(\b2v_inst.reg_ancho_3Z0Z_2 ));
    Odrv12 I__1627 (
            .O(N__11082),
            .I(\b2v_inst.reg_ancho_3Z0Z_2 ));
    CascadeMux I__1626 (
            .O(N__11075),
            .I(N__11071));
    InMux I__1625 (
            .O(N__11074),
            .I(N__11067));
    InMux I__1624 (
            .O(N__11071),
            .I(N__11064));
    InMux I__1623 (
            .O(N__11070),
            .I(N__11061));
    LocalMux I__1622 (
            .O(N__11067),
            .I(N__11057));
    LocalMux I__1621 (
            .O(N__11064),
            .I(N__11051));
    LocalMux I__1620 (
            .O(N__11061),
            .I(N__11051));
    InMux I__1619 (
            .O(N__11060),
            .I(N__11048));
    Span4Mux_h I__1618 (
            .O(N__11057),
            .I(N__11045));
    InMux I__1617 (
            .O(N__11056),
            .I(N__11042));
    Odrv4 I__1616 (
            .O(N__11051),
            .I(\b2v_inst.reg_ancho_1Z0Z_2 ));
    LocalMux I__1615 (
            .O(N__11048),
            .I(\b2v_inst.reg_ancho_1Z0Z_2 ));
    Odrv4 I__1614 (
            .O(N__11045),
            .I(\b2v_inst.reg_ancho_1Z0Z_2 ));
    LocalMux I__1613 (
            .O(N__11042),
            .I(\b2v_inst.reg_ancho_1Z0Z_2 ));
    InMux I__1612 (
            .O(N__11033),
            .I(N__11029));
    InMux I__1611 (
            .O(N__11032),
            .I(N__11026));
    LocalMux I__1610 (
            .O(N__11029),
            .I(N__11023));
    LocalMux I__1609 (
            .O(N__11026),
            .I(N__11018));
    Span4Mux_v I__1608 (
            .O(N__11023),
            .I(N__11015));
    CascadeMux I__1607 (
            .O(N__11022),
            .I(N__11012));
    InMux I__1606 (
            .O(N__11021),
            .I(N__11008));
    Span4Mux_h I__1605 (
            .O(N__11018),
            .I(N__11003));
    Span4Mux_h I__1604 (
            .O(N__11015),
            .I(N__11003));
    InMux I__1603 (
            .O(N__11012),
            .I(N__11000));
    InMux I__1602 (
            .O(N__11011),
            .I(N__10997));
    LocalMux I__1601 (
            .O(N__11008),
            .I(\b2v_inst.reg_ancho_1Z0Z_3 ));
    Odrv4 I__1600 (
            .O(N__11003),
            .I(\b2v_inst.reg_ancho_1Z0Z_3 ));
    LocalMux I__1599 (
            .O(N__11000),
            .I(\b2v_inst.reg_ancho_1Z0Z_3 ));
    LocalMux I__1598 (
            .O(N__10997),
            .I(\b2v_inst.reg_ancho_1Z0Z_3 ));
    InMux I__1597 (
            .O(N__10988),
            .I(N__10985));
    LocalMux I__1596 (
            .O(N__10985),
            .I(N__10981));
    CascadeMux I__1595 (
            .O(N__10984),
            .I(N__10977));
    Span4Mux_v I__1594 (
            .O(N__10981),
            .I(N__10974));
    InMux I__1593 (
            .O(N__10980),
            .I(N__10971));
    InMux I__1592 (
            .O(N__10977),
            .I(N__10968));
    Span4Mux_h I__1591 (
            .O(N__10974),
            .I(N__10963));
    LocalMux I__1590 (
            .O(N__10971),
            .I(N__10963));
    LocalMux I__1589 (
            .O(N__10968),
            .I(\b2v_inst.reg_ancho_3Z0Z_3 ));
    Odrv4 I__1588 (
            .O(N__10963),
            .I(\b2v_inst.reg_ancho_3Z0Z_3 ));
    InMux I__1587 (
            .O(N__10958),
            .I(N__10955));
    LocalMux I__1586 (
            .O(N__10955),
            .I(N__10951));
    InMux I__1585 (
            .O(N__10954),
            .I(N__10947));
    Span4Mux_v I__1584 (
            .O(N__10951),
            .I(N__10943));
    InMux I__1583 (
            .O(N__10950),
            .I(N__10939));
    LocalMux I__1582 (
            .O(N__10947),
            .I(N__10936));
    InMux I__1581 (
            .O(N__10946),
            .I(N__10933));
    Span4Mux_h I__1580 (
            .O(N__10943),
            .I(N__10930));
    InMux I__1579 (
            .O(N__10942),
            .I(N__10927));
    LocalMux I__1578 (
            .O(N__10939),
            .I(\b2v_inst.reg_ancho_1Z0Z_4 ));
    Odrv4 I__1577 (
            .O(N__10936),
            .I(\b2v_inst.reg_ancho_1Z0Z_4 ));
    LocalMux I__1576 (
            .O(N__10933),
            .I(\b2v_inst.reg_ancho_1Z0Z_4 ));
    Odrv4 I__1575 (
            .O(N__10930),
            .I(\b2v_inst.reg_ancho_1Z0Z_4 ));
    LocalMux I__1574 (
            .O(N__10927),
            .I(\b2v_inst.reg_ancho_1Z0Z_4 ));
    InMux I__1573 (
            .O(N__10916),
            .I(N__10913));
    LocalMux I__1572 (
            .O(N__10913),
            .I(N__10910));
    Span4Mux_h I__1571 (
            .O(N__10910),
            .I(N__10906));
    InMux I__1570 (
            .O(N__10909),
            .I(N__10902));
    Span4Mux_v I__1569 (
            .O(N__10906),
            .I(N__10899));
    InMux I__1568 (
            .O(N__10905),
            .I(N__10896));
    LocalMux I__1567 (
            .O(N__10902),
            .I(N__10893));
    Odrv4 I__1566 (
            .O(N__10899),
            .I(\b2v_inst.reg_ancho_3Z0Z_4 ));
    LocalMux I__1565 (
            .O(N__10896),
            .I(\b2v_inst.reg_ancho_3Z0Z_4 ));
    Odrv4 I__1564 (
            .O(N__10893),
            .I(\b2v_inst.reg_ancho_3Z0Z_4 ));
    InMux I__1563 (
            .O(N__10886),
            .I(N__10881));
    InMux I__1562 (
            .O(N__10885),
            .I(N__10878));
    InMux I__1561 (
            .O(N__10884),
            .I(N__10875));
    LocalMux I__1560 (
            .O(N__10881),
            .I(N__10872));
    LocalMux I__1559 (
            .O(N__10878),
            .I(N__10865));
    LocalMux I__1558 (
            .O(N__10875),
            .I(N__10865));
    Span4Mux_h I__1557 (
            .O(N__10872),
            .I(N__10862));
    InMux I__1556 (
            .O(N__10871),
            .I(N__10859));
    InMux I__1555 (
            .O(N__10870),
            .I(N__10856));
    Odrv4 I__1554 (
            .O(N__10865),
            .I(\b2v_inst.reg_ancho_1Z0Z_5 ));
    Odrv4 I__1553 (
            .O(N__10862),
            .I(\b2v_inst.reg_ancho_1Z0Z_5 ));
    LocalMux I__1552 (
            .O(N__10859),
            .I(\b2v_inst.reg_ancho_1Z0Z_5 ));
    LocalMux I__1551 (
            .O(N__10856),
            .I(\b2v_inst.reg_ancho_1Z0Z_5 ));
    InMux I__1550 (
            .O(N__10847),
            .I(N__10842));
    InMux I__1549 (
            .O(N__10846),
            .I(N__10839));
    InMux I__1548 (
            .O(N__10845),
            .I(N__10836));
    LocalMux I__1547 (
            .O(N__10842),
            .I(N__10833));
    LocalMux I__1546 (
            .O(N__10839),
            .I(N__10830));
    LocalMux I__1545 (
            .O(N__10836),
            .I(N__10825));
    Span4Mux_h I__1544 (
            .O(N__10833),
            .I(N__10822));
    Span4Mux_h I__1543 (
            .O(N__10830),
            .I(N__10819));
    InMux I__1542 (
            .O(N__10829),
            .I(N__10816));
    InMux I__1541 (
            .O(N__10828),
            .I(N__10813));
    Odrv12 I__1540 (
            .O(N__10825),
            .I(\b2v_inst.reg_ancho_1Z0Z_6 ));
    Odrv4 I__1539 (
            .O(N__10822),
            .I(\b2v_inst.reg_ancho_1Z0Z_6 ));
    Odrv4 I__1538 (
            .O(N__10819),
            .I(\b2v_inst.reg_ancho_1Z0Z_6 ));
    LocalMux I__1537 (
            .O(N__10816),
            .I(\b2v_inst.reg_ancho_1Z0Z_6 ));
    LocalMux I__1536 (
            .O(N__10813),
            .I(\b2v_inst.reg_ancho_1Z0Z_6 ));
    InMux I__1535 (
            .O(N__10802),
            .I(N__10798));
    InMux I__1534 (
            .O(N__10801),
            .I(N__10795));
    LocalMux I__1533 (
            .O(N__10798),
            .I(N__10790));
    LocalMux I__1532 (
            .O(N__10795),
            .I(N__10787));
    CascadeMux I__1531 (
            .O(N__10794),
            .I(N__10784));
    InMux I__1530 (
            .O(N__10793),
            .I(N__10780));
    Span4Mux_v I__1529 (
            .O(N__10790),
            .I(N__10777));
    Span4Mux_h I__1528 (
            .O(N__10787),
            .I(N__10774));
    InMux I__1527 (
            .O(N__10784),
            .I(N__10771));
    InMux I__1526 (
            .O(N__10783),
            .I(N__10768));
    LocalMux I__1525 (
            .O(N__10780),
            .I(\b2v_inst.reg_ancho_1Z0Z_7 ));
    Odrv4 I__1524 (
            .O(N__10777),
            .I(\b2v_inst.reg_ancho_1Z0Z_7 ));
    Odrv4 I__1523 (
            .O(N__10774),
            .I(\b2v_inst.reg_ancho_1Z0Z_7 ));
    LocalMux I__1522 (
            .O(N__10771),
            .I(\b2v_inst.reg_ancho_1Z0Z_7 ));
    LocalMux I__1521 (
            .O(N__10768),
            .I(\b2v_inst.reg_ancho_1Z0Z_7 ));
    CascadeMux I__1520 (
            .O(N__10757),
            .I(N__10753));
    CascadeMux I__1519 (
            .O(N__10756),
            .I(N__10749));
    InMux I__1518 (
            .O(N__10753),
            .I(N__10746));
    InMux I__1517 (
            .O(N__10752),
            .I(N__10743));
    InMux I__1516 (
            .O(N__10749),
            .I(N__10740));
    LocalMux I__1515 (
            .O(N__10746),
            .I(N__10735));
    LocalMux I__1514 (
            .O(N__10743),
            .I(N__10735));
    LocalMux I__1513 (
            .O(N__10740),
            .I(\b2v_inst.reg_ancho_3Z0Z_7 ));
    Odrv4 I__1512 (
            .O(N__10735),
            .I(\b2v_inst.reg_ancho_3Z0Z_7 ));
    InMux I__1511 (
            .O(N__10730),
            .I(bfn_5_18_0_));
    InMux I__1510 (
            .O(N__10727),
            .I(N__10724));
    LocalMux I__1509 (
            .O(N__10724),
            .I(N__10721));
    Span4Mux_h I__1508 (
            .O(N__10721),
            .I(N__10718));
    Odrv4 I__1507 (
            .O(N__10718),
            .I(\b2v_inst.valor_max_final50_THRU_CO ));
    InMux I__1506 (
            .O(N__10715),
            .I(N__10712));
    LocalMux I__1505 (
            .O(N__10712),
            .I(N__10709));
    Odrv4 I__1504 (
            .O(N__10709),
            .I(\b2v_inst.data_a_escribir9_5_and ));
    InMux I__1503 (
            .O(N__10706),
            .I(N__10702));
    InMux I__1502 (
            .O(N__10705),
            .I(N__10697));
    LocalMux I__1501 (
            .O(N__10702),
            .I(N__10692));
    InMux I__1500 (
            .O(N__10701),
            .I(N__10689));
    InMux I__1499 (
            .O(N__10700),
            .I(N__10685));
    LocalMux I__1498 (
            .O(N__10697),
            .I(N__10682));
    InMux I__1497 (
            .O(N__10696),
            .I(N__10673));
    InMux I__1496 (
            .O(N__10695),
            .I(N__10673));
    Span4Mux_v I__1495 (
            .O(N__10692),
            .I(N__10668));
    LocalMux I__1494 (
            .O(N__10689),
            .I(N__10668));
    InMux I__1493 (
            .O(N__10688),
            .I(N__10665));
    LocalMux I__1492 (
            .O(N__10685),
            .I(N__10662));
    Span4Mux_v I__1491 (
            .O(N__10682),
            .I(N__10659));
    InMux I__1490 (
            .O(N__10681),
            .I(N__10654));
    InMux I__1489 (
            .O(N__10680),
            .I(N__10654));
    InMux I__1488 (
            .O(N__10679),
            .I(N__10649));
    InMux I__1487 (
            .O(N__10678),
            .I(N__10649));
    LocalMux I__1486 (
            .O(N__10673),
            .I(N__10646));
    Span4Mux_h I__1485 (
            .O(N__10668),
            .I(N__10641));
    LocalMux I__1484 (
            .O(N__10665),
            .I(N__10641));
    Odrv4 I__1483 (
            .O(N__10662),
            .I(\b2v_inst.un3_valor_max1_THRU_CO ));
    Odrv4 I__1482 (
            .O(N__10659),
            .I(\b2v_inst.un3_valor_max1_THRU_CO ));
    LocalMux I__1481 (
            .O(N__10654),
            .I(\b2v_inst.un3_valor_max1_THRU_CO ));
    LocalMux I__1480 (
            .O(N__10649),
            .I(\b2v_inst.un3_valor_max1_THRU_CO ));
    Odrv4 I__1479 (
            .O(N__10646),
            .I(\b2v_inst.un3_valor_max1_THRU_CO ));
    Odrv4 I__1478 (
            .O(N__10641),
            .I(\b2v_inst.un3_valor_max1_THRU_CO ));
    InMux I__1477 (
            .O(N__10628),
            .I(N__10625));
    LocalMux I__1476 (
            .O(N__10625),
            .I(N__10622));
    Odrv4 I__1475 (
            .O(N__10622),
            .I(\b2v_inst.data_a_escribir_RNO_3Z0Z_6 ));
    InMux I__1474 (
            .O(N__10619),
            .I(N__10616));
    LocalMux I__1473 (
            .O(N__10616),
            .I(N__10613));
    Span4Mux_h I__1472 (
            .O(N__10613),
            .I(N__10607));
    InMux I__1471 (
            .O(N__10612),
            .I(N__10604));
    InMux I__1470 (
            .O(N__10611),
            .I(N__10601));
    InMux I__1469 (
            .O(N__10610),
            .I(N__10598));
    Odrv4 I__1468 (
            .O(N__10607),
            .I(\b2v_inst.un1_reg_anterior_iv_0_0_a2_6_0_1 ));
    LocalMux I__1467 (
            .O(N__10604),
            .I(\b2v_inst.un1_reg_anterior_iv_0_0_a2_6_0_1 ));
    LocalMux I__1466 (
            .O(N__10601),
            .I(\b2v_inst.un1_reg_anterior_iv_0_0_a2_6_0_1 ));
    LocalMux I__1465 (
            .O(N__10598),
            .I(\b2v_inst.un1_reg_anterior_iv_0_0_a2_6_0_1 ));
    InMux I__1464 (
            .O(N__10589),
            .I(N__10586));
    LocalMux I__1463 (
            .O(N__10586),
            .I(\b2v_inst.un1_m3_0_0 ));
    InMux I__1462 (
            .O(N__10583),
            .I(N__10580));
    LocalMux I__1461 (
            .O(N__10580),
            .I(N__10577));
    Odrv4 I__1460 (
            .O(N__10577),
            .I(\b2v_inst.un1_reg_anterior_iv_0_0_0_6 ));
    CascadeMux I__1459 (
            .O(N__10574),
            .I(\b2v_inst.data_a_escribir_RNO_1Z0Z_6_cascade_ ));
    CascadeMux I__1458 (
            .O(N__10571),
            .I(N__10564));
    CascadeMux I__1457 (
            .O(N__10570),
            .I(N__10559));
    CascadeMux I__1456 (
            .O(N__10569),
            .I(N__10554));
    InMux I__1455 (
            .O(N__10568),
            .I(N__10548));
    InMux I__1454 (
            .O(N__10567),
            .I(N__10548));
    InMux I__1453 (
            .O(N__10564),
            .I(N__10537));
    InMux I__1452 (
            .O(N__10563),
            .I(N__10534));
    InMux I__1451 (
            .O(N__10562),
            .I(N__10531));
    InMux I__1450 (
            .O(N__10559),
            .I(N__10528));
    InMux I__1449 (
            .O(N__10558),
            .I(N__10519));
    InMux I__1448 (
            .O(N__10557),
            .I(N__10519));
    InMux I__1447 (
            .O(N__10554),
            .I(N__10519));
    InMux I__1446 (
            .O(N__10553),
            .I(N__10519));
    LocalMux I__1445 (
            .O(N__10548),
            .I(N__10507));
    InMux I__1444 (
            .O(N__10547),
            .I(N__10494));
    InMux I__1443 (
            .O(N__10546),
            .I(N__10494));
    InMux I__1442 (
            .O(N__10545),
            .I(N__10494));
    InMux I__1441 (
            .O(N__10544),
            .I(N__10494));
    InMux I__1440 (
            .O(N__10543),
            .I(N__10494));
    InMux I__1439 (
            .O(N__10542),
            .I(N__10494));
    InMux I__1438 (
            .O(N__10541),
            .I(N__10489));
    InMux I__1437 (
            .O(N__10540),
            .I(N__10489));
    LocalMux I__1436 (
            .O(N__10537),
            .I(N__10482));
    LocalMux I__1435 (
            .O(N__10534),
            .I(N__10482));
    LocalMux I__1434 (
            .O(N__10531),
            .I(N__10482));
    LocalMux I__1433 (
            .O(N__10528),
            .I(N__10477));
    LocalMux I__1432 (
            .O(N__10519),
            .I(N__10477));
    InMux I__1431 (
            .O(N__10518),
            .I(N__10472));
    InMux I__1430 (
            .O(N__10517),
            .I(N__10472));
    InMux I__1429 (
            .O(N__10516),
            .I(N__10467));
    InMux I__1428 (
            .O(N__10515),
            .I(N__10467));
    InMux I__1427 (
            .O(N__10514),
            .I(N__10456));
    InMux I__1426 (
            .O(N__10513),
            .I(N__10456));
    InMux I__1425 (
            .O(N__10512),
            .I(N__10456));
    InMux I__1424 (
            .O(N__10511),
            .I(N__10456));
    InMux I__1423 (
            .O(N__10510),
            .I(N__10456));
    Span4Mux_h I__1422 (
            .O(N__10507),
            .I(N__10451));
    LocalMux I__1421 (
            .O(N__10494),
            .I(N__10451));
    LocalMux I__1420 (
            .O(N__10489),
            .I(N__10444));
    Span4Mux_v I__1419 (
            .O(N__10482),
            .I(N__10444));
    Span4Mux_h I__1418 (
            .O(N__10477),
            .I(N__10444));
    LocalMux I__1417 (
            .O(N__10472),
            .I(\b2v_inst.data_a_escribir10_THRU_CO ));
    LocalMux I__1416 (
            .O(N__10467),
            .I(\b2v_inst.data_a_escribir10_THRU_CO ));
    LocalMux I__1415 (
            .O(N__10456),
            .I(\b2v_inst.data_a_escribir10_THRU_CO ));
    Odrv4 I__1414 (
            .O(N__10451),
            .I(\b2v_inst.data_a_escribir10_THRU_CO ));
    Odrv4 I__1413 (
            .O(N__10444),
            .I(\b2v_inst.data_a_escribir10_THRU_CO ));
    InMux I__1412 (
            .O(N__10433),
            .I(N__10420));
    InMux I__1411 (
            .O(N__10432),
            .I(N__10420));
    InMux I__1410 (
            .O(N__10431),
            .I(N__10414));
    InMux I__1409 (
            .O(N__10430),
            .I(N__10414));
    InMux I__1408 (
            .O(N__10429),
            .I(N__10411));
    InMux I__1407 (
            .O(N__10428),
            .I(N__10406));
    InMux I__1406 (
            .O(N__10427),
            .I(N__10406));
    InMux I__1405 (
            .O(N__10426),
            .I(N__10401));
    InMux I__1404 (
            .O(N__10425),
            .I(N__10401));
    LocalMux I__1403 (
            .O(N__10420),
            .I(N__10398));
    InMux I__1402 (
            .O(N__10419),
            .I(N__10395));
    LocalMux I__1401 (
            .O(N__10414),
            .I(N__10392));
    LocalMux I__1400 (
            .O(N__10411),
            .I(N__10383));
    LocalMux I__1399 (
            .O(N__10406),
            .I(N__10383));
    LocalMux I__1398 (
            .O(N__10401),
            .I(N__10383));
    Span4Mux_h I__1397 (
            .O(N__10398),
            .I(N__10383));
    LocalMux I__1396 (
            .O(N__10395),
            .I(\b2v_inst.N_264 ));
    Odrv4 I__1395 (
            .O(N__10392),
            .I(\b2v_inst.N_264 ));
    Odrv4 I__1394 (
            .O(N__10383),
            .I(\b2v_inst.N_264 ));
    InMux I__1393 (
            .O(N__10376),
            .I(N__10373));
    LocalMux I__1392 (
            .O(N__10373),
            .I(N__10370));
    Odrv4 I__1391 (
            .O(N__10370),
            .I(\b2v_inst.un1_reg_anterior_iv_0_0_0_7 ));
    CascadeMux I__1390 (
            .O(N__10367),
            .I(\b2v_inst.un1_reg_anterior_iv_0_0_3_0_7_cascade_ ));
    InMux I__1389 (
            .O(N__10364),
            .I(N__10361));
    LocalMux I__1388 (
            .O(N__10361),
            .I(N__10358));
    Span4Mux_h I__1387 (
            .O(N__10358),
            .I(N__10355));
    Odrv4 I__1386 (
            .O(N__10355),
            .I(\b2v_inst.un1_reg_anterior_iv_0_0_2_0_tz_7 ));
    CEMux I__1385 (
            .O(N__10352),
            .I(N__10346));
    CEMux I__1384 (
            .O(N__10351),
            .I(N__10343));
    CEMux I__1383 (
            .O(N__10350),
            .I(N__10340));
    CEMux I__1382 (
            .O(N__10349),
            .I(N__10337));
    LocalMux I__1381 (
            .O(N__10346),
            .I(N__10334));
    LocalMux I__1380 (
            .O(N__10343),
            .I(N__10330));
    LocalMux I__1379 (
            .O(N__10340),
            .I(N__10327));
    LocalMux I__1378 (
            .O(N__10337),
            .I(N__10324));
    Span4Mux_v I__1377 (
            .O(N__10334),
            .I(N__10321));
    CEMux I__1376 (
            .O(N__10333),
            .I(N__10318));
    Span4Mux_h I__1375 (
            .O(N__10330),
            .I(N__10315));
    Span4Mux_h I__1374 (
            .O(N__10327),
            .I(N__10312));
    Span4Mux_h I__1373 (
            .O(N__10324),
            .I(N__10307));
    Span4Mux_v I__1372 (
            .O(N__10321),
            .I(N__10307));
    LocalMux I__1371 (
            .O(N__10318),
            .I(N__10302));
    Span4Mux_h I__1370 (
            .O(N__10315),
            .I(N__10302));
    Odrv4 I__1369 (
            .O(N__10312),
            .I(\b2v_inst.un1_reset_inv_2_0 ));
    Odrv4 I__1368 (
            .O(N__10307),
            .I(\b2v_inst.un1_reset_inv_2_0 ));
    Odrv4 I__1367 (
            .O(N__10302),
            .I(\b2v_inst.un1_reset_inv_2_0 ));
    InMux I__1366 (
            .O(N__10295),
            .I(N__10291));
    InMux I__1365 (
            .O(N__10294),
            .I(N__10288));
    LocalMux I__1364 (
            .O(N__10291),
            .I(N__10283));
    LocalMux I__1363 (
            .O(N__10288),
            .I(N__10279));
    InMux I__1362 (
            .O(N__10287),
            .I(N__10276));
    InMux I__1361 (
            .O(N__10286),
            .I(N__10273));
    Span4Mux_v I__1360 (
            .O(N__10283),
            .I(N__10270));
    InMux I__1359 (
            .O(N__10282),
            .I(N__10267));
    Span4Mux_h I__1358 (
            .O(N__10279),
            .I(N__10264));
    LocalMux I__1357 (
            .O(N__10276),
            .I(N__10259));
    LocalMux I__1356 (
            .O(N__10273),
            .I(N__10259));
    Odrv4 I__1355 (
            .O(N__10270),
            .I(\b2v_inst.reg_ancho_1Z0Z_0 ));
    LocalMux I__1354 (
            .O(N__10267),
            .I(\b2v_inst.reg_ancho_1Z0Z_0 ));
    Odrv4 I__1353 (
            .O(N__10264),
            .I(\b2v_inst.reg_ancho_1Z0Z_0 ));
    Odrv4 I__1352 (
            .O(N__10259),
            .I(\b2v_inst.reg_ancho_1Z0Z_0 ));
    InMux I__1351 (
            .O(N__10250),
            .I(N__10247));
    LocalMux I__1350 (
            .O(N__10247),
            .I(N__10243));
    InMux I__1349 (
            .O(N__10246),
            .I(N__10239));
    Span4Mux_v I__1348 (
            .O(N__10243),
            .I(N__10236));
    InMux I__1347 (
            .O(N__10242),
            .I(N__10233));
    LocalMux I__1346 (
            .O(N__10239),
            .I(N__10230));
    Odrv4 I__1345 (
            .O(N__10236),
            .I(\b2v_inst.reg_ancho_3Z0Z_0 ));
    LocalMux I__1344 (
            .O(N__10233),
            .I(\b2v_inst.reg_ancho_3Z0Z_0 ));
    Odrv4 I__1343 (
            .O(N__10230),
            .I(\b2v_inst.reg_ancho_3Z0Z_0 ));
    CascadeMux I__1342 (
            .O(N__10223),
            .I(N_458_cascade_));
    CascadeMux I__1341 (
            .O(N__10220),
            .I(\b2v_inst.N_429_cascade_ ));
    InMux I__1340 (
            .O(N__10217),
            .I(N__10214));
    LocalMux I__1339 (
            .O(N__10214),
            .I(N__10211));
    Span4Mux_h I__1338 (
            .O(N__10211),
            .I(N__10203));
    InMux I__1337 (
            .O(N__10210),
            .I(N__10198));
    InMux I__1336 (
            .O(N__10209),
            .I(N__10198));
    InMux I__1335 (
            .O(N__10208),
            .I(N__10191));
    InMux I__1334 (
            .O(N__10207),
            .I(N__10191));
    InMux I__1333 (
            .O(N__10206),
            .I(N__10191));
    Odrv4 I__1332 (
            .O(N__10203),
            .I(\b2v_inst.un1_pix_count_anterior_0_N_2_THRU_CO ));
    LocalMux I__1331 (
            .O(N__10198),
            .I(\b2v_inst.un1_pix_count_anterior_0_N_2_THRU_CO ));
    LocalMux I__1330 (
            .O(N__10191),
            .I(\b2v_inst.un1_pix_count_anterior_0_N_2_THRU_CO ));
    InMux I__1329 (
            .O(N__10184),
            .I(N__10175));
    InMux I__1328 (
            .O(N__10183),
            .I(N__10175));
    InMux I__1327 (
            .O(N__10182),
            .I(N__10175));
    LocalMux I__1326 (
            .O(N__10175),
            .I(\b2v_inst.stateZ0Z_3 ));
    CascadeMux I__1325 (
            .O(N__10172),
            .I(N__10168));
    IoInMux I__1324 (
            .O(N__10171),
            .I(N__10165));
    InMux I__1323 (
            .O(N__10168),
            .I(N__10161));
    LocalMux I__1322 (
            .O(N__10165),
            .I(N__10158));
    InMux I__1321 (
            .O(N__10164),
            .I(N__10154));
    LocalMux I__1320 (
            .O(N__10161),
            .I(N__10151));
    IoSpan4Mux I__1319 (
            .O(N__10158),
            .I(N__10148));
    CascadeMux I__1318 (
            .O(N__10157),
            .I(N__10145));
    LocalMux I__1317 (
            .O(N__10154),
            .I(N__10140));
    Span4Mux_v I__1316 (
            .O(N__10151),
            .I(N__10137));
    Sp12to4 I__1315 (
            .O(N__10148),
            .I(N__10134));
    InMux I__1314 (
            .O(N__10145),
            .I(N__10131));
    InMux I__1313 (
            .O(N__10144),
            .I(N__10126));
    InMux I__1312 (
            .O(N__10143),
            .I(N__10126));
    Span4Mux_v I__1311 (
            .O(N__10140),
            .I(N__10123));
    Span4Mux_h I__1310 (
            .O(N__10137),
            .I(N__10120));
    Span12Mux_v I__1309 (
            .O(N__10134),
            .I(N__10117));
    LocalMux I__1308 (
            .O(N__10131),
            .I(\b2v_inst.stateZ0Z_2 ));
    LocalMux I__1307 (
            .O(N__10126),
            .I(\b2v_inst.stateZ0Z_2 ));
    Odrv4 I__1306 (
            .O(N__10123),
            .I(\b2v_inst.stateZ0Z_2 ));
    Odrv4 I__1305 (
            .O(N__10120),
            .I(\b2v_inst.stateZ0Z_2 ));
    Odrv12 I__1304 (
            .O(N__10117),
            .I(\b2v_inst.stateZ0Z_2 ));
    CascadeMux I__1303 (
            .O(N__10106),
            .I(N__10103));
    InMux I__1302 (
            .O(N__10103),
            .I(N__10100));
    LocalMux I__1301 (
            .O(N__10100),
            .I(N__10097));
    Odrv4 I__1300 (
            .O(N__10097),
            .I(\b2v_inst.data_a_escribir9_4_and ));
    InMux I__1299 (
            .O(N__10094),
            .I(N__10091));
    LocalMux I__1298 (
            .O(N__10091),
            .I(N__10088));
    Span4Mux_v I__1297 (
            .O(N__10088),
            .I(N__10085));
    Odrv4 I__1296 (
            .O(N__10085),
            .I(SYNTHESIZED_WIRE_3_3));
    InMux I__1295 (
            .O(N__10082),
            .I(N__10079));
    LocalMux I__1294 (
            .O(N__10079),
            .I(N__10076));
    Span4Mux_h I__1293 (
            .O(N__10076),
            .I(N__10073));
    Odrv4 I__1292 (
            .O(N__10073),
            .I(SYNTHESIZED_WIRE_3_4));
    InMux I__1291 (
            .O(N__10070),
            .I(N__10067));
    LocalMux I__1290 (
            .O(N__10067),
            .I(N__10064));
    Span4Mux_h I__1289 (
            .O(N__10064),
            .I(N__10061));
    Odrv4 I__1288 (
            .O(N__10061),
            .I(SYNTHESIZED_WIRE_3_5));
    CascadeMux I__1287 (
            .O(N__10058),
            .I(N__10055));
    InMux I__1286 (
            .O(N__10055),
            .I(N__10052));
    LocalMux I__1285 (
            .O(N__10052),
            .I(N__10049));
    Span4Mux_h I__1284 (
            .O(N__10049),
            .I(N__10046));
    Odrv4 I__1283 (
            .O(N__10046),
            .I(SYNTHESIZED_WIRE_3_6));
    CascadeMux I__1282 (
            .O(N__10043),
            .I(N__10040));
    InMux I__1281 (
            .O(N__10040),
            .I(N__10037));
    LocalMux I__1280 (
            .O(N__10037),
            .I(N__10034));
    Span4Mux_v I__1279 (
            .O(N__10034),
            .I(N__10031));
    Odrv4 I__1278 (
            .O(N__10031),
            .I(SYNTHESIZED_WIRE_3_7));
    CEMux I__1277 (
            .O(N__10028),
            .I(N__10024));
    CascadeMux I__1276 (
            .O(N__10027),
            .I(N__10020));
    LocalMux I__1275 (
            .O(N__10024),
            .I(N__10017));
    InMux I__1274 (
            .O(N__10023),
            .I(N__10014));
    InMux I__1273 (
            .O(N__10020),
            .I(N__10011));
    Span4Mux_h I__1272 (
            .O(N__10017),
            .I(N__10008));
    LocalMux I__1271 (
            .O(N__10014),
            .I(N__10005));
    LocalMux I__1270 (
            .O(N__10011),
            .I(N__10002));
    Odrv4 I__1269 (
            .O(N__10008),
            .I(\b2v_inst4.pix_count_int_0_sqmuxa ));
    Odrv4 I__1268 (
            .O(N__10005),
            .I(\b2v_inst4.pix_count_int_0_sqmuxa ));
    Odrv4 I__1267 (
            .O(N__10002),
            .I(\b2v_inst4.pix_count_int_0_sqmuxa ));
    CascadeMux I__1266 (
            .O(N__9995),
            .I(\b2v_inst.we_0_a2_0_a2_4_cascade_ ));
    CEMux I__1265 (
            .O(N__9992),
            .I(N__9989));
    LocalMux I__1264 (
            .O(N__9989),
            .I(N__9986));
    Span4Mux_v I__1263 (
            .O(N__9986),
            .I(N__9983));
    Odrv4 I__1262 (
            .O(N__9983),
            .I(SYNTHESIZED_WIRE_4));
    InMux I__1261 (
            .O(N__9980),
            .I(N__9977));
    LocalMux I__1260 (
            .O(N__9977),
            .I(\b2v_inst.we_0_a2_0_a2_3 ));
    CascadeMux I__1259 (
            .O(N__9974),
            .I(\b2v_inst3.un1_m2_0_a2_2_cascade_ ));
    CascadeMux I__1258 (
            .O(N__9971),
            .I(N__9967));
    CascadeMux I__1257 (
            .O(N__9970),
            .I(N__9964));
    InMux I__1256 (
            .O(N__9967),
            .I(N__9959));
    InMux I__1255 (
            .O(N__9964),
            .I(N__9959));
    LocalMux I__1254 (
            .O(N__9959),
            .I(\b2v_inst3.un1_cycle_counter_5_c5 ));
    CascadeMux I__1253 (
            .O(N__9956),
            .I(\b2v_inst3.un1_cycle_counter_5_c5_cascade_ ));
    InMux I__1252 (
            .O(N__9953),
            .I(N__9950));
    LocalMux I__1251 (
            .O(N__9950),
            .I(N__9947));
    Span4Mux_v I__1250 (
            .O(N__9947),
            .I(N__9943));
    InMux I__1249 (
            .O(N__9946),
            .I(N__9940));
    Odrv4 I__1248 (
            .O(N__9943),
            .I(SYNTHESIZED_WIRE_10_0));
    LocalMux I__1247 (
            .O(N__9940),
            .I(SYNTHESIZED_WIRE_10_0));
    InMux I__1246 (
            .O(N__9935),
            .I(N__9932));
    LocalMux I__1245 (
            .O(N__9932),
            .I(N__9929));
    Span4Mux_h I__1244 (
            .O(N__9929),
            .I(N__9926));
    Odrv4 I__1243 (
            .O(N__9926),
            .I(SYNTHESIZED_WIRE_3_0));
    InMux I__1242 (
            .O(N__9923),
            .I(N__9920));
    LocalMux I__1241 (
            .O(N__9920),
            .I(N__9917));
    Span4Mux_h I__1240 (
            .O(N__9917),
            .I(N__9914));
    Odrv4 I__1239 (
            .O(N__9914),
            .I(SYNTHESIZED_WIRE_3_1));
    InMux I__1238 (
            .O(N__9911),
            .I(N__9908));
    LocalMux I__1237 (
            .O(N__9908),
            .I(N__9905));
    Span4Mux_v I__1236 (
            .O(N__9905),
            .I(N__9902));
    Odrv4 I__1235 (
            .O(N__9902),
            .I(SYNTHESIZED_WIRE_3_2));
    InMux I__1234 (
            .O(N__9899),
            .I(N__9896));
    LocalMux I__1233 (
            .O(N__9896),
            .I(\b2v_inst.un1_reg_anterior_iv_0_0_2_tz_4 ));
    CascadeMux I__1232 (
            .O(N__9893),
            .I(\b2v_inst3.fsm_state_ns_0_0_0_1_cascade_ ));
    CascadeMux I__1231 (
            .O(N__9890),
            .I(N_230_cascade_));
    InMux I__1230 (
            .O(N__9887),
            .I(N__9884));
    LocalMux I__1229 (
            .O(N__9884),
            .I(\b2v_inst3.N_434 ));
    InMux I__1228 (
            .O(N__9881),
            .I(N__9878));
    LocalMux I__1227 (
            .O(N__9878),
            .I(\b2v_inst3.N_490 ));
    CascadeMux I__1226 (
            .O(N__9875),
            .I(\b2v_inst3.fsm_state_ns_i_i_1_0_cascade_ ));
    CascadeMux I__1225 (
            .O(N__9872),
            .I(N__9868));
    InMux I__1224 (
            .O(N__9871),
            .I(N__9865));
    InMux I__1223 (
            .O(N__9868),
            .I(N__9862));
    LocalMux I__1222 (
            .O(N__9865),
            .I(N__9859));
    LocalMux I__1221 (
            .O(N__9862),
            .I(\b2v_inst.reg_anterior_i_1 ));
    Odrv4 I__1220 (
            .O(N__9859),
            .I(\b2v_inst.reg_anterior_i_1 ));
    CascadeMux I__1219 (
            .O(N__9854),
            .I(N__9850));
    InMux I__1218 (
            .O(N__9853),
            .I(N__9847));
    InMux I__1217 (
            .O(N__9850),
            .I(N__9844));
    LocalMux I__1216 (
            .O(N__9847),
            .I(N__9841));
    LocalMux I__1215 (
            .O(N__9844),
            .I(\b2v_inst.reg_anterior_i_2 ));
    Odrv4 I__1214 (
            .O(N__9841),
            .I(\b2v_inst.reg_anterior_i_2 ));
    CascadeMux I__1213 (
            .O(N__9836),
            .I(N__9832));
    InMux I__1212 (
            .O(N__9835),
            .I(N__9829));
    InMux I__1211 (
            .O(N__9832),
            .I(N__9826));
    LocalMux I__1210 (
            .O(N__9829),
            .I(N__9823));
    LocalMux I__1209 (
            .O(N__9826),
            .I(\b2v_inst.reg_anterior_i_3 ));
    Odrv4 I__1208 (
            .O(N__9823),
            .I(\b2v_inst.reg_anterior_i_3 ));
    CascadeMux I__1207 (
            .O(N__9818),
            .I(N__9814));
    CascadeMux I__1206 (
            .O(N__9817),
            .I(N__9811));
    InMux I__1205 (
            .O(N__9814),
            .I(N__9808));
    InMux I__1204 (
            .O(N__9811),
            .I(N__9805));
    LocalMux I__1203 (
            .O(N__9808),
            .I(N__9802));
    LocalMux I__1202 (
            .O(N__9805),
            .I(\b2v_inst.reg_anterior_i_4 ));
    Odrv4 I__1201 (
            .O(N__9802),
            .I(\b2v_inst.reg_anterior_i_4 ));
    CascadeMux I__1200 (
            .O(N__9797),
            .I(N__9793));
    CascadeMux I__1199 (
            .O(N__9796),
            .I(N__9790));
    InMux I__1198 (
            .O(N__9793),
            .I(N__9787));
    InMux I__1197 (
            .O(N__9790),
            .I(N__9784));
    LocalMux I__1196 (
            .O(N__9787),
            .I(N__9781));
    LocalMux I__1195 (
            .O(N__9784),
            .I(\b2v_inst.reg_anterior_i_5 ));
    Odrv4 I__1194 (
            .O(N__9781),
            .I(\b2v_inst.reg_anterior_i_5 ));
    CascadeMux I__1193 (
            .O(N__9776),
            .I(N__9772));
    CascadeMux I__1192 (
            .O(N__9775),
            .I(N__9769));
    InMux I__1191 (
            .O(N__9772),
            .I(N__9766));
    InMux I__1190 (
            .O(N__9769),
            .I(N__9763));
    LocalMux I__1189 (
            .O(N__9766),
            .I(N__9760));
    LocalMux I__1188 (
            .O(N__9763),
            .I(N__9757));
    Odrv4 I__1187 (
            .O(N__9760),
            .I(\b2v_inst.reg_anterior_i_6 ));
    Odrv4 I__1186 (
            .O(N__9757),
            .I(\b2v_inst.reg_anterior_i_6 ));
    InMux I__1185 (
            .O(N__9752),
            .I(N__9748));
    CascadeMux I__1184 (
            .O(N__9751),
            .I(N__9745));
    LocalMux I__1183 (
            .O(N__9748),
            .I(N__9742));
    InMux I__1182 (
            .O(N__9745),
            .I(N__9739));
    Span4Mux_h I__1181 (
            .O(N__9742),
            .I(N__9736));
    LocalMux I__1180 (
            .O(N__9739),
            .I(\b2v_inst.reg_anterior_i_7 ));
    Odrv4 I__1179 (
            .O(N__9736),
            .I(\b2v_inst.reg_anterior_i_7 ));
    InMux I__1178 (
            .O(N__9731),
            .I(N__9728));
    LocalMux I__1177 (
            .O(N__9728),
            .I(N__9724));
    InMux I__1176 (
            .O(N__9727),
            .I(N__9721));
    Odrv4 I__1175 (
            .O(N__9724),
            .I(\b2v_inst.valor_max_final53_THRU_CO ));
    LocalMux I__1174 (
            .O(N__9721),
            .I(\b2v_inst.valor_max_final53_THRU_CO ));
    CascadeMux I__1173 (
            .O(N__9716),
            .I(N__9713));
    InMux I__1172 (
            .O(N__9713),
            .I(N__9710));
    LocalMux I__1171 (
            .O(N__9710),
            .I(\b2v_inst.un1_m3_0_m3_ns_1 ));
    InMux I__1170 (
            .O(N__9707),
            .I(bfn_3_20_0_));
    InMux I__1169 (
            .O(N__9704),
            .I(N__9701));
    LocalMux I__1168 (
            .O(N__9701),
            .I(N__9698));
    Odrv12 I__1167 (
            .O(N__9698),
            .I(\b2v_inst.N_497 ));
    InMux I__1166 (
            .O(N__9695),
            .I(N__9692));
    LocalMux I__1165 (
            .O(N__9692),
            .I(N__9689));
    Odrv4 I__1164 (
            .O(N__9689),
            .I(\b2v_inst.un1_reg_anterior_iv_0_0_2_tz_2 ));
    CascadeMux I__1163 (
            .O(N__9686),
            .I(\b2v_inst.data_a_escribir_RNO_1Z0Z_2_cascade_ ));
    InMux I__1162 (
            .O(N__9683),
            .I(N__9680));
    LocalMux I__1161 (
            .O(N__9680),
            .I(\b2v_inst.un1_reg_anterior_iv_0_0_1_2 ));
    CascadeMux I__1160 (
            .O(N__9677),
            .I(\b2v_inst.data_a_escribir_RNO_4Z0Z_5_cascade_ ));
    CascadeMux I__1159 (
            .O(N__9674),
            .I(\b2v_inst.un1_reg_anterior_iv_0_0_2_1_5_cascade_ ));
    InMux I__1158 (
            .O(N__9671),
            .I(N__9663));
    InMux I__1157 (
            .O(N__9670),
            .I(N__9663));
    InMux I__1156 (
            .O(N__9669),
            .I(N__9660));
    InMux I__1155 (
            .O(N__9668),
            .I(N__9657));
    LocalMux I__1154 (
            .O(N__9663),
            .I(\b2v_inst.un1_reg_anterior_iv_0_0_a2_4_0_1 ));
    LocalMux I__1153 (
            .O(N__9660),
            .I(\b2v_inst.un1_reg_anterior_iv_0_0_a2_4_0_1 ));
    LocalMux I__1152 (
            .O(N__9657),
            .I(\b2v_inst.un1_reg_anterior_iv_0_0_a2_4_0_1 ));
    InMux I__1151 (
            .O(N__9650),
            .I(N__9647));
    LocalMux I__1150 (
            .O(N__9647),
            .I(N__9644));
    Span4Mux_h I__1149 (
            .O(N__9644),
            .I(N__9641));
    Odrv4 I__1148 (
            .O(N__9641),
            .I(\b2v_inst.un1_reg_anterior_iv_0_0_0_5 ));
    CascadeMux I__1147 (
            .O(N__9638),
            .I(\b2v_inst.data_a_escribir_RNO_0Z0Z_5_cascade_ ));
    InMux I__1146 (
            .O(N__9635),
            .I(N__9632));
    LocalMux I__1145 (
            .O(N__9632),
            .I(\b2v_inst.data_a_escribir_RNO_1Z0Z_5 ));
    CascadeMux I__1144 (
            .O(N__9629),
            .I(N__9625));
    InMux I__1143 (
            .O(N__9628),
            .I(N__9622));
    InMux I__1142 (
            .O(N__9625),
            .I(N__9619));
    LocalMux I__1141 (
            .O(N__9622),
            .I(N__9616));
    LocalMux I__1140 (
            .O(N__9619),
            .I(\b2v_inst.reg_anterior_i_0 ));
    Odrv4 I__1139 (
            .O(N__9616),
            .I(\b2v_inst.reg_anterior_i_0 ));
    InMux I__1138 (
            .O(N__9611),
            .I(N__9608));
    LocalMux I__1137 (
            .O(N__9608),
            .I(N__9605));
    Span4Mux_h I__1136 (
            .O(N__9605),
            .I(N__9601));
    InMux I__1135 (
            .O(N__9604),
            .I(N__9598));
    Odrv4 I__1134 (
            .O(N__9601),
            .I(\b2v_inst.eventosZ0Z_1 ));
    LocalMux I__1133 (
            .O(N__9598),
            .I(\b2v_inst.eventosZ0Z_1 ));
    InMux I__1132 (
            .O(N__9593),
            .I(N__9590));
    LocalMux I__1131 (
            .O(N__9590),
            .I(N__9586));
    InMux I__1130 (
            .O(N__9589),
            .I(N__9583));
    Span12Mux_s11_v I__1129 (
            .O(N__9586),
            .I(N__9580));
    LocalMux I__1128 (
            .O(N__9583),
            .I(\b2v_inst.eventosZ0Z_6 ));
    Odrv12 I__1127 (
            .O(N__9580),
            .I(\b2v_inst.eventosZ0Z_6 ));
    CascadeMux I__1126 (
            .O(N__9575),
            .I(\b2v_inst.un1_reg_anterior_iv_0_0_2_1_1_cascade_ ));
    CascadeMux I__1125 (
            .O(N__9572),
            .I(\b2v_inst.data_a_escribir_RNO_4Z0Z_1_cascade_ ));
    InMux I__1124 (
            .O(N__9569),
            .I(N__9566));
    LocalMux I__1123 (
            .O(N__9566),
            .I(\b2v_inst.un1_reg_anterior_iv_0_0_0_1 ));
    InMux I__1122 (
            .O(N__9563),
            .I(N__9560));
    LocalMux I__1121 (
            .O(N__9560),
            .I(\b2v_inst.data_a_escribir_RNO_0Z0Z_1 ));
    CascadeMux I__1120 (
            .O(N__9557),
            .I(\b2v_inst.data_a_escribir_RNO_1Z0Z_1_cascade_ ));
    InMux I__1119 (
            .O(N__9554),
            .I(N__9551));
    LocalMux I__1118 (
            .O(N__9551),
            .I(N__9548));
    Span4Mux_h I__1117 (
            .O(N__9548),
            .I(N__9545));
    Odrv4 I__1116 (
            .O(N__9545),
            .I(\b2v_inst.data_a_escribir9_2_and ));
    InMux I__1115 (
            .O(N__9542),
            .I(N__9539));
    LocalMux I__1114 (
            .O(N__9539),
            .I(N__9536));
    Odrv4 I__1113 (
            .O(N__9536),
            .I(\b2v_inst.data_a_escribir9_3_and ));
    InMux I__1112 (
            .O(N__9533),
            .I(bfn_3_16_0_));
    InMux I__1111 (
            .O(N__9530),
            .I(N__9527));
    LocalMux I__1110 (
            .O(N__9527),
            .I(N__9523));
    InMux I__1109 (
            .O(N__9526),
            .I(N__9520));
    Span4Mux_h I__1108 (
            .O(N__9523),
            .I(N__9517));
    LocalMux I__1107 (
            .O(N__9520),
            .I(\b2v_inst.eventosZ0Z_7 ));
    Odrv4 I__1106 (
            .O(N__9517),
            .I(\b2v_inst.eventosZ0Z_7 ));
    InMux I__1105 (
            .O(N__9512),
            .I(N__9506));
    InMux I__1104 (
            .O(N__9511),
            .I(N__9499));
    InMux I__1103 (
            .O(N__9510),
            .I(N__9499));
    InMux I__1102 (
            .O(N__9509),
            .I(N__9499));
    LocalMux I__1101 (
            .O(N__9506),
            .I(SYNTHESIZED_WIRE_2_7));
    LocalMux I__1100 (
            .O(N__9499),
            .I(SYNTHESIZED_WIRE_2_7));
    InMux I__1099 (
            .O(N__9494),
            .I(N__9491));
    LocalMux I__1098 (
            .O(N__9491),
            .I(\b2v_inst4.pix_count_int_RNO_0Z0Z_7 ));
    InMux I__1097 (
            .O(N__9488),
            .I(\b2v_inst4.un1_pix_count_int_cry_6 ));
    InMux I__1096 (
            .O(N__9485),
            .I(N__9479));
    InMux I__1095 (
            .O(N__9484),
            .I(N__9472));
    InMux I__1094 (
            .O(N__9483),
            .I(N__9472));
    InMux I__1093 (
            .O(N__9482),
            .I(N__9472));
    LocalMux I__1092 (
            .O(N__9479),
            .I(SYNTHESIZED_WIRE_2_8));
    LocalMux I__1091 (
            .O(N__9472),
            .I(SYNTHESIZED_WIRE_2_8));
    InMux I__1090 (
            .O(N__9467),
            .I(N__9464));
    LocalMux I__1089 (
            .O(N__9464),
            .I(\b2v_inst4.pix_count_int_RNO_0Z0Z_8 ));
    InMux I__1088 (
            .O(N__9461),
            .I(bfn_3_14_0_));
    InMux I__1087 (
            .O(N__9458),
            .I(\b2v_inst4.un1_pix_count_int_cry_8 ));
    InMux I__1086 (
            .O(N__9455),
            .I(N__9447));
    InMux I__1085 (
            .O(N__9454),
            .I(N__9447));
    InMux I__1084 (
            .O(N__9453),
            .I(N__9444));
    InMux I__1083 (
            .O(N__9452),
            .I(N__9441));
    LocalMux I__1082 (
            .O(N__9447),
            .I(N__9436));
    LocalMux I__1081 (
            .O(N__9444),
            .I(N__9436));
    LocalMux I__1080 (
            .O(N__9441),
            .I(SYNTHESIZED_WIRE_2_10));
    Odrv4 I__1079 (
            .O(N__9436),
            .I(SYNTHESIZED_WIRE_2_10));
    InMux I__1078 (
            .O(N__9431),
            .I(\b2v_inst4.un1_pix_count_int_cry_9 ));
    InMux I__1077 (
            .O(N__9428),
            .I(N__9422));
    InMux I__1076 (
            .O(N__9427),
            .I(N__9419));
    InMux I__1075 (
            .O(N__9426),
            .I(N__9414));
    InMux I__1074 (
            .O(N__9425),
            .I(N__9414));
    LocalMux I__1073 (
            .O(N__9422),
            .I(SYNTHESIZED_WIRE_2_11));
    LocalMux I__1072 (
            .O(N__9419),
            .I(SYNTHESIZED_WIRE_2_11));
    LocalMux I__1071 (
            .O(N__9414),
            .I(SYNTHESIZED_WIRE_2_11));
    InMux I__1070 (
            .O(N__9407),
            .I(N__9404));
    LocalMux I__1069 (
            .O(N__9404),
            .I(\b2v_inst4.pix_count_int_RNO_0Z0Z_11 ));
    InMux I__1068 (
            .O(N__9401),
            .I(\b2v_inst4.un1_pix_count_int_cry_10 ));
    CascadeMux I__1067 (
            .O(N__9398),
            .I(N__9393));
    InMux I__1066 (
            .O(N__9397),
            .I(N__9389));
    InMux I__1065 (
            .O(N__9396),
            .I(N__9386));
    InMux I__1064 (
            .O(N__9393),
            .I(N__9383));
    InMux I__1063 (
            .O(N__9392),
            .I(N__9380));
    LocalMux I__1062 (
            .O(N__9389),
            .I(SYNTHESIZED_WIRE_2_12));
    LocalMux I__1061 (
            .O(N__9386),
            .I(SYNTHESIZED_WIRE_2_12));
    LocalMux I__1060 (
            .O(N__9383),
            .I(SYNTHESIZED_WIRE_2_12));
    LocalMux I__1059 (
            .O(N__9380),
            .I(SYNTHESIZED_WIRE_2_12));
    InMux I__1058 (
            .O(N__9371),
            .I(\b2v_inst4.un1_pix_count_int_cry_11 ));
    InMux I__1057 (
            .O(N__9368),
            .I(N__9365));
    LocalMux I__1056 (
            .O(N__9365),
            .I(\b2v_inst4.pix_count_int_RNO_0Z0Z_12 ));
    InMux I__1055 (
            .O(N__9362),
            .I(N__9359));
    LocalMux I__1054 (
            .O(N__9359),
            .I(\b2v_inst.data_a_escribir9_0_and ));
    InMux I__1053 (
            .O(N__9356),
            .I(N__9353));
    LocalMux I__1052 (
            .O(N__9353),
            .I(\b2v_inst.data_a_escribir9_1_and ));
    CascadeMux I__1051 (
            .O(N__9350),
            .I(N__9347));
    InMux I__1050 (
            .O(N__9347),
            .I(N__9344));
    LocalMux I__1049 (
            .O(N__9344),
            .I(\b2v_inst.pix_count_anteriorZ0Z_11 ));
    CEMux I__1048 (
            .O(N__9341),
            .I(N__9323));
    CEMux I__1047 (
            .O(N__9340),
            .I(N__9323));
    CEMux I__1046 (
            .O(N__9339),
            .I(N__9323));
    CEMux I__1045 (
            .O(N__9338),
            .I(N__9323));
    CEMux I__1044 (
            .O(N__9337),
            .I(N__9323));
    CEMux I__1043 (
            .O(N__9336),
            .I(N__9323));
    GlobalMux I__1042 (
            .O(N__9323),
            .I(N__9320));
    gio2CtrlBuf I__1041 (
            .O(N__9320),
            .I(\b2v_inst.N_254_i_g ));
    CascadeMux I__1040 (
            .O(N__9317),
            .I(N__9314));
    InMux I__1039 (
            .O(N__9314),
            .I(N__9311));
    LocalMux I__1038 (
            .O(N__9311),
            .I(N__9305));
    InMux I__1037 (
            .O(N__9310),
            .I(N__9302));
    InMux I__1036 (
            .O(N__9309),
            .I(N__9297));
    InMux I__1035 (
            .O(N__9308),
            .I(N__9297));
    Odrv4 I__1034 (
            .O(N__9305),
            .I(SYNTHESIZED_WIRE_2_0));
    LocalMux I__1033 (
            .O(N__9302),
            .I(SYNTHESIZED_WIRE_2_0));
    LocalMux I__1032 (
            .O(N__9297),
            .I(SYNTHESIZED_WIRE_2_0));
    InMux I__1031 (
            .O(N__9290),
            .I(N__9287));
    LocalMux I__1030 (
            .O(N__9287),
            .I(\b2v_inst4.pix_count_int_RNO_0Z0Z_0 ));
    InMux I__1029 (
            .O(N__9284),
            .I(N__9278));
    InMux I__1028 (
            .O(N__9283),
            .I(N__9271));
    InMux I__1027 (
            .O(N__9282),
            .I(N__9271));
    InMux I__1026 (
            .O(N__9281),
            .I(N__9271));
    LocalMux I__1025 (
            .O(N__9278),
            .I(SYNTHESIZED_WIRE_2_1));
    LocalMux I__1024 (
            .O(N__9271),
            .I(SYNTHESIZED_WIRE_2_1));
    InMux I__1023 (
            .O(N__9266),
            .I(\b2v_inst4.un1_pix_count_int_cry_0 ));
    CascadeMux I__1022 (
            .O(N__9263),
            .I(N__9259));
    InMux I__1021 (
            .O(N__9262),
            .I(N__9252));
    InMux I__1020 (
            .O(N__9259),
            .I(N__9252));
    InMux I__1019 (
            .O(N__9258),
            .I(N__9249));
    InMux I__1018 (
            .O(N__9257),
            .I(N__9246));
    LocalMux I__1017 (
            .O(N__9252),
            .I(SYNTHESIZED_WIRE_2_2));
    LocalMux I__1016 (
            .O(N__9249),
            .I(SYNTHESIZED_WIRE_2_2));
    LocalMux I__1015 (
            .O(N__9246),
            .I(SYNTHESIZED_WIRE_2_2));
    InMux I__1014 (
            .O(N__9239),
            .I(\b2v_inst4.un1_pix_count_int_cry_1 ));
    InMux I__1013 (
            .O(N__9236),
            .I(N__9230));
    InMux I__1012 (
            .O(N__9235),
            .I(N__9223));
    InMux I__1011 (
            .O(N__9234),
            .I(N__9223));
    InMux I__1010 (
            .O(N__9233),
            .I(N__9223));
    LocalMux I__1009 (
            .O(N__9230),
            .I(SYNTHESIZED_WIRE_2_3));
    LocalMux I__1008 (
            .O(N__9223),
            .I(SYNTHESIZED_WIRE_2_3));
    InMux I__1007 (
            .O(N__9218),
            .I(N__9215));
    LocalMux I__1006 (
            .O(N__9215),
            .I(\b2v_inst4.pix_count_int_RNO_0Z0Z_3 ));
    InMux I__1005 (
            .O(N__9212),
            .I(\b2v_inst4.un1_pix_count_int_cry_2 ));
    InMux I__1004 (
            .O(N__9209),
            .I(N__9203));
    InMux I__1003 (
            .O(N__9208),
            .I(N__9196));
    InMux I__1002 (
            .O(N__9207),
            .I(N__9196));
    InMux I__1001 (
            .O(N__9206),
            .I(N__9196));
    LocalMux I__1000 (
            .O(N__9203),
            .I(SYNTHESIZED_WIRE_2_4));
    LocalMux I__999 (
            .O(N__9196),
            .I(SYNTHESIZED_WIRE_2_4));
    InMux I__998 (
            .O(N__9191),
            .I(\b2v_inst4.un1_pix_count_int_cry_3 ));
    InMux I__997 (
            .O(N__9188),
            .I(N__9182));
    InMux I__996 (
            .O(N__9187),
            .I(N__9179));
    InMux I__995 (
            .O(N__9186),
            .I(N__9174));
    InMux I__994 (
            .O(N__9185),
            .I(N__9174));
    LocalMux I__993 (
            .O(N__9182),
            .I(SYNTHESIZED_WIRE_2_5));
    LocalMux I__992 (
            .O(N__9179),
            .I(SYNTHESIZED_WIRE_2_5));
    LocalMux I__991 (
            .O(N__9174),
            .I(SYNTHESIZED_WIRE_2_5));
    InMux I__990 (
            .O(N__9167),
            .I(N__9164));
    LocalMux I__989 (
            .O(N__9164),
            .I(\b2v_inst4.pix_count_int_RNO_0Z0Z_5 ));
    InMux I__988 (
            .O(N__9161),
            .I(\b2v_inst4.un1_pix_count_int_cry_4 ));
    InMux I__987 (
            .O(N__9158),
            .I(N__9152));
    InMux I__986 (
            .O(N__9157),
            .I(N__9149));
    InMux I__985 (
            .O(N__9156),
            .I(N__9144));
    InMux I__984 (
            .O(N__9155),
            .I(N__9144));
    LocalMux I__983 (
            .O(N__9152),
            .I(SYNTHESIZED_WIRE_2_6));
    LocalMux I__982 (
            .O(N__9149),
            .I(SYNTHESIZED_WIRE_2_6));
    LocalMux I__981 (
            .O(N__9144),
            .I(SYNTHESIZED_WIRE_2_6));
    InMux I__980 (
            .O(N__9137),
            .I(\b2v_inst4.un1_pix_count_int_cry_5 ));
    InMux I__979 (
            .O(N__9134),
            .I(N__9131));
    LocalMux I__978 (
            .O(N__9131),
            .I(N__9128));
    Odrv4 I__977 (
            .O(N__9128),
            .I(\b2v_inst.N_361 ));
    InMux I__976 (
            .O(N__9125),
            .I(N__9119));
    InMux I__975 (
            .O(N__9124),
            .I(N__9119));
    LocalMux I__974 (
            .O(N__9119),
            .I(\b2v_inst.state_ns_i_i_a2_5Z0Z_6 ));
    IoInMux I__973 (
            .O(N__9116),
            .I(N__9113));
    LocalMux I__972 (
            .O(N__9113),
            .I(N__9110));
    Odrv12 I__971 (
            .O(N__9110),
            .I(\b2v_inst.N_254_i ));
    InMux I__970 (
            .O(N__9107),
            .I(N__9104));
    LocalMux I__969 (
            .O(N__9104),
            .I(\b2v_inst.pix_count_anteriorZ0Z_2 ));
    InMux I__968 (
            .O(N__9101),
            .I(N__9098));
    LocalMux I__967 (
            .O(N__9098),
            .I(\b2v_inst.un1_pix_count_anterior_0_I_27_c_RNOZ0 ));
    CascadeMux I__966 (
            .O(N__9095),
            .I(N__9092));
    InMux I__965 (
            .O(N__9092),
            .I(N__9089));
    LocalMux I__964 (
            .O(N__9089),
            .I(\b2v_inst.pix_count_anteriorZ0Z_3 ));
    InMux I__963 (
            .O(N__9086),
            .I(N__9083));
    LocalMux I__962 (
            .O(N__9083),
            .I(\b2v_inst.pix_count_anteriorZ0Z_10 ));
    InMux I__961 (
            .O(N__9080),
            .I(N__9077));
    LocalMux I__960 (
            .O(N__9077),
            .I(\b2v_inst.un1_pix_count_anterior_0_I_9_c_RNOZ0 ));
    InMux I__959 (
            .O(N__9074),
            .I(N__9071));
    LocalMux I__958 (
            .O(N__9071),
            .I(N__9068));
    Odrv12 I__957 (
            .O(N__9068),
            .I(\b2v_inst.data_a_escribir_RNO_0Z0Z_4 ));
    CascadeMux I__956 (
            .O(N__9065),
            .I(N__9062));
    InMux I__955 (
            .O(N__9062),
            .I(N__9059));
    LocalMux I__954 (
            .O(N__9059),
            .I(N__9056));
    Span4Mux_h I__953 (
            .O(N__9056),
            .I(N__9053));
    Span4Mux_v I__952 (
            .O(N__9053),
            .I(N__9050));
    Odrv4 I__951 (
            .O(N__9050),
            .I(\b2v_inst.un1_reg_anterior_iv_0_0_0_4 ));
    InMux I__950 (
            .O(N__9047),
            .I(N__9044));
    LocalMux I__949 (
            .O(N__9044),
            .I(N__9041));
    Span4Mux_h I__948 (
            .O(N__9041),
            .I(N__9038));
    Odrv4 I__947 (
            .O(N__9038),
            .I(N_211_i));
    InMux I__946 (
            .O(N__9035),
            .I(N__9032));
    LocalMux I__945 (
            .O(N__9032),
            .I(N__9029));
    Span4Mux_h I__944 (
            .O(N__9029),
            .I(N__9026));
    Span4Mux_h I__943 (
            .O(N__9026),
            .I(N__9023));
    Odrv4 I__942 (
            .O(N__9023),
            .I(N_219_i));
    InMux I__941 (
            .O(N__9020),
            .I(N__9017));
    LocalMux I__940 (
            .O(N__9017),
            .I(N__9014));
    Span12Mux_v I__939 (
            .O(N__9014),
            .I(N__9011));
    Odrv12 I__938 (
            .O(N__9011),
            .I(N_217_i));
    InMux I__937 (
            .O(N__9008),
            .I(N__9005));
    LocalMux I__936 (
            .O(N__9005),
            .I(N__9002));
    Span4Mux_h I__935 (
            .O(N__9002),
            .I(N__8999));
    Span4Mux_v I__934 (
            .O(N__8999),
            .I(N__8996));
    Odrv4 I__933 (
            .O(N__8996),
            .I(N_215_i));
    CascadeMux I__932 (
            .O(N__8993),
            .I(N__8990));
    InMux I__931 (
            .O(N__8990),
            .I(N__8987));
    LocalMux I__930 (
            .O(N__8987),
            .I(\b2v_inst.state_ns_i_i_a2_4Z0Z_6 ));
    CascadeMux I__929 (
            .O(N__8984),
            .I(\b2v_inst.state_ns_i_i_a2_4Z0Z_6_cascade_ ));
    CascadeMux I__928 (
            .O(N__8981),
            .I(\b2v_inst.N_497_cascade_ ));
    InMux I__927 (
            .O(N__8978),
            .I(N__8975));
    LocalMux I__926 (
            .O(N__8975),
            .I(\b2v_inst.N_317 ));
    InMux I__925 (
            .O(N__8972),
            .I(N__8969));
    LocalMux I__924 (
            .O(N__8969),
            .I(\b2v_inst.un1_reg_anterior_iv_0_0_a2_4_tz_1_2 ));
    InMux I__923 (
            .O(N__8966),
            .I(N__8963));
    LocalMux I__922 (
            .O(N__8963),
            .I(N__8960));
    Span4Mux_v I__921 (
            .O(N__8960),
            .I(N__8956));
    InMux I__920 (
            .O(N__8959),
            .I(N__8953));
    Odrv4 I__919 (
            .O(N__8956),
            .I(\b2v_inst.eventosZ0Z_2 ));
    LocalMux I__918 (
            .O(N__8953),
            .I(\b2v_inst.eventosZ0Z_2 ));
    CascadeMux I__917 (
            .O(N__8948),
            .I(\b2v_inst.N_320_tz_cascade_ ));
    CascadeMux I__916 (
            .O(N__8945),
            .I(\b2v_inst.un1_m3_0_m3_ns_1_cascade_ ));
    InMux I__915 (
            .O(N__8942),
            .I(N__8939));
    LocalMux I__914 (
            .O(N__8939),
            .I(N__8936));
    Odrv4 I__913 (
            .O(N__8936),
            .I(\b2v_inst.N_318 ));
    CascadeMux I__912 (
            .O(N__8933),
            .I(\b2v_inst.data_a_escribir_RNO_3Z0Z_4_cascade_ ));
    CascadeMux I__911 (
            .O(N__8930),
            .I(\b2v_inst.data_a_escribir_RNO_3Z0Z_0_cascade_ ));
    InMux I__910 (
            .O(N__8927),
            .I(N__8924));
    LocalMux I__909 (
            .O(N__8924),
            .I(N__8921));
    Span4Mux_v I__908 (
            .O(N__8921),
            .I(N__8918));
    Odrv4 I__907 (
            .O(N__8918),
            .I(\b2v_inst.un1_reg_anterior_iv_0_0_0_0 ));
    InMux I__906 (
            .O(N__8915),
            .I(N__8912));
    LocalMux I__905 (
            .O(N__8912),
            .I(\b2v_inst.un1_m3_2_0 ));
    CascadeMux I__904 (
            .O(N__8909),
            .I(\b2v_inst.data_a_escribir_RNO_1Z0Z_0_cascade_ ));
    InMux I__903 (
            .O(N__8906),
            .I(N__8903));
    LocalMux I__902 (
            .O(N__8903),
            .I(N__8900));
    Odrv4 I__901 (
            .O(N__8900),
            .I(\b2v_inst.un1_reg_anterior_iv_0_0_1_1_3 ));
    CascadeMux I__900 (
            .O(N__8897),
            .I(\b2v_inst.N_315_cascade_ ));
    InMux I__899 (
            .O(N__8894),
            .I(N__8891));
    LocalMux I__898 (
            .O(N__8891),
            .I(\b2v_inst.un1_reg_anterior_iv_0_0_1_3 ));
    CascadeMux I__897 (
            .O(N__8888),
            .I(\b2v_inst.un1_reg_anterior_iv_0_0_a2_6_0_1_cascade_ ));
    InMux I__896 (
            .O(N__8885),
            .I(N__8873));
    InMux I__895 (
            .O(N__8884),
            .I(N__8873));
    InMux I__894 (
            .O(N__8883),
            .I(N__8860));
    InMux I__893 (
            .O(N__8882),
            .I(N__8860));
    InMux I__892 (
            .O(N__8881),
            .I(N__8860));
    InMux I__891 (
            .O(N__8880),
            .I(N__8860));
    InMux I__890 (
            .O(N__8879),
            .I(N__8860));
    InMux I__889 (
            .O(N__8878),
            .I(N__8860));
    LocalMux I__888 (
            .O(N__8873),
            .I(N__8855));
    LocalMux I__887 (
            .O(N__8860),
            .I(N__8855));
    Odrv4 I__886 (
            .O(N__8855),
            .I(\b2v_inst.ignorar_anchoZ0Z_1 ));
    CascadeMux I__885 (
            .O(N__8852),
            .I(N__8849));
    InMux I__884 (
            .O(N__8849),
            .I(N__8846));
    LocalMux I__883 (
            .O(N__8846),
            .I(\b2v_inst.pix_count_anteriorZ0Z_7 ));
    InMux I__882 (
            .O(N__8843),
            .I(N__8840));
    LocalMux I__881 (
            .O(N__8840),
            .I(\b2v_inst.pix_count_anteriorZ0Z_8 ));
    InMux I__880 (
            .O(N__8837),
            .I(N__8834));
    LocalMux I__879 (
            .O(N__8834),
            .I(N__8831));
    Odrv12 I__878 (
            .O(N__8831),
            .I(\b2v_inst.un1_pix_count_anterior_0_I_51_c_RNOZ0 ));
    CascadeMux I__877 (
            .O(N__8828),
            .I(N__8825));
    InMux I__876 (
            .O(N__8825),
            .I(N__8822));
    LocalMux I__875 (
            .O(N__8822),
            .I(\b2v_inst.pix_count_anteriorZ0Z_9 ));
    CEMux I__874 (
            .O(N__8819),
            .I(N__8816));
    LocalMux I__873 (
            .O(N__8816),
            .I(N__8813));
    Span4Mux_v I__872 (
            .O(N__8813),
            .I(N__8810));
    Odrv4 I__871 (
            .O(N__8810),
            .I(\b2v_inst.un1_state_17_0 ));
    InMux I__870 (
            .O(N__8807),
            .I(N__8804));
    LocalMux I__869 (
            .O(N__8804),
            .I(\b2v_inst.pix_count_anteriorZ0Z_12 ));
    InMux I__868 (
            .O(N__8801),
            .I(N__8798));
    LocalMux I__867 (
            .O(N__8798),
            .I(N__8795));
    Odrv4 I__866 (
            .O(N__8795),
            .I(\b2v_inst.un1_pix_count_anterior_0_I_39_c_RNOZ0 ));
    InMux I__865 (
            .O(N__8792),
            .I(N__8789));
    LocalMux I__864 (
            .O(N__8789),
            .I(N__8786));
    Odrv4 I__863 (
            .O(N__8786),
            .I(\b2v_inst.un1_pix_count_anterior_0_I_21_c_RNOZ0 ));
    InMux I__862 (
            .O(N__8783),
            .I(N__8780));
    LocalMux I__861 (
            .O(N__8780),
            .I(\b2v_inst.pix_count_anteriorZ0Z_6 ));
    CascadeMux I__860 (
            .O(N__8777),
            .I(\b2v_inst4.un1_pix_count_int_0_sqmuxa_8_cascade_ ));
    InMux I__859 (
            .O(N__8774),
            .I(N__8771));
    LocalMux I__858 (
            .O(N__8771),
            .I(\b2v_inst.pix_count_anteriorZ0Z_4 ));
    CascadeMux I__857 (
            .O(N__8768),
            .I(N__8765));
    InMux I__856 (
            .O(N__8765),
            .I(N__8762));
    LocalMux I__855 (
            .O(N__8762),
            .I(\b2v_inst.pix_count_anteriorZ0Z_5 ));
    CascadeMux I__854 (
            .O(N__8759),
            .I(N__8756));
    InMux I__853 (
            .O(N__8756),
            .I(N__8753));
    LocalMux I__852 (
            .O(N__8753),
            .I(\b2v_inst.pix_count_anteriorZ0Z_1 ));
    InMux I__851 (
            .O(N__8750),
            .I(N__8747));
    LocalMux I__850 (
            .O(N__8747),
            .I(\b2v_inst.un1_pix_count_anterior_0_I_1_c_RNOZ0 ));
    InMux I__849 (
            .O(N__8744),
            .I(N__8741));
    LocalMux I__848 (
            .O(N__8741),
            .I(\b2v_inst.pix_count_anteriorZ0Z_0 ));
    InMux I__847 (
            .O(N__8738),
            .I(\b2v_inst.un1_pix_count_anterior_0_N_2 ));
    InMux I__846 (
            .O(N__8735),
            .I(N__8732));
    LocalMux I__845 (
            .O(N__8732),
            .I(\b2v_inst.un1_pix_count_anterior_0_I_15_c_RNOZ0 ));
    InMux I__844 (
            .O(N__8729),
            .I(bfn_1_20_0_));
    InMux I__843 (
            .O(N__8726),
            .I(N__8723));
    LocalMux I__842 (
            .O(N__8723),
            .I(N__8720));
    Span12Mux_v I__841 (
            .O(N__8720),
            .I(N__8717));
    Odrv12 I__840 (
            .O(N__8717),
            .I(\b2v_inst.g0_10_1 ));
    InMux I__839 (
            .O(N__8714),
            .I(N__8711));
    LocalMux I__838 (
            .O(N__8711),
            .I(N__8708));
    Span12Mux_s8_v I__837 (
            .O(N__8708),
            .I(N__8705));
    Odrv12 I__836 (
            .O(N__8705),
            .I(\b2v_inst.g0_10_a3_7 ));
    CascadeMux I__835 (
            .O(N__8702),
            .I(N__8699));
    InMux I__834 (
            .O(N__8699),
            .I(N__8696));
    LocalMux I__833 (
            .O(N__8696),
            .I(\b2v_inst.reg_ancho_1_i_4 ));
    CascadeMux I__832 (
            .O(N__8693),
            .I(N__8690));
    InMux I__831 (
            .O(N__8690),
            .I(N__8687));
    LocalMux I__830 (
            .O(N__8687),
            .I(\b2v_inst.reg_ancho_1_i_5 ));
    CascadeMux I__829 (
            .O(N__8684),
            .I(N__8681));
    InMux I__828 (
            .O(N__8681),
            .I(N__8678));
    LocalMux I__827 (
            .O(N__8678),
            .I(\b2v_inst.reg_ancho_1_i_6 ));
    CascadeMux I__826 (
            .O(N__8675),
            .I(N__8672));
    InMux I__825 (
            .O(N__8672),
            .I(N__8669));
    LocalMux I__824 (
            .O(N__8669),
            .I(\b2v_inst.reg_ancho_1_i_7 ));
    InMux I__823 (
            .O(N__8666),
            .I(bfn_1_18_0_));
    CascadeMux I__822 (
            .O(N__8663),
            .I(N__8659));
    InMux I__821 (
            .O(N__8662),
            .I(N__8656));
    InMux I__820 (
            .O(N__8659),
            .I(N__8653));
    LocalMux I__819 (
            .O(N__8656),
            .I(\b2v_inst.eventosZ0Z_3 ));
    LocalMux I__818 (
            .O(N__8653),
            .I(\b2v_inst.eventosZ0Z_3 ));
    InMux I__817 (
            .O(N__8648),
            .I(N__8644));
    InMux I__816 (
            .O(N__8647),
            .I(N__8641));
    LocalMux I__815 (
            .O(N__8644),
            .I(\b2v_inst.eventosZ0Z_4 ));
    LocalMux I__814 (
            .O(N__8641),
            .I(\b2v_inst.eventosZ0Z_4 ));
    InMux I__813 (
            .O(N__8636),
            .I(N__8632));
    InMux I__812 (
            .O(N__8635),
            .I(N__8629));
    LocalMux I__811 (
            .O(N__8632),
            .I(\b2v_inst.eventosZ0Z_0 ));
    LocalMux I__810 (
            .O(N__8629),
            .I(\b2v_inst.eventosZ0Z_0 ));
    InMux I__809 (
            .O(N__8624),
            .I(N__8620));
    InMux I__808 (
            .O(N__8623),
            .I(N__8617));
    LocalMux I__807 (
            .O(N__8620),
            .I(\b2v_inst.eventosZ0Z_5 ));
    LocalMux I__806 (
            .O(N__8617),
            .I(\b2v_inst.eventosZ0Z_5 ));
    CEMux I__805 (
            .O(N__8612),
            .I(N__8609));
    LocalMux I__804 (
            .O(N__8609),
            .I(N__8606));
    Odrv4 I__803 (
            .O(N__8606),
            .I(\b2v_inst.N_47_i ));
    CascadeMux I__802 (
            .O(N__8603),
            .I(N__8600));
    InMux I__801 (
            .O(N__8600),
            .I(N__8597));
    LocalMux I__800 (
            .O(N__8597),
            .I(\b2v_inst.reg_ancho_1_i_0 ));
    CascadeMux I__799 (
            .O(N__8594),
            .I(N__8591));
    InMux I__798 (
            .O(N__8591),
            .I(N__8588));
    LocalMux I__797 (
            .O(N__8588),
            .I(\b2v_inst.reg_ancho_1_i_1 ));
    CascadeMux I__796 (
            .O(N__8585),
            .I(N__8582));
    InMux I__795 (
            .O(N__8582),
            .I(N__8579));
    LocalMux I__794 (
            .O(N__8579),
            .I(\b2v_inst.reg_ancho_1_i_2 ));
    CascadeMux I__793 (
            .O(N__8576),
            .I(N__8573));
    InMux I__792 (
            .O(N__8573),
            .I(N__8570));
    LocalMux I__791 (
            .O(N__8570),
            .I(N__8567));
    Odrv4 I__790 (
            .O(N__8567),
            .I(\b2v_inst.reg_ancho_1_i_3 ));
    InMux I__789 (
            .O(N__8564),
            .I(\b2v_inst.eventos_cry_0 ));
    InMux I__788 (
            .O(N__8561),
            .I(\b2v_inst.eventos_cry_1 ));
    InMux I__787 (
            .O(N__8558),
            .I(\b2v_inst.eventos_cry_2 ));
    InMux I__786 (
            .O(N__8555),
            .I(\b2v_inst.eventos_cry_3 ));
    InMux I__785 (
            .O(N__8552),
            .I(\b2v_inst.eventos_cry_4 ));
    InMux I__784 (
            .O(N__8549),
            .I(\b2v_inst.eventos_cry_5 ));
    InMux I__783 (
            .O(N__8546),
            .I(\b2v_inst.eventos_cry_6 ));
    CascadeMux I__782 (
            .O(N__8543),
            .I(N__8539));
    CascadeMux I__781 (
            .O(N__8542),
            .I(N__8536));
    InMux I__780 (
            .O(N__8539),
            .I(N__8526));
    InMux I__779 (
            .O(N__8536),
            .I(N__8526));
    InMux I__778 (
            .O(N__8535),
            .I(N__8526));
    InMux I__777 (
            .O(N__8534),
            .I(N__8521));
    InMux I__776 (
            .O(N__8533),
            .I(N__8521));
    LocalMux I__775 (
            .O(N__8526),
            .I(\b2v_inst.cuenta_pixelZ0Z_7 ));
    LocalMux I__774 (
            .O(N__8521),
            .I(\b2v_inst.cuenta_pixelZ0Z_7 ));
    InMux I__773 (
            .O(N__8516),
            .I(N__8513));
    LocalMux I__772 (
            .O(N__8513),
            .I(N__8505));
    InMux I__771 (
            .O(N__8512),
            .I(N__8496));
    InMux I__770 (
            .O(N__8511),
            .I(N__8496));
    InMux I__769 (
            .O(N__8510),
            .I(N__8496));
    InMux I__768 (
            .O(N__8509),
            .I(N__8496));
    InMux I__767 (
            .O(N__8508),
            .I(N__8493));
    Odrv4 I__766 (
            .O(N__8505),
            .I(\b2v_inst.cuenta_pixelZ0Z_2 ));
    LocalMux I__765 (
            .O(N__8496),
            .I(\b2v_inst.cuenta_pixelZ0Z_2 ));
    LocalMux I__764 (
            .O(N__8493),
            .I(\b2v_inst.cuenta_pixelZ0Z_2 ));
    InMux I__763 (
            .O(N__8486),
            .I(N__8483));
    LocalMux I__762 (
            .O(N__8483),
            .I(\b2v_inst.N_6_i ));
    CascadeMux I__761 (
            .O(N__8480),
            .I(\b2v_inst.g0_6_1_cascade_ ));
    InMux I__760 (
            .O(N__8477),
            .I(N__8474));
    LocalMux I__759 (
            .O(N__8474),
            .I(N__8471));
    Odrv4 I__758 (
            .O(N__8471),
            .I(\b2v_inst.N_4 ));
    CascadeMux I__757 (
            .O(N__8468),
            .I(\b2v_inst.un11_cuenta_pixel_6_cascade_ ));
    InMux I__756 (
            .O(N__8465),
            .I(N__8462));
    LocalMux I__755 (
            .O(N__8462),
            .I(N__8457));
    InMux I__754 (
            .O(N__8461),
            .I(N__8452));
    InMux I__753 (
            .O(N__8460),
            .I(N__8452));
    Odrv4 I__752 (
            .O(N__8457),
            .I(\b2v_inst.un11_cuenta_pixel_6 ));
    LocalMux I__751 (
            .O(N__8452),
            .I(\b2v_inst.un11_cuenta_pixel_6 ));
    InMux I__750 (
            .O(N__8447),
            .I(N__8441));
    InMux I__749 (
            .O(N__8446),
            .I(N__8436));
    InMux I__748 (
            .O(N__8445),
            .I(N__8436));
    InMux I__747 (
            .O(N__8444),
            .I(N__8433));
    LocalMux I__746 (
            .O(N__8441),
            .I(\b2v_inst.cuenta_pixel_RNI3FD32_0Z0Z_5 ));
    LocalMux I__745 (
            .O(N__8436),
            .I(\b2v_inst.cuenta_pixel_RNI3FD32_0Z0Z_5 ));
    LocalMux I__744 (
            .O(N__8433),
            .I(\b2v_inst.cuenta_pixel_RNI3FD32_0Z0Z_5 ));
    InMux I__743 (
            .O(N__8426),
            .I(N__8420));
    InMux I__742 (
            .O(N__8425),
            .I(N__8415));
    InMux I__741 (
            .O(N__8424),
            .I(N__8415));
    InMux I__740 (
            .O(N__8423),
            .I(N__8408));
    LocalMux I__739 (
            .O(N__8420),
            .I(N__8403));
    LocalMux I__738 (
            .O(N__8415),
            .I(N__8403));
    InMux I__737 (
            .O(N__8414),
            .I(N__8394));
    InMux I__736 (
            .O(N__8413),
            .I(N__8394));
    InMux I__735 (
            .O(N__8412),
            .I(N__8394));
    InMux I__734 (
            .O(N__8411),
            .I(N__8394));
    LocalMux I__733 (
            .O(N__8408),
            .I(\b2v_inst.cuenta_pixelZ0Z_3 ));
    Odrv4 I__732 (
            .O(N__8403),
            .I(\b2v_inst.cuenta_pixelZ0Z_3 ));
    LocalMux I__731 (
            .O(N__8394),
            .I(\b2v_inst.cuenta_pixelZ0Z_3 ));
    InMux I__730 (
            .O(N__8387),
            .I(N__8383));
    InMux I__729 (
            .O(N__8386),
            .I(N__8380));
    LocalMux I__728 (
            .O(N__8383),
            .I(N__8373));
    LocalMux I__727 (
            .O(N__8380),
            .I(N__8373));
    InMux I__726 (
            .O(N__8379),
            .I(N__8368));
    InMux I__725 (
            .O(N__8378),
            .I(N__8368));
    Odrv4 I__724 (
            .O(N__8373),
            .I(\b2v_inst.un1_cuenta_pixel_c3 ));
    LocalMux I__723 (
            .O(N__8368),
            .I(\b2v_inst.un1_cuenta_pixel_c3 ));
    CascadeMux I__722 (
            .O(N__8363),
            .I(N__8359));
    CascadeMux I__721 (
            .O(N__8362),
            .I(N__8356));
    InMux I__720 (
            .O(N__8359),
            .I(N__8341));
    InMux I__719 (
            .O(N__8356),
            .I(N__8341));
    InMux I__718 (
            .O(N__8355),
            .I(N__8341));
    InMux I__717 (
            .O(N__8354),
            .I(N__8341));
    InMux I__716 (
            .O(N__8353),
            .I(N__8338));
    InMux I__715 (
            .O(N__8352),
            .I(N__8331));
    InMux I__714 (
            .O(N__8351),
            .I(N__8331));
    InMux I__713 (
            .O(N__8350),
            .I(N__8331));
    LocalMux I__712 (
            .O(N__8341),
            .I(N__8328));
    LocalMux I__711 (
            .O(N__8338),
            .I(\b2v_inst.cuenta_pixelZ0Z_4 ));
    LocalMux I__710 (
            .O(N__8331),
            .I(\b2v_inst.cuenta_pixelZ0Z_4 ));
    Odrv4 I__709 (
            .O(N__8328),
            .I(\b2v_inst.cuenta_pixelZ0Z_4 ));
    InMux I__708 (
            .O(N__8321),
            .I(bfn_1_15_0_));
    CascadeMux I__707 (
            .O(N__8318),
            .I(\b2v_inst.g0_10_a3_0_7_cascade_ ));
    InMux I__706 (
            .O(N__8315),
            .I(N__8312));
    LocalMux I__705 (
            .O(N__8312),
            .I(\b2v_inst.g0_10_a3_0_5 ));
    CascadeMux I__704 (
            .O(N__8309),
            .I(\b2v_inst.g0_10_a3_5_cascade_ ));
    InMux I__703 (
            .O(N__8306),
            .I(N__8303));
    LocalMux I__702 (
            .O(N__8303),
            .I(\b2v_inst.g0_10_a3_4 ));
    InMux I__701 (
            .O(N__8300),
            .I(N__8297));
    LocalMux I__700 (
            .O(N__8297),
            .I(\b2v_inst.un1_cuenta_pixel_c6 ));
    CascadeMux I__699 (
            .O(N__8294),
            .I(\b2v_inst.un1_cuenta_pixel_c6_cascade_ ));
    InMux I__698 (
            .O(N__8291),
            .I(N__8288));
    LocalMux I__697 (
            .O(N__8288),
            .I(\b2v_inst.cuenta_pixel_RNO_0Z0Z_1 ));
    InMux I__696 (
            .O(N__8285),
            .I(N__8282));
    LocalMux I__695 (
            .O(N__8282),
            .I(\b2v_inst.g0_10_a3_0_4 ));
    defparam IN_MUX_bfv_2_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_11_0_));
    defparam IN_MUX_bfv_1_19_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_19_0_));
    defparam IN_MUX_bfv_1_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_20_0_ (
            .carryinitin(\b2v_inst.valor_max_final53 ),
            .carryinitout(bfn_1_20_0_));
    defparam IN_MUX_bfv_5_19_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_19_0_));
    defparam IN_MUX_bfv_5_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_20_0_ (
            .carryinitin(\b2v_inst.valor_max_final52 ),
            .carryinitout(bfn_5_20_0_));
    defparam IN_MUX_bfv_6_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_17_0_));
    defparam IN_MUX_bfv_6_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_18_0_ (
            .carryinitin(\b2v_inst.un3_valor_max2 ),
            .carryinitout(bfn_6_18_0_));
    defparam IN_MUX_bfv_10_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_10_0_));
    defparam IN_MUX_bfv_3_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_15_0_));
    defparam IN_MUX_bfv_3_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_16_0_ (
            .carryinitin(\b2v_inst.data_a_escribir10 ),
            .carryinitout(bfn_3_16_0_));
    defparam IN_MUX_bfv_3_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_13_0_));
    defparam IN_MUX_bfv_3_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_14_0_ (
            .carryinitin(\b2v_inst4.un1_pix_count_int_cry_7 ),
            .carryinitout(bfn_3_14_0_));
    defparam IN_MUX_bfv_1_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_15_0_));
    defparam IN_MUX_bfv_3_19_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_19_0_));
    defparam IN_MUX_bfv_3_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_20_0_ (
            .carryinitin(\b2v_inst.valor_max_final51 ),
            .carryinitout(bfn_3_20_0_));
    defparam IN_MUX_bfv_5_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_17_0_));
    defparam IN_MUX_bfv_5_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_18_0_ (
            .carryinitin(\b2v_inst.valor_max_final50 ),
            .carryinitout(bfn_5_18_0_));
    defparam IN_MUX_bfv_1_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_17_0_));
    defparam IN_MUX_bfv_1_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_18_0_ (
            .carryinitin(\b2v_inst.un3_valor_max1 ),
            .carryinitout(bfn_1_18_0_));
    ICE_GB reset_i_g_gb (
            .USERSIGNALTOGLOBALBUFFER(N__13151),
            .GLOBALBUFFEROUTPUT(reset_i_g));
    ICE_GB \b2v_inst.un1_pix_count_anterior_0_I_39_c_RNIT6R7_0  (
            .USERSIGNALTOGLOBALBUFFER(N__9116),
            .GLOBALBUFFEROUTPUT(\b2v_inst.N_254_i_g ));
    ICE_GB \b2v_inst.state_RNI0PU5_2  (
            .USERSIGNALTOGLOBALBUFFER(N__10171),
            .GLOBALBUFFEROUTPUT(\b2v_inst.state_g_2 ));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \b2v_inst.cuenta_pixel_1_LC_1_11_0 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_pixel_1_LC_1_11_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.cuenta_pixel_1_LC_1_11_0 .LUT_INIT=16'b1010001010101010;
    LogicCell40 \b2v_inst.cuenta_pixel_1_LC_1_11_0  (
            .in0(N__8291),
            .in1(N__8465),
            .in2(N__11801),
            .in3(N__8447),
            .lcout(\b2v_inst.cuenta_pixelZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22410),
            .ce(N__9336),
            .sr(N__22875));
    defparam \b2v_inst.ignorar_ancho_1_RNO_1_LC_1_11_1 .C_ON=1'b0;
    defparam \b2v_inst.ignorar_ancho_1_RNO_1_LC_1_11_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.ignorar_ancho_1_RNO_1_LC_1_11_1 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \b2v_inst.ignorar_ancho_1_RNO_1_LC_1_11_1  (
            .in0(N__8509),
            .in1(N__12422),
            .in2(N__11846),
            .in3(N__12493),
            .lcout(\b2v_inst.g0_10_a3_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.cuenta_pixel_2_LC_1_11_2 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_pixel_2_LC_1_11_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.cuenta_pixel_2_LC_1_11_2 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \b2v_inst.cuenta_pixel_2_LC_1_11_2  (
            .in0(N__12497),
            .in1(_gnd_net_),
            .in2(N__12438),
            .in3(N__8511),
            .lcout(\b2v_inst.cuenta_pixelZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22410),
            .ce(N__9336),
            .sr(N__22875));
    defparam \b2v_inst.cuenta_pixel_RNITIM11_2_LC_1_11_4 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_pixel_RNITIM11_2_LC_1_11_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.cuenta_pixel_RNITIM11_2_LC_1_11_4 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \b2v_inst.cuenta_pixel_RNITIM11_2_LC_1_11_4  (
            .in0(N__12494),
            .in1(_gnd_net_),
            .in2(N__12437),
            .in3(N__8510),
            .lcout(\b2v_inst.un1_cuenta_pixel_c3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.cuenta_pixel_RNIT0FM_1_LC_1_11_5 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_pixel_RNIT0FM_1_LC_1_11_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.cuenta_pixel_RNIT0FM_1_LC_1_11_5 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \b2v_inst.cuenta_pixel_RNIT0FM_1_LC_1_11_5  (
            .in0(_gnd_net_),
            .in1(N__12426),
            .in2(_gnd_net_),
            .in3(N__12495),
            .lcout(\b2v_inst.N_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.cuenta_pixel_3_LC_1_11_6 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_pixel_3_LC_1_11_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.cuenta_pixel_3_LC_1_11_6 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \b2v_inst.cuenta_pixel_3_LC_1_11_6  (
            .in0(N__12498),
            .in1(N__8423),
            .in2(N__12439),
            .in3(N__8512),
            .lcout(\b2v_inst.cuenta_pixelZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22410),
            .ce(N__9336),
            .sr(N__22875));
    defparam \b2v_inst.cuenta_pixel_RNO_0_1_LC_1_11_7 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_pixel_RNO_0_1_LC_1_11_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.cuenta_pixel_RNO_0_1_LC_1_11_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \b2v_inst.cuenta_pixel_RNO_0_1_LC_1_11_7  (
            .in0(_gnd_net_),
            .in1(N__12427),
            .in2(_gnd_net_),
            .in3(N__12496),
            .lcout(\b2v_inst.cuenta_pixel_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.ignorar_ancho_1_RNO_0_LC_1_12_0 .C_ON=1'b0;
    defparam \b2v_inst.ignorar_ancho_1_RNO_0_LC_1_12_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.ignorar_ancho_1_RNO_0_LC_1_12_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \b2v_inst.ignorar_ancho_1_RNO_0_LC_1_12_0  (
            .in0(N__8315),
            .in1(N__8285),
            .in2(_gnd_net_),
            .in3(N__10210),
            .lcout(),
            .ltout(\b2v_inst.g0_10_a3_0_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.ignorar_ancho_1_RNO_LC_1_12_1 .C_ON=1'b0;
    defparam \b2v_inst.ignorar_ancho_1_RNO_LC_1_12_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.ignorar_ancho_1_RNO_LC_1_12_1 .LUT_INIT=16'b1111010001000100;
    LogicCell40 \b2v_inst.ignorar_ancho_1_RNO_LC_1_12_1  (
            .in0(N__15677),
            .in1(N__10164),
            .in2(N__8318),
            .in3(N__8444),
            .lcout(\b2v_inst.un1_state_17_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.cuenta_pixel_RNI3FD32_0_5_LC_1_12_2 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_pixel_RNI3FD32_0_5_LC_1_12_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.cuenta_pixel_RNI3FD32_0_5_LC_1_12_2 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \b2v_inst.cuenta_pixel_RNI3FD32_0_5_LC_1_12_2  (
            .in0(N__8413),
            .in1(N__11759),
            .in2(N__8362),
            .in3(N__8378),
            .lcout(\b2v_inst.cuenta_pixel_RNI3FD32_0Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.ignorar_ancho_1_RNO_2_LC_1_12_3 .C_ON=1'b0;
    defparam \b2v_inst.ignorar_ancho_1_RNO_2_LC_1_12_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.ignorar_ancho_1_RNO_2_LC_1_12_3 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \b2v_inst.ignorar_ancho_1_RNO_2_LC_1_12_3  (
            .in0(N__8533),
            .in1(N__8354),
            .in2(N__15685),
            .in3(N__8411),
            .lcout(\b2v_inst.g0_10_a3_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.ignorar_anterior_RNO_0_LC_1_12_4 .C_ON=1'b0;
    defparam \b2v_inst.ignorar_anterior_RNO_0_LC_1_12_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.ignorar_anterior_RNO_0_LC_1_12_4 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \b2v_inst.ignorar_anterior_RNO_0_LC_1_12_4  (
            .in0(N__8414),
            .in1(N__11760),
            .in2(N__8363),
            .in3(N__8379),
            .lcout(\b2v_inst.g0_10_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.ignorar_anterior_RNO_3_LC_1_12_5 .C_ON=1'b0;
    defparam \b2v_inst.ignorar_anterior_RNO_3_LC_1_12_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.ignorar_anterior_RNO_3_LC_1_12_5 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \b2v_inst.ignorar_anterior_RNO_3_LC_1_12_5  (
            .in0(N__8534),
            .in1(N__8355),
            .in2(N__15686),
            .in3(N__8412),
            .lcout(),
            .ltout(\b2v_inst.g0_10_a3_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.ignorar_anterior_RNO_1_LC_1_12_6 .C_ON=1'b0;
    defparam \b2v_inst.ignorar_anterior_RNO_1_LC_1_12_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.ignorar_anterior_RNO_1_LC_1_12_6 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \b2v_inst.ignorar_anterior_RNO_1_LC_1_12_6  (
            .in0(_gnd_net_),
            .in1(N__8306),
            .in2(N__8309),
            .in3(N__10209),
            .lcout(\b2v_inst.g0_10_a3_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.ignorar_anterior_RNO_2_LC_1_12_7 .C_ON=1'b0;
    defparam \b2v_inst.ignorar_anterior_RNO_2_LC_1_12_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.ignorar_anterior_RNO_2_LC_1_12_7 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \b2v_inst.ignorar_anterior_RNO_2_LC_1_12_7  (
            .in0(N__8508),
            .in1(N__12421),
            .in2(N__11845),
            .in3(N__12473),
            .lcout(\b2v_inst.g0_10_a3_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.cuenta_pixel_7_LC_1_13_0 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_pixel_7_LC_1_13_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.cuenta_pixel_7_LC_1_13_0 .LUT_INIT=16'b0101101011110000;
    LogicCell40 \b2v_inst.cuenta_pixel_7_LC_1_13_0  (
            .in0(N__11834),
            .in1(_gnd_net_),
            .in2(N__8543),
            .in3(N__8300),
            .lcout(\b2v_inst.cuenta_pixelZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22562),
            .ce(N__9337),
            .sr(N__22876));
    defparam \b2v_inst.cuenta_pixel_RNI3FD32_5_LC_1_13_1 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_pixel_RNI3FD32_5_LC_1_13_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.cuenta_pixel_RNI3FD32_5_LC_1_13_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst.cuenta_pixel_RNI3FD32_5_LC_1_13_1  (
            .in0(N__8351),
            .in1(N__8386),
            .in2(N__11764),
            .in3(N__8425),
            .lcout(\b2v_inst.un1_cuenta_pixel_c6 ),
            .ltout(\b2v_inst.un1_cuenta_pixel_c6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.cuenta_pixel_6_LC_1_13_2 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_pixel_6_LC_1_13_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.cuenta_pixel_6_LC_1_13_2 .LUT_INIT=16'b0001001001011010;
    LogicCell40 \b2v_inst.cuenta_pixel_6_LC_1_13_2  (
            .in0(N__11833),
            .in1(N__12395),
            .in2(N__8294),
            .in3(N__8461),
            .lcout(\b2v_inst.cuenta_pixelZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22562),
            .ce(N__9337),
            .sr(N__22876));
    defparam \b2v_inst.cuenta_pixel_RNIC2N11_5_LC_1_13_3 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_pixel_RNIC2N11_5_LC_1_13_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.cuenta_pixel_RNIC2N11_5_LC_1_13_3 .LUT_INIT=16'b1001100100110011;
    LogicCell40 \b2v_inst.cuenta_pixel_RNIC2N11_5_LC_1_13_3  (
            .in0(N__11755),
            .in1(N__8535),
            .in2(_gnd_net_),
            .in3(N__11832),
            .lcout(\b2v_inst.N_6_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.cuenta_pixel_RNI8GUC1_7_LC_1_13_4 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_pixel_RNI8GUC1_7_LC_1_13_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.cuenta_pixel_RNI8GUC1_7_LC_1_13_4 .LUT_INIT=16'b0100010011001101;
    LogicCell40 \b2v_inst.cuenta_pixel_RNI8GUC1_7_LC_1_13_4  (
            .in0(N__8424),
            .in1(N__8350),
            .in2(N__8542),
            .in3(N__8516),
            .lcout(),
            .ltout(\b2v_inst.g0_6_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.cuenta_pixel_RNIJ7CG3_4_LC_1_13_5 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_pixel_RNIJ7CG3_4_LC_1_13_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.cuenta_pixel_RNIJ7CG3_4_LC_1_13_5 .LUT_INIT=16'b0101000000001000;
    LogicCell40 \b2v_inst.cuenta_pixel_RNIJ7CG3_4_LC_1_13_5  (
            .in0(N__8352),
            .in1(N__8486),
            .in2(N__8480),
            .in3(N__8477),
            .lcout(\b2v_inst.un11_cuenta_pixel_6 ),
            .ltout(\b2v_inst.un11_cuenta_pixel_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.cuenta_pixel_5_LC_1_13_6 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_pixel_5_LC_1_13_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.cuenta_pixel_5_LC_1_13_6 .LUT_INIT=16'b1010101000001010;
    LogicCell40 \b2v_inst.cuenta_pixel_5_LC_1_13_6  (
            .in0(N__8446),
            .in1(_gnd_net_),
            .in2(N__8468),
            .in3(N__11787),
            .lcout(\b2v_inst.cuenta_pixelZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22562),
            .ce(N__9337),
            .sr(N__22876));
    defparam \b2v_inst.cuenta_pixel_0_LC_1_13_7 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_pixel_0_LC_1_13_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.cuenta_pixel_0_LC_1_13_7 .LUT_INIT=16'b0000100011111111;
    LogicCell40 \b2v_inst.cuenta_pixel_0_LC_1_13_7  (
            .in0(N__8460),
            .in1(N__8445),
            .in2(N__11794),
            .in3(N__12492),
            .lcout(\b2v_inst.cuenta_pixelZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22562),
            .ce(N__9337),
            .sr(N__22876));
    defparam \b2v_inst.cuenta_pixel_4_LC_1_14_0 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_pixel_4_LC_1_14_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.cuenta_pixel_4_LC_1_14_0 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \b2v_inst.cuenta_pixel_4_LC_1_14_0  (
            .in0(N__8353),
            .in1(N__8426),
            .in2(_gnd_net_),
            .in3(N__8387),
            .lcout(\b2v_inst.cuenta_pixelZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22598),
            .ce(N__9339),
            .sr(N__22879));
    defparam \b2v_inst.pix_count_anterior_12_LC_1_14_1 .C_ON=1'b0;
    defparam \b2v_inst.pix_count_anterior_12_LC_1_14_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.pix_count_anterior_12_LC_1_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.pix_count_anterior_12_LC_1_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9397),
            .lcout(\b2v_inst.pix_count_anteriorZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22598),
            .ce(N__9339),
            .sr(N__22879));
    defparam \b2v_inst.eventos_0_LC_1_15_0 .C_ON=1'b1;
    defparam \b2v_inst.eventos_0_LC_1_15_0 .SEQ_MODE=4'b1011;
    defparam \b2v_inst.eventos_0_LC_1_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.eventos_0_LC_1_15_0  (
            .in0(_gnd_net_),
            .in1(N__8635),
            .in2(_gnd_net_),
            .in3(N__8321),
            .lcout(\b2v_inst.eventosZ0Z_0 ),
            .ltout(),
            .carryin(bfn_1_15_0_),
            .carryout(\b2v_inst.eventos_cry_0 ),
            .clk(N__22509),
            .ce(N__8612),
            .sr(N__22882));
    defparam \b2v_inst.eventos_1_LC_1_15_1 .C_ON=1'b1;
    defparam \b2v_inst.eventos_1_LC_1_15_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.eventos_1_LC_1_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.eventos_1_LC_1_15_1  (
            .in0(_gnd_net_),
            .in1(N__9604),
            .in2(_gnd_net_),
            .in3(N__8564),
            .lcout(\b2v_inst.eventosZ0Z_1 ),
            .ltout(),
            .carryin(\b2v_inst.eventos_cry_0 ),
            .carryout(\b2v_inst.eventos_cry_1 ),
            .clk(N__22509),
            .ce(N__8612),
            .sr(N__22882));
    defparam \b2v_inst.eventos_2_LC_1_15_2 .C_ON=1'b1;
    defparam \b2v_inst.eventos_2_LC_1_15_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.eventos_2_LC_1_15_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.eventos_2_LC_1_15_2  (
            .in0(_gnd_net_),
            .in1(N__8959),
            .in2(_gnd_net_),
            .in3(N__8561),
            .lcout(\b2v_inst.eventosZ0Z_2 ),
            .ltout(),
            .carryin(\b2v_inst.eventos_cry_1 ),
            .carryout(\b2v_inst.eventos_cry_2 ),
            .clk(N__22509),
            .ce(N__8612),
            .sr(N__22882));
    defparam \b2v_inst.eventos_3_LC_1_15_3 .C_ON=1'b1;
    defparam \b2v_inst.eventos_3_LC_1_15_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.eventos_3_LC_1_15_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.eventos_3_LC_1_15_3  (
            .in0(_gnd_net_),
            .in1(N__8662),
            .in2(_gnd_net_),
            .in3(N__8558),
            .lcout(\b2v_inst.eventosZ0Z_3 ),
            .ltout(),
            .carryin(\b2v_inst.eventos_cry_2 ),
            .carryout(\b2v_inst.eventos_cry_3 ),
            .clk(N__22509),
            .ce(N__8612),
            .sr(N__22882));
    defparam \b2v_inst.eventos_4_LC_1_15_4 .C_ON=1'b1;
    defparam \b2v_inst.eventos_4_LC_1_15_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.eventos_4_LC_1_15_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.eventos_4_LC_1_15_4  (
            .in0(_gnd_net_),
            .in1(N__8647),
            .in2(_gnd_net_),
            .in3(N__8555),
            .lcout(\b2v_inst.eventosZ0Z_4 ),
            .ltout(),
            .carryin(\b2v_inst.eventos_cry_3 ),
            .carryout(\b2v_inst.eventos_cry_4 ),
            .clk(N__22509),
            .ce(N__8612),
            .sr(N__22882));
    defparam \b2v_inst.eventos_5_LC_1_15_5 .C_ON=1'b1;
    defparam \b2v_inst.eventos_5_LC_1_15_5 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.eventos_5_LC_1_15_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.eventos_5_LC_1_15_5  (
            .in0(_gnd_net_),
            .in1(N__8624),
            .in2(_gnd_net_),
            .in3(N__8552),
            .lcout(\b2v_inst.eventosZ0Z_5 ),
            .ltout(),
            .carryin(\b2v_inst.eventos_cry_4 ),
            .carryout(\b2v_inst.eventos_cry_5 ),
            .clk(N__22509),
            .ce(N__8612),
            .sr(N__22882));
    defparam \b2v_inst.eventos_6_LC_1_15_6 .C_ON=1'b1;
    defparam \b2v_inst.eventos_6_LC_1_15_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.eventos_6_LC_1_15_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst.eventos_6_LC_1_15_6  (
            .in0(_gnd_net_),
            .in1(N__9589),
            .in2(_gnd_net_),
            .in3(N__8549),
            .lcout(\b2v_inst.eventosZ0Z_6 ),
            .ltout(),
            .carryin(\b2v_inst.eventos_cry_5 ),
            .carryout(\b2v_inst.eventos_cry_6 ),
            .clk(N__22509),
            .ce(N__8612),
            .sr(N__22882));
    defparam \b2v_inst.eventos_7_LC_1_15_7 .C_ON=1'b0;
    defparam \b2v_inst.eventos_7_LC_1_15_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.eventos_7_LC_1_15_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \b2v_inst.eventos_7_LC_1_15_7  (
            .in0(_gnd_net_),
            .in1(N__9526),
            .in2(_gnd_net_),
            .in3(N__8546),
            .lcout(\b2v_inst.eventosZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22509),
            .ce(N__8612),
            .sr(N__22882));
    defparam \b2v_inst.data_a_escribir_RNO_1_7_LC_1_16_0 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_1_7_LC_1_16_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_1_7_LC_1_16_0 .LUT_INIT=16'b0000001000010011;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_1_7_LC_1_16_0  (
            .in0(N__10695),
            .in1(N__10543),
            .in2(N__11222),
            .in3(N__10793),
            .lcout(\b2v_inst.un1_reg_anterior_iv_0_0_2_0_tz_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.reg_ancho_1_7_LC_1_16_1 .C_ON=1'b0;
    defparam \b2v_inst.reg_ancho_1_7_LC_1_16_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_ancho_1_7_LC_1_16_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \b2v_inst.reg_ancho_1_7_LC_1_16_1  (
            .in0(_gnd_net_),
            .in1(N__8885),
            .in2(_gnd_net_),
            .in3(N__13638),
            .lcout(\b2v_inst.reg_ancho_1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22570),
            .ce(N__13913),
            .sr(N__22886));
    defparam \b2v_inst.reg_ancho_1_6_LC_1_16_2 .C_ON=1'b0;
    defparam \b2v_inst.reg_ancho_1_6_LC_1_16_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_ancho_1_6_LC_1_16_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \b2v_inst.reg_ancho_1_6_LC_1_16_2  (
            .in0(N__8884),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14241),
            .lcout(\b2v_inst.reg_ancho_1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22570),
            .ce(N__13913),
            .sr(N__22886));
    defparam \b2v_inst.data_a_escribir_RNO_4_3_LC_1_16_3 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_4_3_LC_1_16_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_4_3_LC_1_16_3 .LUT_INIT=16'b0000101000011011;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_4_3_LC_1_16_3  (
            .in0(N__10542),
            .in1(N__11021),
            .in2(N__8663),
            .in3(N__10696),
            .lcout(\b2v_inst.un1_reg_anterior_iv_0_0_1_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_1_4_LC_1_16_4 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_1_4_LC_1_16_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_1_4_LC_1_16_4 .LUT_INIT=16'b0111011101010101;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_1_4_LC_1_16_4  (
            .in0(N__14795),
            .in1(N__8648),
            .in2(_gnd_net_),
            .in3(N__10547),
            .lcout(\b2v_inst.un1_reg_anterior_iv_0_0_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_2_0_LC_1_16_5 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_2_0_LC_1_16_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_2_0_LC_1_16_5 .LUT_INIT=16'b0010001011111111;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_2_0_LC_1_16_5  (
            .in0(N__10545),
            .in1(N__8636),
            .in2(_gnd_net_),
            .in3(N__14793),
            .lcout(\b2v_inst.un1_reg_anterior_iv_0_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_2_5_LC_1_16_6 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_2_5_LC_1_16_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_2_5_LC_1_16_6 .LUT_INIT=16'b0111011101010101;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_2_5_LC_1_16_6  (
            .in0(N__14794),
            .in1(N__8623),
            .in2(_gnd_net_),
            .in3(N__10546),
            .lcout(\b2v_inst.un1_reg_anterior_iv_0_0_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNIN3GK_7_LC_1_16_7 .C_ON=1'b0;
    defparam \b2v_inst.state_RNIN3GK_7_LC_1_16_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNIN3GK_7_LC_1_16_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \b2v_inst.state_RNIN3GK_7_LC_1_16_7  (
            .in0(N__10544),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14792),
            .lcout(\b2v_inst.N_47_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_un3_valor_max1_cry_0_c_inv_LC_1_17_0 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_un3_valor_max1_cry_0_c_inv_LC_1_17_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_un3_valor_max1_cry_0_c_inv_LC_1_17_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst.encontrar_maximo_un3_valor_max1_cry_0_c_inv_LC_1_17_0  (
            .in0(N__10286),
            .in1(N__11511),
            .in2(N__8603),
            .in3(_gnd_net_),
            .lcout(\b2v_inst.reg_ancho_1_i_0 ),
            .ltout(),
            .carryin(bfn_1_17_0_),
            .carryout(\b2v_inst.un3_valor_max1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_un3_valor_max1_cry_1_c_inv_LC_1_17_1 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_un3_valor_max1_cry_1_c_inv_LC_1_17_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_un3_valor_max1_cry_1_c_inv_LC_1_17_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst.encontrar_maximo_un3_valor_max1_cry_1_c_inv_LC_1_17_1  (
            .in0(_gnd_net_),
            .in1(N__11473),
            .in2(N__8594),
            .in3(N__11155),
            .lcout(\b2v_inst.reg_ancho_1_i_1 ),
            .ltout(),
            .carryin(\b2v_inst.un3_valor_max1_cry_0 ),
            .carryout(\b2v_inst.un3_valor_max1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_un3_valor_max1_cry_2_c_inv_LC_1_17_2 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_un3_valor_max1_cry_2_c_inv_LC_1_17_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_un3_valor_max1_cry_2_c_inv_LC_1_17_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst.encontrar_maximo_un3_valor_max1_cry_2_c_inv_LC_1_17_2  (
            .in0(_gnd_net_),
            .in1(N__11427),
            .in2(N__8585),
            .in3(N__11056),
            .lcout(\b2v_inst.reg_ancho_1_i_2 ),
            .ltout(),
            .carryin(\b2v_inst.un3_valor_max1_cry_1 ),
            .carryout(\b2v_inst.un3_valor_max1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_un3_valor_max1_cry_3_c_inv_LC_1_17_3 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_un3_valor_max1_cry_3_c_inv_LC_1_17_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_un3_valor_max1_cry_3_c_inv_LC_1_17_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst.encontrar_maximo_un3_valor_max1_cry_3_c_inv_LC_1_17_3  (
            .in0(_gnd_net_),
            .in1(N__11386),
            .in2(N__8576),
            .in3(N__11011),
            .lcout(\b2v_inst.reg_ancho_1_i_3 ),
            .ltout(),
            .carryin(\b2v_inst.un3_valor_max1_cry_2 ),
            .carryout(\b2v_inst.un3_valor_max1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_un3_valor_max1_cry_4_c_inv_LC_1_17_4 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_un3_valor_max1_cry_4_c_inv_LC_1_17_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_un3_valor_max1_cry_4_c_inv_LC_1_17_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst.encontrar_maximo_un3_valor_max1_cry_4_c_inv_LC_1_17_4  (
            .in0(_gnd_net_),
            .in1(N__11337),
            .in2(N__8702),
            .in3(N__10942),
            .lcout(\b2v_inst.reg_ancho_1_i_4 ),
            .ltout(),
            .carryin(\b2v_inst.un3_valor_max1_cry_3 ),
            .carryout(\b2v_inst.un3_valor_max1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_un3_valor_max1_cry_5_c_inv_LC_1_17_5 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_un3_valor_max1_cry_5_c_inv_LC_1_17_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_un3_valor_max1_cry_5_c_inv_LC_1_17_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst.encontrar_maximo_un3_valor_max1_cry_5_c_inv_LC_1_17_5  (
            .in0(_gnd_net_),
            .in1(N__11304),
            .in2(N__8693),
            .in3(N__10870),
            .lcout(\b2v_inst.reg_ancho_1_i_5 ),
            .ltout(),
            .carryin(\b2v_inst.un3_valor_max1_cry_4 ),
            .carryout(\b2v_inst.un3_valor_max1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_un3_valor_max1_cry_6_c_inv_LC_1_17_6 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_un3_valor_max1_cry_6_c_inv_LC_1_17_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_un3_valor_max1_cry_6_c_inv_LC_1_17_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst.encontrar_maximo_un3_valor_max1_cry_6_c_inv_LC_1_17_6  (
            .in0(_gnd_net_),
            .in1(N__11243),
            .in2(N__8684),
            .in3(N__10828),
            .lcout(\b2v_inst.reg_ancho_1_i_6 ),
            .ltout(),
            .carryin(\b2v_inst.un3_valor_max1_cry_5 ),
            .carryout(\b2v_inst.un3_valor_max1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_un3_valor_max1_cry_7_c_inv_LC_1_17_7 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_un3_valor_max1_cry_7_c_inv_LC_1_17_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_un3_valor_max1_cry_7_c_inv_LC_1_17_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst.encontrar_maximo_un3_valor_max1_cry_7_c_inv_LC_1_17_7  (
            .in0(_gnd_net_),
            .in1(N__11213),
            .in2(N__8675),
            .in3(N__10783),
            .lcout(\b2v_inst.reg_ancho_1_i_7 ),
            .ltout(),
            .carryin(\b2v_inst.un3_valor_max1_cry_6 ),
            .carryout(\b2v_inst.un3_valor_max1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un3_valor_max1_THRU_LUT4_0_LC_1_18_0 .C_ON=1'b0;
    defparam \b2v_inst.un3_valor_max1_THRU_LUT4_0_LC_1_18_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un3_valor_max1_THRU_LUT4_0_LC_1_18_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.un3_valor_max1_THRU_LUT4_0_LC_1_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8666),
            .lcout(\b2v_inst.un3_valor_max1_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_0_0_LC_1_18_2 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_0_0_LC_1_18_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_0_0_LC_1_18_2 .LUT_INIT=16'b1111110011111010;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_0_0_LC_1_18_2  (
            .in0(N__10287),
            .in1(N__11510),
            .in2(N__10570),
            .in3(N__10681),
            .lcout(\b2v_inst.un1_m3_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_4_2_LC_1_18_4 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_4_2_LC_1_18_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_4_2_LC_1_18_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_4_2_LC_1_18_4  (
            .in0(_gnd_net_),
            .in1(N__11426),
            .in2(_gnd_net_),
            .in3(N__10680),
            .lcout(\b2v_inst.un1_reg_anterior_iv_0_0_a2_4_tz_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst3.reset_i_LC_1_18_6 .C_ON=1'b0;
    defparam \b2v_inst3.reset_i_LC_1_18_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst3.reset_i_LC_1_18_6 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \b2v_inst3.reset_i_LC_1_18_6  (
            .in0(_gnd_net_),
            .in1(N__18933),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(reset_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_3_cry_0_c_LC_1_19_0 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_3_cry_0_c_LC_1_19_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_3_cry_0_c_LC_1_19_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final5_3_cry_0_c_LC_1_19_0  (
            .in0(_gnd_net_),
            .in1(N__9628),
            .in2(N__11513),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_19_0_),
            .carryout(\b2v_inst.valor_max_final5_3_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_3_cry_1_c_LC_1_19_1 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_3_cry_1_c_LC_1_19_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_3_cry_1_c_LC_1_19_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final5_3_cry_1_c_LC_1_19_1  (
            .in0(_gnd_net_),
            .in1(N__9871),
            .in2(N__11471),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.valor_max_final5_3_cry_0 ),
            .carryout(\b2v_inst.valor_max_final5_3_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_3_cry_2_c_LC_1_19_2 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_3_cry_2_c_LC_1_19_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_3_cry_2_c_LC_1_19_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final5_3_cry_2_c_LC_1_19_2  (
            .in0(_gnd_net_),
            .in1(N__9853),
            .in2(N__11429),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.valor_max_final5_3_cry_1 ),
            .carryout(\b2v_inst.valor_max_final5_3_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_3_cry_3_c_LC_1_19_3 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_3_cry_3_c_LC_1_19_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_3_cry_3_c_LC_1_19_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final5_3_cry_3_c_LC_1_19_3  (
            .in0(_gnd_net_),
            .in1(N__9835),
            .in2(N__11389),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.valor_max_final5_3_cry_2 ),
            .carryout(\b2v_inst.valor_max_final5_3_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_3_cry_4_c_LC_1_19_4 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_3_cry_4_c_LC_1_19_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_3_cry_4_c_LC_1_19_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final5_3_cry_4_c_LC_1_19_4  (
            .in0(_gnd_net_),
            .in1(N__11345),
            .in2(N__9818),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.valor_max_final5_3_cry_3 ),
            .carryout(\b2v_inst.valor_max_final5_3_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_3_cry_5_c_LC_1_19_5 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_3_cry_5_c_LC_1_19_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_3_cry_5_c_LC_1_19_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final5_3_cry_5_c_LC_1_19_5  (
            .in0(_gnd_net_),
            .in1(N__11308),
            .in2(N__9797),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.valor_max_final5_3_cry_4 ),
            .carryout(\b2v_inst.valor_max_final5_3_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_3_cry_6_c_LC_1_19_6 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_3_cry_6_c_LC_1_19_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_3_cry_6_c_LC_1_19_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final5_3_cry_6_c_LC_1_19_6  (
            .in0(_gnd_net_),
            .in1(N__11263),
            .in2(N__9775),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.valor_max_final5_3_cry_5 ),
            .carryout(\b2v_inst.valor_max_final5_3_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_3_cry_7_c_LC_1_19_7 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_3_cry_7_c_LC_1_19_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_3_cry_7_c_LC_1_19_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final5_3_cry_7_c_LC_1_19_7  (
            .in0(_gnd_net_),
            .in1(N__9752),
            .in2(N__11217),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.valor_max_final5_3_cry_6 ),
            .carryout(\b2v_inst.valor_max_final53 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.valor_max_final53_THRU_LUT4_0_LC_1_20_0 .C_ON=1'b0;
    defparam \b2v_inst.valor_max_final53_THRU_LUT4_0_LC_1_20_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.valor_max_final53_THRU_LUT4_0_LC_1_20_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.valor_max_final53_THRU_LUT4_0_LC_1_20_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8729),
            .lcout(\b2v_inst.valor_max_final53_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.ignorar_anterior_RNO_LC_1_20_4 .C_ON=1'b0;
    defparam \b2v_inst.ignorar_anterior_RNO_LC_1_20_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.ignorar_anterior_RNO_LC_1_20_4 .LUT_INIT=16'b1101110001010000;
    LogicCell40 \b2v_inst.ignorar_anterior_RNO_LC_1_20_4  (
            .in0(N__15683),
            .in1(N__8726),
            .in2(N__10172),
            .in3(N__8714),
            .lcout(\b2v_inst.un1_state_19_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un1_pix_count_anterior_0_I_1_c_LC_2_11_0 .C_ON=1'b1;
    defparam \b2v_inst.un1_pix_count_anterior_0_I_1_c_LC_2_11_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un1_pix_count_anterior_0_I_1_c_LC_2_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.un1_pix_count_anterior_0_I_1_c_LC_2_11_0  (
            .in0(_gnd_net_),
            .in1(N__8750),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_11_0_),
            .carryout(\b2v_inst.un1_pix_count_anterior_0_data_tmp_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un1_pix_count_anterior_0_I_27_c_LC_2_11_1 .C_ON=1'b1;
    defparam \b2v_inst.un1_pix_count_anterior_0_I_27_c_LC_2_11_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un1_pix_count_anterior_0_I_27_c_LC_2_11_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.un1_pix_count_anterior_0_I_27_c_LC_2_11_1  (
            .in0(_gnd_net_),
            .in1(N__9101),
            .in2(N__18605),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.un1_pix_count_anterior_0_data_tmp_0 ),
            .carryout(\b2v_inst.un1_pix_count_anterior_0_data_tmp_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un1_pix_count_anterior_0_I_15_c_LC_2_11_2 .C_ON=1'b1;
    defparam \b2v_inst.un1_pix_count_anterior_0_I_15_c_LC_2_11_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un1_pix_count_anterior_0_I_15_c_LC_2_11_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.un1_pix_count_anterior_0_I_15_c_LC_2_11_2  (
            .in0(_gnd_net_),
            .in1(N__8735),
            .in2(N__18601),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.un1_pix_count_anterior_0_data_tmp_1 ),
            .carryout(\b2v_inst.un1_pix_count_anterior_0_data_tmp_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un1_pix_count_anterior_0_I_21_c_LC_2_11_3 .C_ON=1'b1;
    defparam \b2v_inst.un1_pix_count_anterior_0_I_21_c_LC_2_11_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un1_pix_count_anterior_0_I_21_c_LC_2_11_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.un1_pix_count_anterior_0_I_21_c_LC_2_11_3  (
            .in0(_gnd_net_),
            .in1(N__8792),
            .in2(N__18604),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.un1_pix_count_anterior_0_data_tmp_2 ),
            .carryout(\b2v_inst.un1_pix_count_anterior_0_data_tmp_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un1_pix_count_anterior_0_I_51_c_LC_2_11_4 .C_ON=1'b1;
    defparam \b2v_inst.un1_pix_count_anterior_0_I_51_c_LC_2_11_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un1_pix_count_anterior_0_I_51_c_LC_2_11_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.un1_pix_count_anterior_0_I_51_c_LC_2_11_4  (
            .in0(_gnd_net_),
            .in1(N__8837),
            .in2(N__18603),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.un1_pix_count_anterior_0_data_tmp_3 ),
            .carryout(\b2v_inst.un1_pix_count_anterior_0_data_tmp_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un1_pix_count_anterior_0_I_9_c_LC_2_11_5 .C_ON=1'b1;
    defparam \b2v_inst.un1_pix_count_anterior_0_I_9_c_LC_2_11_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un1_pix_count_anterior_0_I_9_c_LC_2_11_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.un1_pix_count_anterior_0_I_9_c_LC_2_11_5  (
            .in0(_gnd_net_),
            .in1(N__9080),
            .in2(N__18606),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.un1_pix_count_anterior_0_data_tmp_4 ),
            .carryout(\b2v_inst.un1_pix_count_anterior_0_data_tmp_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un1_pix_count_anterior_0_I_39_c_LC_2_11_6 .C_ON=1'b1;
    defparam \b2v_inst.un1_pix_count_anterior_0_I_39_c_LC_2_11_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un1_pix_count_anterior_0_I_39_c_LC_2_11_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.un1_pix_count_anterior_0_I_39_c_LC_2_11_6  (
            .in0(_gnd_net_),
            .in1(N__8801),
            .in2(N__18602),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.un1_pix_count_anterior_0_data_tmp_5 ),
            .carryout(\b2v_inst.un1_pix_count_anterior_0_N_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un1_pix_count_anterior_0_N_2_THRU_LUT4_0_LC_2_11_7 .C_ON=1'b0;
    defparam \b2v_inst.un1_pix_count_anterior_0_N_2_THRU_LUT4_0_LC_2_11_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un1_pix_count_anterior_0_N_2_THRU_LUT4_0_LC_2_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.un1_pix_count_anterior_0_N_2_THRU_LUT4_0_LC_2_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8738),
            .lcout(\b2v_inst.un1_pix_count_anterior_0_N_2_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un1_pix_count_anterior_0_I_15_c_RNO_LC_2_12_0 .C_ON=1'b0;
    defparam \b2v_inst.un1_pix_count_anterior_0_I_15_c_RNO_LC_2_12_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un1_pix_count_anterior_0_I_15_c_RNO_LC_2_12_0 .LUT_INIT=16'b0110111111110110;
    LogicCell40 \b2v_inst.un1_pix_count_anterior_0_I_15_c_RNO_LC_2_12_0  (
            .in0(N__9206),
            .in1(N__8774),
            .in2(N__8768),
            .in3(N__9185),
            .lcout(\b2v_inst.un1_pix_count_anterior_0_I_15_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.pix_count_anterior_4_LC_2_12_1 .C_ON=1'b0;
    defparam \b2v_inst.pix_count_anterior_4_LC_2_12_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.pix_count_anterior_4_LC_2_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.pix_count_anterior_4_LC_2_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9208),
            .lcout(\b2v_inst.pix_count_anteriorZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22587),
            .ce(N__9338),
            .sr(N__22877));
    defparam \b2v_inst.pix_count_anterior_5_LC_2_12_2 .C_ON=1'b0;
    defparam \b2v_inst.pix_count_anterior_5_LC_2_12_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.pix_count_anterior_5_LC_2_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.pix_count_anterior_5_LC_2_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9186),
            .lcout(\b2v_inst.pix_count_anteriorZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22587),
            .ce(N__9338),
            .sr(N__22877));
    defparam \b2v_inst4.pix_count_int_RNITN3K1_1_LC_2_12_3 .C_ON=1'b0;
    defparam \b2v_inst4.pix_count_int_RNITN3K1_1_LC_2_12_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst4.pix_count_int_RNITN3K1_1_LC_2_12_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst4.pix_count_int_RNITN3K1_1_LC_2_12_3  (
            .in0(N__9158),
            .in1(N__9282),
            .in2(N__9263),
            .in3(N__9207),
            .lcout(\b2v_inst4.un1_pix_count_int_0_sqmuxa_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.pix_count_anterior_1_LC_2_12_4 .C_ON=1'b0;
    defparam \b2v_inst.pix_count_anterior_1_LC_2_12_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.pix_count_anterior_1_LC_2_12_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst.pix_count_anterior_1_LC_2_12_4  (
            .in0(N__9283),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst.pix_count_anteriorZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22587),
            .ce(N__9338),
            .sr(N__22877));
    defparam \b2v_inst.un1_pix_count_anterior_0_I_1_c_RNO_LC_2_12_5 .C_ON=1'b0;
    defparam \b2v_inst.un1_pix_count_anterior_0_I_1_c_RNO_LC_2_12_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un1_pix_count_anterior_0_I_1_c_RNO_LC_2_12_5 .LUT_INIT=16'b0110111111110110;
    LogicCell40 \b2v_inst.un1_pix_count_anterior_0_I_1_c_RNO_LC_2_12_5  (
            .in0(N__8744),
            .in1(N__9308),
            .in2(N__8759),
            .in3(N__9281),
            .lcout(\b2v_inst.un1_pix_count_anterior_0_I_1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.pix_count_anterior_0_LC_2_12_6 .C_ON=1'b0;
    defparam \b2v_inst.pix_count_anterior_0_LC_2_12_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.pix_count_anterior_0_LC_2_12_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst.pix_count_anterior_0_LC_2_12_6  (
            .in0(N__9309),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst.pix_count_anteriorZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22587),
            .ce(N__9338),
            .sr(N__22877));
    defparam \b2v_inst.pix_count_anterior_2_LC_2_12_7 .C_ON=1'b0;
    defparam \b2v_inst.pix_count_anterior_2_LC_2_12_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.pix_count_anterior_2_LC_2_12_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst.pix_count_anterior_2_LC_2_12_7  (
            .in0(N__9262),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst.pix_count_anteriorZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22587),
            .ce(N__9338),
            .sr(N__22877));
    defparam \b2v_inst4.pix_count_int_0_LC_2_13_0 .C_ON=1'b0;
    defparam \b2v_inst4.pix_count_int_0_LC_2_13_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst4.pix_count_int_0_LC_2_13_0 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \b2v_inst4.pix_count_int_0_LC_2_13_0  (
            .in0(N__12007),
            .in1(N__11971),
            .in2(N__11944),
            .in3(N__9290),
            .lcout(SYNTHESIZED_WIRE_2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22496),
            .ce(),
            .sr(N__22880));
    defparam \b2v_inst4.pix_count_int_11_LC_2_13_1 .C_ON=1'b0;
    defparam \b2v_inst4.pix_count_int_11_LC_2_13_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst4.pix_count_int_11_LC_2_13_1 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \b2v_inst4.pix_count_int_11_LC_2_13_1  (
            .in0(N__11972),
            .in1(N__12008),
            .in2(N__11923),
            .in3(N__9407),
            .lcout(SYNTHESIZED_WIRE_2_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22496),
            .ce(),
            .sr(N__22880));
    defparam \b2v_inst4.pix_count_int_12_LC_2_13_2 .C_ON=1'b0;
    defparam \b2v_inst4.pix_count_int_12_LC_2_13_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst4.pix_count_int_12_LC_2_13_2 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \b2v_inst4.pix_count_int_12_LC_2_13_2  (
            .in0(N__12009),
            .in1(N__11973),
            .in2(N__11945),
            .in3(N__9368),
            .lcout(SYNTHESIZED_WIRE_2_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22496),
            .ce(),
            .sr(N__22880));
    defparam \b2v_inst.un1_pix_count_anterior_0_I_39_c_RNO_LC_2_13_3 .C_ON=1'b0;
    defparam \b2v_inst.un1_pix_count_anterior_0_I_39_c_RNO_LC_2_13_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un1_pix_count_anterior_0_I_39_c_RNO_LC_2_13_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \b2v_inst.un1_pix_count_anterior_0_I_39_c_RNO_LC_2_13_3  (
            .in0(_gnd_net_),
            .in1(N__8807),
            .in2(_gnd_net_),
            .in3(N__9392),
            .lcout(\b2v_inst.un1_pix_count_anterior_0_I_39_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst4.pix_count_int_3_LC_2_13_4 .C_ON=1'b0;
    defparam \b2v_inst4.pix_count_int_3_LC_2_13_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst4.pix_count_int_3_LC_2_13_4 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \b2v_inst4.pix_count_int_3_LC_2_13_4  (
            .in0(N__12010),
            .in1(N__11974),
            .in2(N__11946),
            .in3(N__9218),
            .lcout(SYNTHESIZED_WIRE_2_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22496),
            .ce(),
            .sr(N__22880));
    defparam \b2v_inst4.pix_count_int_5_LC_2_13_5 .C_ON=1'b0;
    defparam \b2v_inst4.pix_count_int_5_LC_2_13_5 .SEQ_MODE=4'b1010;
    defparam \b2v_inst4.pix_count_int_5_LC_2_13_5 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \b2v_inst4.pix_count_int_5_LC_2_13_5  (
            .in0(N__11975),
            .in1(N__12011),
            .in2(N__11924),
            .in3(N__9167),
            .lcout(SYNTHESIZED_WIRE_2_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22496),
            .ce(),
            .sr(N__22880));
    defparam \b2v_inst4.pix_count_int_7_LC_2_13_6 .C_ON=1'b0;
    defparam \b2v_inst4.pix_count_int_7_LC_2_13_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst4.pix_count_int_7_LC_2_13_6 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \b2v_inst4.pix_count_int_7_LC_2_13_6  (
            .in0(N__12012),
            .in1(N__11976),
            .in2(N__11947),
            .in3(N__9494),
            .lcout(SYNTHESIZED_WIRE_2_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22496),
            .ce(),
            .sr(N__22880));
    defparam \b2v_inst4.pix_count_int_8_LC_2_13_7 .C_ON=1'b0;
    defparam \b2v_inst4.pix_count_int_8_LC_2_13_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst4.pix_count_int_8_LC_2_13_7 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \b2v_inst4.pix_count_int_8_LC_2_13_7  (
            .in0(N__11977),
            .in1(N__12013),
            .in2(N__11925),
            .in3(N__9467),
            .lcout(SYNTHESIZED_WIRE_2_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22496),
            .ce(),
            .sr(N__22880));
    defparam \b2v_inst.un1_pix_count_anterior_0_I_21_c_RNO_LC_2_14_0 .C_ON=1'b0;
    defparam \b2v_inst.un1_pix_count_anterior_0_I_21_c_RNO_LC_2_14_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un1_pix_count_anterior_0_I_21_c_RNO_LC_2_14_0 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \b2v_inst.un1_pix_count_anterior_0_I_21_c_RNO_LC_2_14_0  (
            .in0(N__9509),
            .in1(N__8783),
            .in2(N__8852),
            .in3(N__9155),
            .lcout(\b2v_inst.un1_pix_count_anterior_0_I_21_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.pix_count_anterior_6_LC_2_14_1 .C_ON=1'b0;
    defparam \b2v_inst.pix_count_anterior_6_LC_2_14_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.pix_count_anterior_6_LC_2_14_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst.pix_count_anterior_6_LC_2_14_1  (
            .in0(N__9156),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst.pix_count_anteriorZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22588),
            .ce(N__9341),
            .sr(N__22883));
    defparam \b2v_inst4.pix_count_int_RNI6KOL1_12_LC_2_14_2 .C_ON=1'b0;
    defparam \b2v_inst4.pix_count_int_RNI6KOL1_12_LC_2_14_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst4.pix_count_int_RNI6KOL1_12_LC_2_14_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst4.pix_count_int_RNI6KOL1_12_LC_2_14_2  (
            .in0(N__9428),
            .in1(N__11868),
            .in2(N__9398),
            .in3(N__9483),
            .lcout(),
            .ltout(\b2v_inst4.un1_pix_count_int_0_sqmuxa_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst4.state_RNIC9UM2_0_LC_2_14_3 .C_ON=1'b0;
    defparam \b2v_inst4.state_RNIC9UM2_0_LC_2_14_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst4.state_RNIC9UM2_0_LC_2_14_3 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \b2v_inst4.state_RNIC9UM2_0_LC_2_14_3  (
            .in0(N__11714),
            .in1(N__9510),
            .in2(N__8777),
            .in3(N__9188),
            .lcout(\b2v_inst4.un1_pix_count_int_0_sqmuxa_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.pix_count_anterior_7_LC_2_14_4 .C_ON=1'b0;
    defparam \b2v_inst.pix_count_anterior_7_LC_2_14_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.pix_count_anterior_7_LC_2_14_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst.pix_count_anterior_7_LC_2_14_4  (
            .in0(N__9511),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst.pix_count_anteriorZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22588),
            .ce(N__9341),
            .sr(N__22883));
    defparam \b2v_inst.pix_count_anterior_8_LC_2_14_5 .C_ON=1'b0;
    defparam \b2v_inst.pix_count_anterior_8_LC_2_14_5 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.pix_count_anterior_8_LC_2_14_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst.pix_count_anterior_8_LC_2_14_5  (
            .in0(N__9484),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst.pix_count_anteriorZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22588),
            .ce(N__9341),
            .sr(N__22883));
    defparam \b2v_inst.un1_pix_count_anterior_0_I_51_c_RNO_LC_2_14_6 .C_ON=1'b0;
    defparam \b2v_inst.un1_pix_count_anterior_0_I_51_c_RNO_LC_2_14_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un1_pix_count_anterior_0_I_51_c_RNO_LC_2_14_6 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \b2v_inst.un1_pix_count_anterior_0_I_51_c_RNO_LC_2_14_6  (
            .in0(N__8843),
            .in1(N__11867),
            .in2(N__8828),
            .in3(N__9482),
            .lcout(\b2v_inst.un1_pix_count_anterior_0_I_51_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.pix_count_anterior_9_LC_2_14_7 .C_ON=1'b0;
    defparam \b2v_inst.pix_count_anterior_9_LC_2_14_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.pix_count_anterior_9_LC_2_14_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst.pix_count_anterior_9_LC_2_14_7  (
            .in0(N__11869),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst.pix_count_anteriorZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22588),
            .ce(N__9341),
            .sr(N__22883));
    defparam \b2v_inst.ignorar_ancho_1_LC_2_15_0 .C_ON=1'b0;
    defparam \b2v_inst.ignorar_ancho_1_LC_2_15_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.ignorar_ancho_1_LC_2_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.ignorar_ancho_1_LC_2_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15678),
            .lcout(\b2v_inst.ignorar_anchoZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22578),
            .ce(N__8819),
            .sr(N__22887));
    defparam \b2v_inst.data_a_escribir9_0_c_RNO_LC_2_16_0 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir9_0_c_RNO_LC_2_16_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir9_0_c_RNO_LC_2_16_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst.data_a_escribir9_0_c_RNO_LC_2_16_0  (
            .in0(N__11060),
            .in1(N__11156),
            .in2(N__11022),
            .in3(N__10282),
            .lcout(\b2v_inst.data_a_escribir9_0_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.reg_ancho_1_0_LC_2_16_1 .C_ON=1'b0;
    defparam \b2v_inst.reg_ancho_1_0_LC_2_16_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_ancho_1_0_LC_2_16_1 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \b2v_inst.reg_ancho_1_0_LC_2_16_1  (
            .in0(N__13095),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8878),
            .lcout(\b2v_inst.reg_ancho_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22606),
            .ce(N__13912),
            .sr(N__22892));
    defparam \b2v_inst.reg_ancho_1_1_LC_2_16_2 .C_ON=1'b0;
    defparam \b2v_inst.reg_ancho_1_1_LC_2_16_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_ancho_1_1_LC_2_16_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \b2v_inst.reg_ancho_1_1_LC_2_16_2  (
            .in0(N__8879),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13020),
            .lcout(\b2v_inst.reg_ancho_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22606),
            .ce(N__13912),
            .sr(N__22892));
    defparam \b2v_inst.reg_ancho_1_2_LC_2_16_3 .C_ON=1'b0;
    defparam \b2v_inst.reg_ancho_1_2_LC_2_16_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_ancho_1_2_LC_2_16_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \b2v_inst.reg_ancho_1_2_LC_2_16_3  (
            .in0(_gnd_net_),
            .in1(N__8880),
            .in2(_gnd_net_),
            .in3(N__12951),
            .lcout(\b2v_inst.reg_ancho_1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22606),
            .ce(N__13912),
            .sr(N__22892));
    defparam \b2v_inst.reg_ancho_1_3_LC_2_16_4 .C_ON=1'b0;
    defparam \b2v_inst.reg_ancho_1_3_LC_2_16_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_ancho_1_3_LC_2_16_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \b2v_inst.reg_ancho_1_3_LC_2_16_4  (
            .in0(N__8881),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12879),
            .lcout(\b2v_inst.reg_ancho_1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22606),
            .ce(N__13912),
            .sr(N__22892));
    defparam \b2v_inst.reg_ancho_1_4_LC_2_16_5 .C_ON=1'b0;
    defparam \b2v_inst.reg_ancho_1_4_LC_2_16_5 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_ancho_1_4_LC_2_16_5 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \b2v_inst.reg_ancho_1_4_LC_2_16_5  (
            .in0(N__13545),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8882),
            .lcout(\b2v_inst.reg_ancho_1Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22606),
            .ce(N__13912),
            .sr(N__22892));
    defparam \b2v_inst.data_a_escribir9_1_c_RNO_LC_2_16_6 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir9_1_c_RNO_LC_2_16_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir9_1_c_RNO_LC_2_16_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst.data_a_escribir9_1_c_RNO_LC_2_16_6  (
            .in0(N__10829),
            .in1(N__10871),
            .in2(N__10794),
            .in3(N__10946),
            .lcout(\b2v_inst.data_a_escribir9_1_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.reg_ancho_1_5_LC_2_16_7 .C_ON=1'b0;
    defparam \b2v_inst.reg_ancho_1_5_LC_2_16_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_ancho_1_5_LC_2_16_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \b2v_inst.reg_ancho_1_5_LC_2_16_7  (
            .in0(_gnd_net_),
            .in1(N__14693),
            .in2(_gnd_net_),
            .in3(N__8883),
            .lcout(\b2v_inst.reg_ancho_1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22606),
            .ce(N__13912),
            .sr(N__22892));
    defparam \b2v_inst.data_a_escribir9_3_c_RNO_LC_2_17_0 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir9_3_c_RNO_LC_2_17_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir9_3_c_RNO_LC_2_17_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst.data_a_escribir9_3_c_RNO_LC_2_17_0  (
            .in0(N__11242),
            .in1(N__11293),
            .in2(N__11203),
            .in3(N__11326),
            .lcout(\b2v_inst.data_a_escribir9_3_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.reg_ancho_2_4_LC_2_17_1 .C_ON=1'b0;
    defparam \b2v_inst.reg_ancho_2_4_LC_2_17_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_ancho_2_4_LC_2_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.reg_ancho_2_4_LC_2_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13553),
            .lcout(\b2v_inst.reg_ancho_2Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22564),
            .ce(N__15490),
            .sr(N__22897));
    defparam \b2v_inst.reg_ancho_2_5_LC_2_17_2 .C_ON=1'b0;
    defparam \b2v_inst.reg_ancho_2_5_LC_2_17_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_ancho_2_5_LC_2_17_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.reg_ancho_2_5_LC_2_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14704),
            .lcout(\b2v_inst.reg_ancho_2Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22564),
            .ce(N__15490),
            .sr(N__22897));
    defparam \b2v_inst.reg_ancho_2_6_LC_2_17_3 .C_ON=1'b0;
    defparam \b2v_inst.reg_ancho_2_6_LC_2_17_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_ancho_2_6_LC_2_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.reg_ancho_2_6_LC_2_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14243),
            .lcout(\b2v_inst.reg_ancho_2Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22564),
            .ce(N__15490),
            .sr(N__22897));
    defparam \b2v_inst.reg_ancho_2_7_LC_2_17_4 .C_ON=1'b0;
    defparam \b2v_inst.reg_ancho_2_7_LC_2_17_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_ancho_2_7_LC_2_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.reg_ancho_2_7_LC_2_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13642),
            .lcout(\b2v_inst.reg_ancho_2Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22564),
            .ce(N__15490),
            .sr(N__22897));
    defparam \b2v_inst.data_a_escribir_RNO_3_4_LC_2_17_5 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_3_4_LC_2_17_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_3_4_LC_2_17_5 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_3_4_LC_2_17_5  (
            .in0(N__11327),
            .in1(N__10516),
            .in2(_gnd_net_),
            .in3(N__10679),
            .lcout(),
            .ltout(\b2v_inst.data_a_escribir_RNO_3Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_0_4_LC_2_17_6 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_0_4_LC_2_17_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_0_4_LC_2_17_6 .LUT_INIT=16'b0000111100000011;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_0_4_LC_2_17_6  (
            .in0(_gnd_net_),
            .in1(N__9668),
            .in2(N__8933),
            .in3(N__10950),
            .lcout(\b2v_inst.data_a_escribir_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_un3_valor_max1_cry_7_c_RNIV45S_LC_2_17_7 .C_ON=1'b0;
    defparam \b2v_inst.encontrar_maximo_un3_valor_max1_cry_7_c_RNIV45S_LC_2_17_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_un3_valor_max1_cry_7_c_RNIV45S_LC_2_17_7 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \b2v_inst.encontrar_maximo_un3_valor_max1_cry_7_c_RNIV45S_LC_2_17_7  (
            .in0(_gnd_net_),
            .in1(N__10515),
            .in2(_gnd_net_),
            .in3(N__10678),
            .lcout(\b2v_inst.un1_reg_anterior_iv_0_0_a2_4_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_3_0_LC_2_18_0 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_3_0_LC_2_18_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_3_0_LC_2_18_0 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_3_0_LC_2_18_0  (
            .in0(N__10250),
            .in1(N__10557),
            .in2(_gnd_net_),
            .in3(N__13219),
            .lcout(),
            .ltout(\b2v_inst.data_a_escribir_RNO_3Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_1_0_LC_2_18_1 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_1_0_LC_2_18_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_1_0_LC_2_18_1 .LUT_INIT=16'b0000111100000011;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_1_0_LC_2_18_1  (
            .in0(_gnd_net_),
            .in1(N__10611),
            .in2(N__8930),
            .in3(N__13067),
            .lcout(),
            .ltout(\b2v_inst.data_a_escribir_RNO_1Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_0_LC_2_18_2 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_0_LC_2_18_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.data_a_escribir_0_LC_2_18_2 .LUT_INIT=16'b0100010001010000;
    LogicCell40 \b2v_inst.data_a_escribir_0_LC_2_18_2  (
            .in0(N__8927),
            .in1(N__8915),
            .in2(N__8909),
            .in3(N__10431),
            .lcout(b2v_inst_data_a_escribir_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22607),
            .ce(N__10350),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_3_3_LC_2_18_3 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_3_3_LC_2_18_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_3_3_LC_2_18_3 .LUT_INIT=16'b1010100011111111;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_3_3_LC_2_18_3  (
            .in0(N__8906),
            .in1(N__10426),
            .in2(N__10569),
            .in3(N__14797),
            .lcout(\b2v_inst.un1_reg_anterior_iv_0_0_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_0_3_LC_2_18_4 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_0_3_LC_2_18_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_0_3_LC_2_18_4 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_0_3_LC_2_18_4  (
            .in0(N__10706),
            .in1(N__10558),
            .in2(N__11390),
            .in3(N__10430),
            .lcout(),
            .ltout(\b2v_inst.N_315_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_3_LC_2_18_5 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_3_LC_2_18_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.data_a_escribir_3_LC_2_18_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst.data_a_escribir_3_LC_2_18_5  (
            .in0(N__8978),
            .in1(N__8942),
            .in2(N__8897),
            .in3(N__8894),
            .lcout(b2v_inst_data_a_escribir_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22607),
            .ce(N__10350),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_un3_valor_max2_cry_7_c_RNI0D1L_LC_2_18_6 .C_ON=1'b0;
    defparam \b2v_inst.encontrar_maximo_un3_valor_max2_cry_7_c_RNI0D1L_LC_2_18_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_un3_valor_max2_cry_7_c_RNI0D1L_LC_2_18_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \b2v_inst.encontrar_maximo_un3_valor_max2_cry_7_c_RNI0D1L_LC_2_18_6  (
            .in0(_gnd_net_),
            .in1(N__10553),
            .in2(_gnd_net_),
            .in3(N__13218),
            .lcout(\b2v_inst.un1_reg_anterior_iv_0_0_a2_6_0_1 ),
            .ltout(\b2v_inst.un1_reg_anterior_iv_0_0_a2_6_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_1_3_LC_2_18_7 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_1_3_LC_2_18_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_1_3_LC_2_18_7 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_1_3_LC_2_18_7  (
            .in0(_gnd_net_),
            .in1(N__10425),
            .in2(N__8888),
            .in3(N__12851),
            .lcout(\b2v_inst.N_317 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir9_2_c_RNO_LC_2_19_0 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir9_2_c_RNO_LC_2_19_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir9_2_c_RNO_LC_2_19_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst.data_a_escribir9_2_c_RNO_LC_2_19_0  (
            .in0(N__11419),
            .in1(N__11458),
            .in2(N__11387),
            .in3(N__11506),
            .lcout(\b2v_inst.data_a_escribir9_2_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.reg_ancho_2_0_LC_2_19_1 .C_ON=1'b0;
    defparam \b2v_inst.reg_ancho_2_0_LC_2_19_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_ancho_2_0_LC_2_19_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.reg_ancho_2_0_LC_2_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13103),
            .lcout(\b2v_inst.reg_ancho_2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22597),
            .ce(N__15491),
            .sr(N__22907));
    defparam \b2v_inst.reg_ancho_2_1_LC_2_19_2 .C_ON=1'b0;
    defparam \b2v_inst.reg_ancho_2_1_LC_2_19_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_ancho_2_1_LC_2_19_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.reg_ancho_2_1_LC_2_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13031),
            .lcout(\b2v_inst.reg_ancho_2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22597),
            .ce(N__15491),
            .sr(N__22907));
    defparam \b2v_inst.reg_ancho_2_2_LC_2_19_3 .C_ON=1'b0;
    defparam \b2v_inst.reg_ancho_2_2_LC_2_19_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_ancho_2_2_LC_2_19_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.reg_ancho_2_2_LC_2_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12959),
            .lcout(\b2v_inst.reg_ancho_2Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22597),
            .ce(N__15491),
            .sr(N__22907));
    defparam \b2v_inst.reg_ancho_2_3_LC_2_19_4 .C_ON=1'b0;
    defparam \b2v_inst.reg_ancho_2_3_LC_2_19_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_ancho_2_3_LC_2_19_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.reg_ancho_2_3_LC_2_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12887),
            .lcout(\b2v_inst.reg_ancho_2Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22597),
            .ce(N__15491),
            .sr(N__22907));
    defparam \b2v_inst.data_a_escribir_RNO_2_2_LC_2_19_6 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_2_2_LC_2_19_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_2_2_LC_2_19_6 .LUT_INIT=16'b1100101000000000;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_2_2_LC_2_19_6  (
            .in0(N__11635),
            .in1(N__9727),
            .in2(N__13238),
            .in3(N__8972),
            .lcout(),
            .ltout(\b2v_inst.N_320_tz_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_0_2_LC_2_19_7 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_0_2_LC_2_19_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_0_2_LC_2_19_7 .LUT_INIT=16'b0111011111110011;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_0_2_LC_2_19_7  (
            .in0(N__8966),
            .in1(N__14798),
            .in2(N__8948),
            .in3(N__10563),
            .lcout(\b2v_inst.un1_reg_anterior_iv_0_0_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_0_cry_7_c_RNI5KAH1_LC_2_20_1 .C_ON=1'b0;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_0_cry_7_c_RNI5KAH1_LC_2_20_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_0_cry_7_c_RNI5KAH1_LC_2_20_1 .LUT_INIT=16'b0101010100011011;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final5_0_cry_7_c_RNI5KAH1_LC_2_20_1  (
            .in0(N__10688),
            .in1(N__10727),
            .in2(N__11636),
            .in3(N__13227),
            .lcout(\b2v_inst.un1_m3_0_m3_ns_1 ),
            .ltout(\b2v_inst.un1_m3_0_m3_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_2_3_LC_2_20_2 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_2_3_LC_2_20_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_2_3_LC_2_20_2 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_2_3_LC_2_20_2  (
            .in0(N__13228),
            .in1(N__10562),
            .in2(N__8945),
            .in3(N__10988),
            .lcout(\b2v_inst.N_318 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_4_LC_2_20_3 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_4_LC_2_20_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.data_a_escribir_4_LC_2_20_3 .LUT_INIT=16'b0000110000000101;
    LogicCell40 \b2v_inst.data_a_escribir_4_LC_2_20_3  (
            .in0(N__9899),
            .in1(N__9074),
            .in2(N__9065),
            .in3(N__10419),
            .lcout(b2v_inst_data_a_escribir_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22596),
            .ce(N__10349),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNIA6JL_4_LC_2_20_4 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNIA6JL_4_LC_2_20_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNIA6JL_4_LC_2_20_4 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \b2v_inst.data_a_escribir_RNIA6JL_4_LC_2_20_4  (
            .in0(N__17717),
            .in1(N__17033),
            .in2(_gnd_net_),
            .in3(N__14509),
            .lcout(N_211_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNI62JL_0_LC_2_20_5 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNI62JL_0_LC_2_20_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNI62JL_0_LC_2_20_5 .LUT_INIT=16'b1111000010100000;
    LogicCell40 \b2v_inst.data_a_escribir_RNI62JL_0_LC_2_20_5  (
            .in0(N__17031),
            .in1(_gnd_net_),
            .in2(N__13459),
            .in3(N__17716),
            .lcout(N_219_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNI73JL_1_LC_2_20_6 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNI73JL_1_LC_2_20_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNI73JL_1_LC_2_20_6 .LUT_INIT=16'b1111000011000000;
    LogicCell40 \b2v_inst.data_a_escribir_RNI73JL_1_LC_2_20_6  (
            .in0(_gnd_net_),
            .in1(N__17032),
            .in2(N__13480),
            .in3(N__17714),
            .lcout(N_217_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNI84JL_2_LC_2_20_7 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNI84JL_2_LC_2_20_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNI84JL_2_LC_2_20_7 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \b2v_inst.data_a_escribir_RNI84JL_2_LC_2_20_7  (
            .in0(N__17030),
            .in1(N__13411),
            .in2(_gnd_net_),
            .in3(N__17715),
            .lcout(N_215_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_11_LC_3_11_0 .C_ON=1'b0;
    defparam \b2v_inst.state_11_LC_3_11_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.state_11_LC_3_11_0 .LUT_INIT=16'b0010101000000000;
    LogicCell40 \b2v_inst.state_11_LC_3_11_0  (
            .in0(N__15682),
            .in1(N__9125),
            .in2(N__8993),
            .in3(N__10208),
            .lcout(\b2v_inst.stateZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22481),
            .ce(),
            .sr(N__22878));
    defparam \b2v_inst.state_ns_i_i_a2_4_6_LC_3_11_1 .C_ON=1'b0;
    defparam \b2v_inst.state_ns_i_i_a2_4_6_LC_3_11_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_ns_i_i_a2_4_6_LC_3_11_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst.state_ns_i_i_a2_4_6_LC_3_11_1  (
            .in0(N__10070),
            .in1(N__10082),
            .in2(N__10058),
            .in3(N__10094),
            .lcout(\b2v_inst.state_ns_i_i_a2_4Z0Z_6 ),
            .ltout(\b2v_inst.state_ns_i_i_a2_4Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un1_pix_count_anterior_0_I_39_c_RNIP5QR3_LC_3_11_2 .C_ON=1'b0;
    defparam \b2v_inst.un1_pix_count_anterior_0_I_39_c_RNIP5QR3_LC_3_11_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un1_pix_count_anterior_0_I_39_c_RNIP5QR3_LC_3_11_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst.un1_pix_count_anterior_0_I_39_c_RNIP5QR3_LC_3_11_2  (
            .in0(N__15681),
            .in1(N__9124),
            .in2(N__8984),
            .in3(N__10207),
            .lcout(\b2v_inst.N_497 ),
            .ltout(\b2v_inst.N_497_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_6_LC_3_11_3 .C_ON=1'b0;
    defparam \b2v_inst.state_6_LC_3_11_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.state_6_LC_3_11_3 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \b2v_inst.state_6_LC_3_11_3  (
            .in0(N__9134),
            .in1(N__14791),
            .in2(N__8981),
            .in3(N__14873),
            .lcout(\b2v_inst.stateZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22481),
            .ce(),
            .sr(N__22878));
    defparam \b2v_inst.state_RNO_0_6_LC_3_11_4 .C_ON=1'b0;
    defparam \b2v_inst.state_RNO_0_6_LC_3_11_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNO_0_6_LC_3_11_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst.state_RNO_0_6_LC_3_11_4  (
            .in0(_gnd_net_),
            .in1(N__17702),
            .in2(_gnd_net_),
            .in3(N__15680),
            .lcout(\b2v_inst.N_361 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_ns_i_i_a2_5_6_LC_3_11_5 .C_ON=1'b0;
    defparam \b2v_inst.state_ns_i_i_a2_5_6_LC_3_11_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_ns_i_i_a2_5_6_LC_3_11_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst.state_ns_i_i_a2_5_6_LC_3_11_5  (
            .in0(N__9911),
            .in1(N__9923),
            .in2(N__10043),
            .in3(N__9935),
            .lcout(\b2v_inst.state_ns_i_i_a2_5Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un1_pix_count_anterior_0_I_39_c_RNIT6R7_LC_3_11_6 .C_ON=1'b0;
    defparam \b2v_inst.un1_pix_count_anterior_0_I_39_c_RNIT6R7_LC_3_11_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un1_pix_count_anterior_0_I_39_c_RNIT6R7_LC_3_11_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst.un1_pix_count_anterior_0_I_39_c_RNIT6R7_LC_3_11_6  (
            .in0(_gnd_net_),
            .in1(N__15679),
            .in2(_gnd_net_),
            .in3(N__10206),
            .lcout(\b2v_inst.N_254_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.borrado_LC_3_11_7 .C_ON=1'b0;
    defparam \b2v_inst.borrado_LC_3_11_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.borrado_LC_3_11_7 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \b2v_inst.borrado_LC_3_11_7  (
            .in0(N__17703),
            .in1(N__15901),
            .in2(_gnd_net_),
            .in3(N__18776),
            .lcout(\b2v_inst.borradoZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22481),
            .ce(),
            .sr(N__22878));
    defparam \b2v_inst.un1_pix_count_anterior_0_I_27_c_RNO_LC_3_12_0 .C_ON=1'b0;
    defparam \b2v_inst.un1_pix_count_anterior_0_I_27_c_RNO_LC_3_12_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un1_pix_count_anterior_0_I_27_c_RNO_LC_3_12_0 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \b2v_inst.un1_pix_count_anterior_0_I_27_c_RNO_LC_3_12_0  (
            .in0(N__9107),
            .in1(N__9233),
            .in2(N__9095),
            .in3(N__9257),
            .lcout(\b2v_inst.un1_pix_count_anterior_0_I_27_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.pix_count_anterior_3_LC_3_12_1 .C_ON=1'b0;
    defparam \b2v_inst.pix_count_anterior_3_LC_3_12_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.pix_count_anterior_3_LC_3_12_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst.pix_count_anterior_3_LC_3_12_1  (
            .in0(N__9235),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst.pix_count_anteriorZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22380),
            .ce(N__9340),
            .sr(N__22881));
    defparam \b2v_inst4.pix_count_int_RNIATHH1_0_LC_3_12_2 .C_ON=1'b0;
    defparam \b2v_inst4.pix_count_int_RNIATHH1_0_LC_3_12_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst4.pix_count_int_RNIATHH1_0_LC_3_12_2 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \b2v_inst4.pix_count_int_RNIATHH1_0_LC_3_12_2  (
            .in0(N__9454),
            .in1(N__9234),
            .in2(N__9317),
            .in3(N__15721),
            .lcout(\b2v_inst4.un1_pix_count_int_0_sqmuxa_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.pix_count_anterior_10_LC_3_12_3 .C_ON=1'b0;
    defparam \b2v_inst.pix_count_anterior_10_LC_3_12_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.pix_count_anterior_10_LC_3_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.pix_count_anterior_10_LC_3_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9455),
            .lcout(\b2v_inst.pix_count_anteriorZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22380),
            .ce(N__9340),
            .sr(N__22881));
    defparam \b2v_inst.un1_pix_count_anterior_0_I_9_c_RNO_LC_3_12_4 .C_ON=1'b0;
    defparam \b2v_inst.un1_pix_count_anterior_0_I_9_c_RNO_LC_3_12_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un1_pix_count_anterior_0_I_9_c_RNO_LC_3_12_4 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \b2v_inst.un1_pix_count_anterior_0_I_9_c_RNO_LC_3_12_4  (
            .in0(N__9086),
            .in1(N__9425),
            .in2(N__9350),
            .in3(N__9453),
            .lcout(\b2v_inst.un1_pix_count_anterior_0_I_9_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.pix_count_anterior_11_LC_3_12_5 .C_ON=1'b0;
    defparam \b2v_inst.pix_count_anterior_11_LC_3_12_5 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.pix_count_anterior_11_LC_3_12_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst.pix_count_anterior_11_LC_3_12_5  (
            .in0(N__9426),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst.pix_count_anteriorZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22380),
            .ce(N__9340),
            .sr(N__22881));
    defparam \b2v_inst4.state_RNICJOG_0_LC_3_12_6 .C_ON=1'b0;
    defparam \b2v_inst4.state_RNICJOG_0_LC_3_12_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst4.state_RNICJOG_0_LC_3_12_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \b2v_inst4.state_RNICJOG_0_LC_3_12_6  (
            .in0(_gnd_net_),
            .in1(N__11713),
            .in2(_gnd_net_),
            .in3(N__15720),
            .lcout(\b2v_inst4.pix_count_int_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst4.pix_count_int_RNO_0_0_LC_3_13_0 .C_ON=1'b1;
    defparam \b2v_inst4.pix_count_int_RNO_0_0_LC_3_13_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst4.pix_count_int_RNO_0_0_LC_3_13_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst4.pix_count_int_RNO_0_0_LC_3_13_0  (
            .in0(_gnd_net_),
            .in1(N__9310),
            .in2(N__10027),
            .in3(N__10023),
            .lcout(\b2v_inst4.pix_count_int_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(bfn_3_13_0_),
            .carryout(\b2v_inst4.un1_pix_count_int_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst4.pix_count_int_1_LC_3_13_1 .C_ON=1'b1;
    defparam \b2v_inst4.pix_count_int_1_LC_3_13_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst4.pix_count_int_1_LC_3_13_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst4.pix_count_int_1_LC_3_13_1  (
            .in0(_gnd_net_),
            .in1(N__9284),
            .in2(_gnd_net_),
            .in3(N__9266),
            .lcout(SYNTHESIZED_WIRE_2_1),
            .ltout(),
            .carryin(\b2v_inst4.un1_pix_count_int_cry_0 ),
            .carryout(\b2v_inst4.un1_pix_count_int_cry_1 ),
            .clk(N__22482),
            .ce(),
            .sr(N__22884));
    defparam \b2v_inst4.pix_count_int_2_LC_3_13_2 .C_ON=1'b1;
    defparam \b2v_inst4.pix_count_int_2_LC_3_13_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst4.pix_count_int_2_LC_3_13_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst4.pix_count_int_2_LC_3_13_2  (
            .in0(_gnd_net_),
            .in1(N__9258),
            .in2(_gnd_net_),
            .in3(N__9239),
            .lcout(SYNTHESIZED_WIRE_2_2),
            .ltout(),
            .carryin(\b2v_inst4.un1_pix_count_int_cry_1 ),
            .carryout(\b2v_inst4.un1_pix_count_int_cry_2 ),
            .clk(N__22482),
            .ce(),
            .sr(N__22884));
    defparam \b2v_inst4.pix_count_int_RNO_0_3_LC_3_13_3 .C_ON=1'b1;
    defparam \b2v_inst4.pix_count_int_RNO_0_3_LC_3_13_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst4.pix_count_int_RNO_0_3_LC_3_13_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst4.pix_count_int_RNO_0_3_LC_3_13_3  (
            .in0(_gnd_net_),
            .in1(N__9236),
            .in2(_gnd_net_),
            .in3(N__9212),
            .lcout(\b2v_inst4.pix_count_int_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(\b2v_inst4.un1_pix_count_int_cry_2 ),
            .carryout(\b2v_inst4.un1_pix_count_int_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst4.pix_count_int_4_LC_3_13_4 .C_ON=1'b1;
    defparam \b2v_inst4.pix_count_int_4_LC_3_13_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst4.pix_count_int_4_LC_3_13_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst4.pix_count_int_4_LC_3_13_4  (
            .in0(_gnd_net_),
            .in1(N__9209),
            .in2(_gnd_net_),
            .in3(N__9191),
            .lcout(SYNTHESIZED_WIRE_2_4),
            .ltout(),
            .carryin(\b2v_inst4.un1_pix_count_int_cry_3 ),
            .carryout(\b2v_inst4.un1_pix_count_int_cry_4 ),
            .clk(N__22482),
            .ce(),
            .sr(N__22884));
    defparam \b2v_inst4.pix_count_int_RNO_0_5_LC_3_13_5 .C_ON=1'b1;
    defparam \b2v_inst4.pix_count_int_RNO_0_5_LC_3_13_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst4.pix_count_int_RNO_0_5_LC_3_13_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst4.pix_count_int_RNO_0_5_LC_3_13_5  (
            .in0(_gnd_net_),
            .in1(N__9187),
            .in2(_gnd_net_),
            .in3(N__9161),
            .lcout(\b2v_inst4.pix_count_int_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\b2v_inst4.un1_pix_count_int_cry_4 ),
            .carryout(\b2v_inst4.un1_pix_count_int_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst4.pix_count_int_6_LC_3_13_6 .C_ON=1'b1;
    defparam \b2v_inst4.pix_count_int_6_LC_3_13_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst4.pix_count_int_6_LC_3_13_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst4.pix_count_int_6_LC_3_13_6  (
            .in0(_gnd_net_),
            .in1(N__9157),
            .in2(_gnd_net_),
            .in3(N__9137),
            .lcout(SYNTHESIZED_WIRE_2_6),
            .ltout(),
            .carryin(\b2v_inst4.un1_pix_count_int_cry_5 ),
            .carryout(\b2v_inst4.un1_pix_count_int_cry_6 ),
            .clk(N__22482),
            .ce(),
            .sr(N__22884));
    defparam \b2v_inst4.pix_count_int_RNO_0_7_LC_3_13_7 .C_ON=1'b1;
    defparam \b2v_inst4.pix_count_int_RNO_0_7_LC_3_13_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst4.pix_count_int_RNO_0_7_LC_3_13_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst4.pix_count_int_RNO_0_7_LC_3_13_7  (
            .in0(_gnd_net_),
            .in1(N__9512),
            .in2(_gnd_net_),
            .in3(N__9488),
            .lcout(\b2v_inst4.pix_count_int_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(\b2v_inst4.un1_pix_count_int_cry_6 ),
            .carryout(\b2v_inst4.un1_pix_count_int_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst4.pix_count_int_RNO_0_8_LC_3_14_0 .C_ON=1'b1;
    defparam \b2v_inst4.pix_count_int_RNO_0_8_LC_3_14_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst4.pix_count_int_RNO_0_8_LC_3_14_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst4.pix_count_int_RNO_0_8_LC_3_14_0  (
            .in0(_gnd_net_),
            .in1(N__9485),
            .in2(_gnd_net_),
            .in3(N__9461),
            .lcout(\b2v_inst4.pix_count_int_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(bfn_3_14_0_),
            .carryout(\b2v_inst4.un1_pix_count_int_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst4.pix_count_int_RNO_0_9_LC_3_14_1 .C_ON=1'b1;
    defparam \b2v_inst4.pix_count_int_RNO_0_9_LC_3_14_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst4.pix_count_int_RNO_0_9_LC_3_14_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst4.pix_count_int_RNO_0_9_LC_3_14_1  (
            .in0(_gnd_net_),
            .in1(N__11870),
            .in2(_gnd_net_),
            .in3(N__9458),
            .lcout(\b2v_inst4.pix_count_int_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(\b2v_inst4.un1_pix_count_int_cry_8 ),
            .carryout(\b2v_inst4.un1_pix_count_int_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst4.pix_count_int_10_LC_3_14_2 .C_ON=1'b1;
    defparam \b2v_inst4.pix_count_int_10_LC_3_14_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst4.pix_count_int_10_LC_3_14_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst4.pix_count_int_10_LC_3_14_2  (
            .in0(_gnd_net_),
            .in1(N__9452),
            .in2(_gnd_net_),
            .in3(N__9431),
            .lcout(SYNTHESIZED_WIRE_2_10),
            .ltout(),
            .carryin(\b2v_inst4.un1_pix_count_int_cry_9 ),
            .carryout(\b2v_inst4.un1_pix_count_int_cry_10 ),
            .clk(N__22381),
            .ce(),
            .sr(N__22888));
    defparam \b2v_inst4.pix_count_int_RNO_0_11_LC_3_14_3 .C_ON=1'b1;
    defparam \b2v_inst4.pix_count_int_RNO_0_11_LC_3_14_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst4.pix_count_int_RNO_0_11_LC_3_14_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst4.pix_count_int_RNO_0_11_LC_3_14_3  (
            .in0(_gnd_net_),
            .in1(N__9427),
            .in2(_gnd_net_),
            .in3(N__9401),
            .lcout(\b2v_inst4.pix_count_int_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(\b2v_inst4.un1_pix_count_int_cry_10 ),
            .carryout(\b2v_inst4.un1_pix_count_int_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst4.pix_count_int_RNO_0_12_LC_3_14_4 .C_ON=1'b0;
    defparam \b2v_inst4.pix_count_int_RNO_0_12_LC_3_14_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst4.pix_count_int_RNO_0_12_LC_3_14_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \b2v_inst4.pix_count_int_RNO_0_12_LC_3_14_4  (
            .in0(_gnd_net_),
            .in1(N__9396),
            .in2(_gnd_net_),
            .in3(N__9371),
            .lcout(\b2v_inst4.pix_count_int_RNO_0Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir9_0_c_LC_3_15_0 .C_ON=1'b1;
    defparam \b2v_inst.data_a_escribir9_0_c_LC_3_15_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir9_0_c_LC_3_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.data_a_escribir9_0_c_LC_3_15_0  (
            .in0(_gnd_net_),
            .in1(N__9362),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_3_15_0_),
            .carryout(\b2v_inst.data_a_escribir9_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir9_1_c_LC_3_15_1 .C_ON=1'b1;
    defparam \b2v_inst.data_a_escribir9_1_c_LC_3_15_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir9_1_c_LC_3_15_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.data_a_escribir9_1_c_LC_3_15_1  (
            .in0(_gnd_net_),
            .in1(N__9356),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.data_a_escribir9_0 ),
            .carryout(\b2v_inst.data_a_escribir9_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir9_2_c_LC_3_15_2 .C_ON=1'b1;
    defparam \b2v_inst.data_a_escribir9_2_c_LC_3_15_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir9_2_c_LC_3_15_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.data_a_escribir9_2_c_LC_3_15_2  (
            .in0(_gnd_net_),
            .in1(N__9554),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.data_a_escribir9_1 ),
            .carryout(\b2v_inst.data_a_escribir9_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir9_3_c_LC_3_15_3 .C_ON=1'b1;
    defparam \b2v_inst.data_a_escribir9_3_c_LC_3_15_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir9_3_c_LC_3_15_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.data_a_escribir9_3_c_LC_3_15_3  (
            .in0(_gnd_net_),
            .in1(N__9542),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.data_a_escribir9_2 ),
            .carryout(\b2v_inst.data_a_escribir9_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir9_4_c_LC_3_15_4 .C_ON=1'b1;
    defparam \b2v_inst.data_a_escribir9_4_c_LC_3_15_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir9_4_c_LC_3_15_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.data_a_escribir9_4_c_LC_3_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10106),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.data_a_escribir9_3 ),
            .carryout(\b2v_inst.data_a_escribir9_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir9_5_c_LC_3_15_5 .C_ON=1'b1;
    defparam \b2v_inst.data_a_escribir9_5_c_LC_3_15_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir9_5_c_LC_3_15_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.data_a_escribir9_5_c_LC_3_15_5  (
            .in0(_gnd_net_),
            .in1(N__10715),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.data_a_escribir9_4 ),
            .carryout(\b2v_inst.data_a_escribir9_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir9_6_c_LC_3_15_6 .C_ON=1'b1;
    defparam \b2v_inst.data_a_escribir9_6_c_LC_3_15_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir9_6_c_LC_3_15_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.data_a_escribir9_6_c_LC_3_15_6  (
            .in0(_gnd_net_),
            .in1(N__11525),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.data_a_escribir9_5 ),
            .carryout(\b2v_inst.data_a_escribir9_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir9_7_c_LC_3_15_7 .C_ON=1'b1;
    defparam \b2v_inst.data_a_escribir9_7_c_LC_3_15_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir9_7_c_LC_3_15_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.data_a_escribir9_7_c_LC_3_15_7  (
            .in0(_gnd_net_),
            .in1(N__13568),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.data_a_escribir9_6 ),
            .carryout(\b2v_inst.data_a_escribir10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir10_THRU_LUT4_0_LC_3_16_0 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir10_THRU_LUT4_0_LC_3_16_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir10_THRU_LUT4_0_LC_3_16_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.data_a_escribir10_THRU_LUT4_0_LC_3_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9533),
            .lcout(\b2v_inst.data_a_escribir10_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_RX_Byte_0_LC_3_16_1 .C_ON=1'b0;
    defparam \b2v_inst1.r_RX_Byte_0_LC_3_16_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst1.r_RX_Byte_0_LC_3_16_1 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \b2v_inst1.r_RX_Byte_0_LC_3_16_1  (
            .in0(N__17126),
            .in1(N__9946),
            .in2(N__22751),
            .in3(N__17177),
            .lcout(SYNTHESIZED_WIRE_10_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22605),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_0_7_LC_3_16_3 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_0_7_LC_3_16_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_0_7_LC_3_16_3 .LUT_INIT=16'b0010001011111111;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_0_7_LC_3_16_3  (
            .in0(N__10511),
            .in1(N__9530),
            .in2(_gnd_net_),
            .in3(N__14785),
            .lcout(\b2v_inst.un1_reg_anterior_iv_0_0_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_2_1_LC_3_16_4 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_2_1_LC_3_16_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_2_1_LC_3_16_4 .LUT_INIT=16'b0111011101010101;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_2_1_LC_3_16_4  (
            .in0(N__14787),
            .in1(N__9611),
            .in2(_gnd_net_),
            .in3(N__10514),
            .lcout(\b2v_inst.un1_reg_anterior_iv_0_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_3_2_LC_3_16_5 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_3_2_LC_3_16_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_3_2_LC_3_16_5 .LUT_INIT=16'b0000010100010001;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_3_2_LC_3_16_5  (
            .in0(N__10513),
            .in1(N__11102),
            .in2(N__12923),
            .in3(N__13232),
            .lcout(\b2v_inst.un1_reg_anterior_iv_0_0_2_tz_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_3_6_LC_3_16_6 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_3_6_LC_3_16_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_3_6_LC_3_16_6 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_3_6_LC_3_16_6  (
            .in0(N__13231),
            .in1(N__10510),
            .in2(_gnd_net_),
            .in3(N__12812),
            .lcout(\b2v_inst.data_a_escribir_RNO_3Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_2_6_LC_3_16_7 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_2_6_LC_3_16_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_2_6_LC_3_16_7 .LUT_INIT=16'b0010001011111111;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_2_6_LC_3_16_7  (
            .in0(N__10512),
            .in1(N__9593),
            .in2(_gnd_net_),
            .in3(N__14786),
            .lcout(\b2v_inst.un1_reg_anterior_iv_0_0_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_3_1_LC_3_17_1 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_3_1_LC_3_17_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_3_1_LC_3_17_1 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_3_1_LC_3_17_1  (
            .in0(N__11472),
            .in1(N__10517),
            .in2(_gnd_net_),
            .in3(N__10705),
            .lcout(),
            .ltout(\b2v_inst.un1_reg_anterior_iv_0_0_2_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_0_1_LC_3_17_2 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_0_1_LC_3_17_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_0_1_LC_3_17_2 .LUT_INIT=16'b0000111100000011;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_0_1_LC_3_17_2  (
            .in0(_gnd_net_),
            .in1(N__9669),
            .in2(N__9575),
            .in3(N__11163),
            .lcout(\b2v_inst.data_a_escribir_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_4_1_LC_3_17_3 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_4_1_LC_3_17_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_4_1_LC_3_17_3 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_4_1_LC_3_17_3  (
            .in0(N__11129),
            .in1(N__10518),
            .in2(_gnd_net_),
            .in3(N__13237),
            .lcout(),
            .ltout(\b2v_inst.data_a_escribir_RNO_4Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_1_1_LC_3_17_4 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_1_1_LC_3_17_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_1_1_LC_3_17_4 .LUT_INIT=16'b0000110000001111;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_1_1_LC_3_17_4  (
            .in0(_gnd_net_),
            .in1(N__12992),
            .in2(N__9572),
            .in3(N__10612),
            .lcout(),
            .ltout(\b2v_inst.data_a_escribir_RNO_1Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_1_LC_3_17_5 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_1_LC_3_17_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.data_a_escribir_1_LC_3_17_5 .LUT_INIT=16'b0100010001010000;
    LogicCell40 \b2v_inst.data_a_escribir_1_LC_3_17_5  (
            .in0(N__9569),
            .in1(N__9563),
            .in2(N__9557),
            .in3(N__10429),
            .lcout(b2v_inst_data_a_escribir_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22563),
            .ce(N__10352),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNI9HNM5_7_LC_3_17_7 .C_ON=1'b0;
    defparam \b2v_inst.state_RNI9HNM5_7_LC_3_17_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNI9HNM5_7_LC_3_17_7 .LUT_INIT=16'b1111000010110000;
    LogicCell40 \b2v_inst.state_RNI9HNM5_7_LC_3_17_7  (
            .in0(N__14781),
            .in1(N__14872),
            .in2(N__18941),
            .in3(N__9704),
            .lcout(\b2v_inst.un1_reset_inv_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_1_2_LC_3_18_0 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_1_2_LC_3_18_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_1_2_LC_3_18_0 .LUT_INIT=16'b1111001101010101;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_1_2_LC_3_18_0  (
            .in0(N__9695),
            .in1(N__9670),
            .in2(N__11075),
            .in3(N__10427),
            .lcout(),
            .ltout(\b2v_inst.data_a_escribir_RNO_1Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_2_LC_3_18_1 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_2_LC_3_18_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.data_a_escribir_2_LC_3_18_1 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \b2v_inst.data_a_escribir_2_LC_3_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9686),
            .in3(N__9683),
            .lcout(b2v_inst_data_a_escribir_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22565),
            .ce(N__10333),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_4_5_LC_3_18_3 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_4_5_LC_3_18_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_4_5_LC_3_18_3 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_4_5_LC_3_18_3  (
            .in0(N__10540),
            .in1(N__12791),
            .in2(_gnd_net_),
            .in3(N__13223),
            .lcout(),
            .ltout(\b2v_inst.data_a_escribir_RNO_4Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_1_5_LC_3_18_4 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_1_5_LC_3_18_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_1_5_LC_3_18_4 .LUT_INIT=16'b0000110000001111;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_1_5_LC_3_18_4  (
            .in0(_gnd_net_),
            .in1(N__14663),
            .in2(N__9677),
            .in3(N__10610),
            .lcout(\b2v_inst.data_a_escribir_RNO_1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_3_5_LC_3_18_5 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_3_5_LC_3_18_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_3_5_LC_3_18_5 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_3_5_LC_3_18_5  (
            .in0(N__10541),
            .in1(N__11303),
            .in2(_gnd_net_),
            .in3(N__10700),
            .lcout(),
            .ltout(\b2v_inst.un1_reg_anterior_iv_0_0_2_1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_0_5_LC_3_18_6 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_0_5_LC_3_18_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_0_5_LC_3_18_6 .LUT_INIT=16'b0000110000001111;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_0_5_LC_3_18_6  (
            .in0(_gnd_net_),
            .in1(N__10885),
            .in2(N__9674),
            .in3(N__9671),
            .lcout(),
            .ltout(\b2v_inst.data_a_escribir_RNO_0Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_5_LC_3_18_7 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_5_LC_3_18_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.data_a_escribir_5_LC_3_18_7 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \b2v_inst.data_a_escribir_5_LC_3_18_7  (
            .in0(N__10428),
            .in1(N__9650),
            .in2(N__9638),
            .in3(N__9635),
            .lcout(b2v_inst_data_a_escribir_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22565),
            .ce(N__10333),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_1_cry_0_c_inv_LC_3_19_0 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_1_cry_0_c_inv_LC_3_19_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_1_cry_0_c_inv_LC_3_19_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final5_1_cry_0_c_inv_LC_3_19_0  (
            .in0(_gnd_net_),
            .in1(N__10295),
            .in2(N__9629),
            .in3(N__13059),
            .lcout(\b2v_inst.reg_anterior_i_0 ),
            .ltout(),
            .carryin(bfn_3_19_0_),
            .carryout(\b2v_inst.valor_max_final5_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_1_cry_1_c_inv_LC_3_19_1 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_1_cry_1_c_inv_LC_3_19_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_1_cry_1_c_inv_LC_3_19_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final5_1_cry_1_c_inv_LC_3_19_1  (
            .in0(_gnd_net_),
            .in1(N__11167),
            .in2(N__9872),
            .in3(N__12987),
            .lcout(\b2v_inst.reg_anterior_i_1 ),
            .ltout(),
            .carryin(\b2v_inst.valor_max_final5_1_cry_0 ),
            .carryout(\b2v_inst.valor_max_final5_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_1_cry_2_c_inv_LC_3_19_2 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_1_cry_2_c_inv_LC_3_19_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_1_cry_2_c_inv_LC_3_19_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final5_1_cry_2_c_inv_LC_3_19_2  (
            .in0(_gnd_net_),
            .in1(N__11070),
            .in2(N__9854),
            .in3(N__12915),
            .lcout(\b2v_inst.reg_anterior_i_2 ),
            .ltout(),
            .carryin(\b2v_inst.valor_max_final5_1_cry_1 ),
            .carryout(\b2v_inst.valor_max_final5_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_1_cry_3_c_inv_LC_3_19_3 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_1_cry_3_c_inv_LC_3_19_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_1_cry_3_c_inv_LC_3_19_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final5_1_cry_3_c_inv_LC_3_19_3  (
            .in0(_gnd_net_),
            .in1(N__11032),
            .in2(N__9836),
            .in3(N__12845),
            .lcout(\b2v_inst.reg_anterior_i_3 ),
            .ltout(),
            .carryin(\b2v_inst.valor_max_final5_1_cry_2 ),
            .carryout(\b2v_inst.valor_max_final5_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_1_cry_4_c_inv_LC_3_19_4 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_1_cry_4_c_inv_LC_3_19_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_1_cry_4_c_inv_LC_3_19_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final5_1_cry_4_c_inv_LC_3_19_4  (
            .in0(N__13509),
            .in1(N__10954),
            .in2(N__9817),
            .in3(_gnd_net_),
            .lcout(\b2v_inst.reg_anterior_i_4 ),
            .ltout(),
            .carryin(\b2v_inst.valor_max_final5_1_cry_3 ),
            .carryout(\b2v_inst.valor_max_final5_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_1_cry_5_c_inv_LC_3_19_5 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_1_cry_5_c_inv_LC_3_19_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_1_cry_5_c_inv_LC_3_19_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final5_1_cry_5_c_inv_LC_3_19_5  (
            .in0(_gnd_net_),
            .in1(N__10884),
            .in2(N__9796),
            .in3(N__14658),
            .lcout(\b2v_inst.reg_anterior_i_5 ),
            .ltout(),
            .carryin(\b2v_inst.valor_max_final5_1_cry_4 ),
            .carryout(\b2v_inst.valor_max_final5_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_1_cry_6_c_inv_LC_3_19_6 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_1_cry_6_c_inv_LC_3_19_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_1_cry_6_c_inv_LC_3_19_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final5_1_cry_6_c_inv_LC_3_19_6  (
            .in0(_gnd_net_),
            .in1(N__10847),
            .in2(N__9776),
            .in3(N__14199),
            .lcout(\b2v_inst.reg_anterior_i_6 ),
            .ltout(),
            .carryin(\b2v_inst.valor_max_final5_1_cry_5 ),
            .carryout(\b2v_inst.valor_max_final5_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_1_cry_7_c_inv_LC_3_19_7 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_1_cry_7_c_inv_LC_3_19_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_1_cry_7_c_inv_LC_3_19_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final5_1_cry_7_c_inv_LC_3_19_7  (
            .in0(_gnd_net_),
            .in1(N__10802),
            .in2(N__9751),
            .in3(N__13604),
            .lcout(\b2v_inst.reg_anterior_i_7 ),
            .ltout(),
            .carryin(\b2v_inst.valor_max_final5_1_cry_6 ),
            .carryout(\b2v_inst.valor_max_final51 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_1_cry_7_c_RNIVOP62_LC_3_20_0 .C_ON=1'b0;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_1_cry_7_c_RNIVOP62_LC_3_20_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_1_cry_7_c_RNIVOP62_LC_3_20_0 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final5_1_cry_7_c_RNIVOP62_LC_3_20_0  (
            .in0(N__13229),
            .in1(N__9731),
            .in2(N__9716),
            .in3(N__9707),
            .lcout(\b2v_inst.N_264 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_2_4_LC_3_20_3 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_2_4_LC_3_20_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_2_4_LC_3_20_3 .LUT_INIT=16'b0000001000000111;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_2_4_LC_3_20_3  (
            .in0(N__13230),
            .in1(N__13514),
            .in2(N__10571),
            .in3(N__10916),
            .lcout(\b2v_inst.un1_reg_anterior_iv_0_0_2_tz_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst3.fsm_state_RNO_2_0_LC_5_10_3 .C_ON=1'b0;
    defparam \b2v_inst3.fsm_state_RNO_2_0_LC_5_10_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst3.fsm_state_RNO_2_0_LC_5_10_3 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \b2v_inst3.fsm_state_RNO_2_0_LC_5_10_3  (
            .in0(N__12157),
            .in1(N__12234),
            .in2(_gnd_net_),
            .in3(N__11600),
            .lcout(\b2v_inst3.N_434 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst3.fsm_state_RNO_0_1_LC_5_10_6 .C_ON=1'b0;
    defparam \b2v_inst3.fsm_state_RNO_0_1_LC_5_10_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst3.fsm_state_RNO_0_1_LC_5_10_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \b2v_inst3.fsm_state_RNO_0_1_LC_5_10_6  (
            .in0(N__12235),
            .in1(N__12158),
            .in2(_gnd_net_),
            .in3(N__11536),
            .lcout(),
            .ltout(\b2v_inst3.fsm_state_ns_0_0_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst3.fsm_state_1_LC_5_10_7 .C_ON=1'b0;
    defparam \b2v_inst3.fsm_state_1_LC_5_10_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst3.fsm_state_1_LC_5_10_7 .LUT_INIT=16'b0000110000001000;
    LogicCell40 \b2v_inst3.fsm_state_1_LC_5_10_7  (
            .in0(N__12159),
            .in1(N__18863),
            .in2(N__9893),
            .in3(N__13357),
            .lcout(\b2v_inst3.fsm_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22447),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst3.fsm_state_RNO_0_0_LC_5_11_0 .C_ON=1'b0;
    defparam \b2v_inst3.fsm_state_RNO_0_0_LC_5_11_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst3.fsm_state_RNO_0_0_LC_5_11_0 .LUT_INIT=16'b0000101000001010;
    LogicCell40 \b2v_inst3.fsm_state_RNO_0_0_LC_5_11_0  (
            .in0(N__12233),
            .in1(_gnd_net_),
            .in2(N__12166),
            .in3(_gnd_net_),
            .lcout(\b2v_inst3.N_490 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst3.fsm_state_RNIDA67_0_LC_5_11_1 .C_ON=1'b0;
    defparam \b2v_inst3.fsm_state_RNIDA67_0_LC_5_11_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst3.fsm_state_RNIDA67_0_LC_5_11_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \b2v_inst3.fsm_state_RNIDA67_0_LC_5_11_1  (
            .in0(_gnd_net_),
            .in1(N__12153),
            .in2(_gnd_net_),
            .in3(N__12232),
            .lcout(N_230),
            .ltout(N_230_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst3.fsm_state_RNO_1_0_LC_5_11_2 .C_ON=1'b0;
    defparam \b2v_inst3.fsm_state_RNO_1_0_LC_5_11_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst3.fsm_state_RNO_1_0_LC_5_11_2 .LUT_INIT=16'b1111111111001101;
    LogicCell40 \b2v_inst3.fsm_state_RNO_1_0_LC_5_11_2  (
            .in0(N__12265),
            .in1(N__11537),
            .in2(N__9890),
            .in3(N__9887),
            .lcout(),
            .ltout(\b2v_inst3.fsm_state_ns_i_i_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst3.fsm_state_0_LC_5_11_3 .C_ON=1'b0;
    defparam \b2v_inst3.fsm_state_0_LC_5_11_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst3.fsm_state_0_LC_5_11_3 .LUT_INIT=16'b0000001000001010;
    LogicCell40 \b2v_inst3.fsm_state_0_LC_5_11_3  (
            .in0(N__18915),
            .in1(N__9881),
            .in2(N__9875),
            .in3(N__13351),
            .lcout(\b2v_inst3.fsm_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22267),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNIAJF6_9_LC_5_11_6 .C_ON=1'b0;
    defparam \b2v_inst.state_RNIAJF6_9_LC_5_11_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNIAJF6_9_LC_5_11_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \b2v_inst.state_RNIAJF6_9_LC_5_11_6  (
            .in0(N__18914),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13970),
            .lcout(\b2v_inst.N_138_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst3.cycle_counter_6_LC_5_12_0 .C_ON=1'b0;
    defparam \b2v_inst3.cycle_counter_6_LC_5_12_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst3.cycle_counter_6_LC_5_12_0 .LUT_INIT=16'b0001010001000100;
    LogicCell40 \b2v_inst3.cycle_counter_6_LC_5_12_0  (
            .in0(N__13349),
            .in1(N__11690),
            .in2(N__9970),
            .in3(N__11672),
            .lcout(\b2v_inst3.cycle_counterZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22515),
            .ce(),
            .sr(N__22889));
    defparam \b2v_inst3.cycle_counter_7_LC_5_12_2 .C_ON=1'b0;
    defparam \b2v_inst3.cycle_counter_7_LC_5_12_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst3.cycle_counter_7_LC_5_12_2 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \b2v_inst3.cycle_counter_7_LC_5_12_2  (
            .in0(N__11653),
            .in1(N__11689),
            .in2(N__9971),
            .in3(N__11670),
            .lcout(\b2v_inst3.cycle_counterZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22515),
            .ce(),
            .sr(N__22889));
    defparam \b2v_inst3.cycle_counter_RNI4OAT_4_LC_5_12_3 .C_ON=1'b0;
    defparam \b2v_inst3.cycle_counter_RNI4OAT_4_LC_5_12_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst3.cycle_counter_RNI4OAT_4_LC_5_12_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \b2v_inst3.cycle_counter_RNI4OAT_4_LC_5_12_3  (
            .in0(N__12058),
            .in1(N__12035),
            .in2(_gnd_net_),
            .in3(N__12118),
            .lcout(),
            .ltout(\b2v_inst3.un1_m2_0_a2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst3.cycle_counter_RNIIR2O1_1_LC_5_12_4 .C_ON=1'b0;
    defparam \b2v_inst3.cycle_counter_RNIIR2O1_1_LC_5_12_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst3.cycle_counter_RNIIR2O1_1_LC_5_12_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst3.cycle_counter_RNIIR2O1_1_LC_5_12_4  (
            .in0(N__14298),
            .in1(N__12081),
            .in2(N__9974),
            .in3(N__12198),
            .lcout(\b2v_inst3.un1_cycle_counter_5_c5 ),
            .ltout(\b2v_inst3.un1_cycle_counter_5_c5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst3.cycle_counter_5_LC_5_12_5 .C_ON=1'b0;
    defparam \b2v_inst3.cycle_counter_5_LC_5_12_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst3.cycle_counter_5_LC_5_12_5 .LUT_INIT=16'b0000000001011010;
    LogicCell40 \b2v_inst3.cycle_counter_5_LC_5_12_5  (
            .in0(N__11671),
            .in1(_gnd_net_),
            .in2(N__9956),
            .in3(N__13348),
            .lcout(\b2v_inst3.cycle_counterZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22515),
            .ce(),
            .sr(N__22889));
    defparam \b2v_inst3.cycle_counter_3_LC_5_12_6 .C_ON=1'b0;
    defparam \b2v_inst3.cycle_counter_3_LC_5_12_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst3.cycle_counter_3_LC_5_12_6 .LUT_INIT=16'b0000000001101010;
    LogicCell40 \b2v_inst3.cycle_counter_3_LC_5_12_6  (
            .in0(N__12059),
            .in1(N__12095),
            .in2(N__12089),
            .in3(N__13347),
            .lcout(\b2v_inst3.cycle_counterZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22515),
            .ce(),
            .sr(N__22889));
    defparam \b2v_inst3.cycle_counter_2_LC_5_12_7 .C_ON=1'b0;
    defparam \b2v_inst3.cycle_counter_2_LC_5_12_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst3.cycle_counter_2_LC_5_12_7 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \b2v_inst3.cycle_counter_2_LC_5_12_7  (
            .in0(N__12199),
            .in1(N__14299),
            .in2(N__12088),
            .in3(N__12119),
            .lcout(\b2v_inst3.cycle_counterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22515),
            .ce(),
            .sr(N__22889));
    defparam \b2v_inst4.reg_data_0_LC_5_13_0 .C_ON=1'b0;
    defparam \b2v_inst4.reg_data_0_LC_5_13_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst4.reg_data_0_LC_5_13_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst4.reg_data_0_LC_5_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9953),
            .lcout(SYNTHESIZED_WIRE_3_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22405),
            .ce(N__10028),
            .sr(N__22893));
    defparam \b2v_inst4.reg_data_1_LC_5_13_1 .C_ON=1'b0;
    defparam \b2v_inst4.reg_data_1_LC_5_13_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst4.reg_data_1_LC_5_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst4.reg_data_1_LC_5_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15749),
            .lcout(SYNTHESIZED_WIRE_3_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22405),
            .ce(N__10028),
            .sr(N__22893));
    defparam \b2v_inst4.reg_data_2_LC_5_13_2 .C_ON=1'b0;
    defparam \b2v_inst4.reg_data_2_LC_5_13_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst4.reg_data_2_LC_5_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst4.reg_data_2_LC_5_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12350),
            .lcout(SYNTHESIZED_WIRE_3_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22405),
            .ce(N__10028),
            .sr(N__22893));
    defparam \b2v_inst4.reg_data_3_LC_5_13_3 .C_ON=1'b0;
    defparam \b2v_inst4.reg_data_3_LC_5_13_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst4.reg_data_3_LC_5_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst4.reg_data_3_LC_5_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12338),
            .lcout(SYNTHESIZED_WIRE_3_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22405),
            .ce(N__10028),
            .sr(N__22893));
    defparam \b2v_inst4.reg_data_4_LC_5_13_4 .C_ON=1'b0;
    defparam \b2v_inst4.reg_data_4_LC_5_13_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst4.reg_data_4_LC_5_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst4.reg_data_4_LC_5_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12326),
            .lcout(SYNTHESIZED_WIRE_3_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22405),
            .ce(N__10028),
            .sr(N__22893));
    defparam \b2v_inst4.reg_data_5_LC_5_13_5 .C_ON=1'b0;
    defparam \b2v_inst4.reg_data_5_LC_5_13_5 .SEQ_MODE=4'b1010;
    defparam \b2v_inst4.reg_data_5_LC_5_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst4.reg_data_5_LC_5_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12314),
            .lcout(SYNTHESIZED_WIRE_3_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22405),
            .ce(N__10028),
            .sr(N__22893));
    defparam \b2v_inst4.reg_data_6_LC_5_13_6 .C_ON=1'b0;
    defparam \b2v_inst4.reg_data_6_LC_5_13_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst4.reg_data_6_LC_5_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst4.reg_data_6_LC_5_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12301),
            .lcout(SYNTHESIZED_WIRE_3_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22405),
            .ce(N__10028),
            .sr(N__22893));
    defparam \b2v_inst4.reg_data_7_LC_5_13_7 .C_ON=1'b0;
    defparam \b2v_inst4.reg_data_7_LC_5_13_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst4.reg_data_7_LC_5_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst4.reg_data_7_LC_5_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12557),
            .lcout(SYNTHESIZED_WIRE_3_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22405),
            .ce(N__10028),
            .sr(N__22893));
    defparam \b2v_inst.state_RNINUTP_2_LC_5_14_0 .C_ON=1'b0;
    defparam \b2v_inst.state_RNINUTP_2_LC_5_14_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNINUTP_2_LC_5_14_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst.state_RNINUTP_2_LC_5_14_0  (
            .in0(N__10143),
            .in1(N__16481),
            .in2(N__14796),
            .in3(N__15234),
            .lcout(),
            .ltout(\b2v_inst.we_0_a2_0_a2_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNIJHF42_2_LC_5_14_1 .C_ON=1'b0;
    defparam \b2v_inst.state_RNIJHF42_2_LC_5_14_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNIJHF42_2_LC_5_14_1 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \b2v_inst.state_RNIJHF42_2_LC_5_14_1  (
            .in0(N__9980),
            .in1(N__16958),
            .in2(N__9995),
            .in3(N__15380),
            .lcout(SYNTHESIZED_WIRE_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNICN8L_3_LC_5_14_2 .C_ON=1'b0;
    defparam \b2v_inst.state_RNICN8L_3_LC_5_14_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNICN8L_3_LC_5_14_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst.state_RNICN8L_3_LC_5_14_2  (
            .in0(N__10182),
            .in1(N__15632),
            .in2(N__12278),
            .in3(N__18998),
            .lcout(\b2v_inst.we_0_a2_0_a2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNI3LTB_3_LC_5_14_3 .C_ON=1'b0;
    defparam \b2v_inst.state_RNI3LTB_3_LC_5_14_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNI3LTB_3_LC_5_14_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \b2v_inst.state_RNI3LTB_3_LC_5_14_3  (
            .in0(_gnd_net_),
            .in1(N__12276),
            .in2(_gnd_net_),
            .in3(N__10183),
            .lcout(N_458),
            .ltout(N_458_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_3_LC_5_14_4 .C_ON=1'b0;
    defparam \b2v_inst.state_3_LC_5_14_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.state_3_LC_5_14_4 .LUT_INIT=16'b0000111100001010;
    LogicCell40 \b2v_inst.state_3_LC_5_14_4  (
            .in0(N__12277),
            .in1(_gnd_net_),
            .in2(N__10223),
            .in3(N__14322),
            .lcout(\b2v_inst.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22517),
            .ce(),
            .sr(N__22898));
    defparam \b2v_inst.state_RNO_0_16_LC_5_14_5 .C_ON=1'b0;
    defparam \b2v_inst.state_RNO_0_16_LC_5_14_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNO_0_16_LC_5_14_5 .LUT_INIT=16'b0000000100000101;
    LogicCell40 \b2v_inst.state_RNO_0_16_LC_5_14_5  (
            .in0(N__15633),
            .in1(N__17698),
            .in2(N__10157),
            .in3(N__18774),
            .lcout(),
            .ltout(\b2v_inst.N_429_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_16_LC_5_14_6 .C_ON=1'b0;
    defparam \b2v_inst.state_16_LC_5_14_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.state_16_LC_5_14_6 .LUT_INIT=16'b0000101100001111;
    LogicCell40 \b2v_inst.state_16_LC_5_14_6  (
            .in0(N__10144),
            .in1(N__13709),
            .in2(N__10220),
            .in3(N__10217),
            .lcout(\b2v_inst.stateZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22517),
            .ce(),
            .sr(N__22898));
    defparam \b2v_inst.state_2_LC_5_14_7 .C_ON=1'b0;
    defparam \b2v_inst.state_2_LC_5_14_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.state_2_LC_5_14_7 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \b2v_inst.state_2_LC_5_14_7  (
            .in0(N__14321),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10184),
            .lcout(\b2v_inst.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22517),
            .ce(),
            .sr(N__22898));
    defparam \b2v_inst.data_a_escribir9_4_c_RNO_LC_5_15_0 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir9_4_c_RNO_LC_5_15_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir9_4_c_RNO_LC_5_15_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst.data_a_escribir9_4_c_RNO_LC_5_15_0  (
            .in0(N__11094),
            .in1(N__11121),
            .in2(N__10984),
            .in3(N__10242),
            .lcout(\b2v_inst.data_a_escribir9_4_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.reg_ancho_3_0_LC_5_15_1 .C_ON=1'b0;
    defparam \b2v_inst.reg_ancho_3_0_LC_5_15_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_ancho_3_0_LC_5_15_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \b2v_inst.reg_ancho_3_0_LC_5_15_1  (
            .in0(_gnd_net_),
            .in1(N__15594),
            .in2(_gnd_net_),
            .in3(N__13085),
            .lcout(\b2v_inst.reg_ancho_3Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22406),
            .ce(N__16045),
            .sr(N__22902));
    defparam \b2v_inst.reg_ancho_3_1_LC_5_15_2 .C_ON=1'b0;
    defparam \b2v_inst.reg_ancho_3_1_LC_5_15_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_ancho_3_1_LC_5_15_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \b2v_inst.reg_ancho_3_1_LC_5_15_2  (
            .in0(N__15595),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13010),
            .lcout(\b2v_inst.reg_ancho_3Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22406),
            .ce(N__16045),
            .sr(N__22902));
    defparam \b2v_inst.reg_ancho_3_2_LC_5_15_3 .C_ON=1'b0;
    defparam \b2v_inst.reg_ancho_3_2_LC_5_15_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_ancho_3_2_LC_5_15_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \b2v_inst.reg_ancho_3_2_LC_5_15_3  (
            .in0(_gnd_net_),
            .in1(N__15596),
            .in2(_gnd_net_),
            .in3(N__12941),
            .lcout(\b2v_inst.reg_ancho_3Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22406),
            .ce(N__16045),
            .sr(N__22902));
    defparam \b2v_inst.reg_ancho_3_3_LC_5_15_4 .C_ON=1'b0;
    defparam \b2v_inst.reg_ancho_3_3_LC_5_15_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_ancho_3_3_LC_5_15_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \b2v_inst.reg_ancho_3_3_LC_5_15_4  (
            .in0(N__15597),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12869),
            .lcout(\b2v_inst.reg_ancho_3Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22406),
            .ce(N__16045),
            .sr(N__22902));
    defparam \b2v_inst.reg_ancho_3_7_LC_5_15_5 .C_ON=1'b0;
    defparam \b2v_inst.reg_ancho_3_7_LC_5_15_5 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_ancho_3_7_LC_5_15_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \b2v_inst.reg_ancho_3_7_LC_5_15_5  (
            .in0(_gnd_net_),
            .in1(N__15599),
            .in2(_gnd_net_),
            .in3(N__13619),
            .lcout(\b2v_inst.reg_ancho_3Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22406),
            .ce(N__16045),
            .sr(N__22902));
    defparam \b2v_inst.data_a_escribir9_5_c_RNO_LC_5_15_6 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir9_5_c_RNO_LC_5_15_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir9_5_c_RNO_LC_5_15_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst.data_a_escribir9_5_c_RNO_LC_5_15_6  (
            .in0(N__12784),
            .in1(N__12808),
            .in2(N__10756),
            .in3(N__10905),
            .lcout(\b2v_inst.data_a_escribir9_5_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.reg_ancho_3_4_LC_5_15_7 .C_ON=1'b0;
    defparam \b2v_inst.reg_ancho_3_4_LC_5_15_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_ancho_3_4_LC_5_15_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \b2v_inst.reg_ancho_3_4_LC_5_15_7  (
            .in0(_gnd_net_),
            .in1(N__15598),
            .in2(_gnd_net_),
            .in3(N__13535),
            .lcout(\b2v_inst.reg_ancho_3Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22406),
            .ce(N__16045),
            .sr(N__22902));
    defparam \b2v_inst.data_a_escribir_RNO_0_6_LC_5_16_0 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_0_6_LC_5_16_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_0_6_LC_5_16_0 .LUT_INIT=16'b1111101011101110;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_0_6_LC_5_16_0  (
            .in0(N__10567),
            .in1(N__10845),
            .in2(N__11267),
            .in3(N__10701),
            .lcout(\b2v_inst.un1_m3_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_1_6_LC_5_16_2 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_1_6_LC_5_16_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_1_6_LC_5_16_2 .LUT_INIT=16'b0100010001010101;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_1_6_LC_5_16_2  (
            .in0(N__10628),
            .in1(N__14204),
            .in2(_gnd_net_),
            .in3(N__10619),
            .lcout(),
            .ltout(\b2v_inst.data_a_escribir_RNO_1Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_6_LC_5_16_3 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_6_LC_5_16_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.data_a_escribir_6_LC_5_16_3 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \b2v_inst.data_a_escribir_6_LC_5_16_3  (
            .in0(N__10589),
            .in1(N__10583),
            .in2(N__10574),
            .in3(N__10433),
            .lcout(b2v_inst_data_a_escribir_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22573),
            .ce(N__10351),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNO_2_7_LC_5_16_5 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNO_2_7_LC_5_16_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNO_2_7_LC_5_16_5 .LUT_INIT=16'b0000000100100011;
    LogicCell40 \b2v_inst.data_a_escribir_RNO_2_7_LC_5_16_5  (
            .in0(N__13233),
            .in1(N__10568),
            .in2(N__10757),
            .in3(N__13602),
            .lcout(),
            .ltout(\b2v_inst.un1_reg_anterior_iv_0_0_3_0_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_7_LC_5_16_6 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_7_LC_5_16_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.data_a_escribir_7_LC_5_16_6 .LUT_INIT=16'b0000000100100011;
    LogicCell40 \b2v_inst.data_a_escribir_7_LC_5_16_6  (
            .in0(N__10432),
            .in1(N__10376),
            .in2(N__10367),
            .in3(N__10364),
            .lcout(b2v_inst_data_a_escribir_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22573),
            .ce(N__10351),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_0_cry_0_c_inv_LC_5_17_0 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_0_cry_0_c_inv_LC_5_17_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_0_cry_0_c_inv_LC_5_17_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final5_0_cry_0_c_inv_LC_5_17_0  (
            .in0(_gnd_net_),
            .in1(N__10294),
            .in2(N__12763),
            .in3(N__10246),
            .lcout(\b2v_inst.reg_ancho_3_i_0 ),
            .ltout(),
            .carryin(bfn_5_17_0_),
            .carryout(\b2v_inst.valor_max_final5_0_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_0_cry_1_c_inv_LC_5_17_1 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_0_cry_1_c_inv_LC_5_17_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_0_cry_1_c_inv_LC_5_17_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final5_0_cry_1_c_inv_LC_5_17_1  (
            .in0(_gnd_net_),
            .in1(N__11168),
            .in2(N__12736),
            .in3(N__11125),
            .lcout(\b2v_inst.reg_ancho_3_i_1 ),
            .ltout(),
            .carryin(\b2v_inst.valor_max_final5_0_cry_0 ),
            .carryout(\b2v_inst.valor_max_final5_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_0_cry_2_c_inv_LC_5_17_2 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_0_cry_2_c_inv_LC_5_17_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_0_cry_2_c_inv_LC_5_17_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final5_0_cry_2_c_inv_LC_5_17_2  (
            .in0(N__11098),
            .in1(N__11074),
            .in2(N__12703),
            .in3(_gnd_net_),
            .lcout(\b2v_inst.reg_ancho_3_i_2 ),
            .ltout(),
            .carryin(\b2v_inst.valor_max_final5_0_cry_1 ),
            .carryout(\b2v_inst.valor_max_final5_0_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_0_cry_3_c_inv_LC_5_17_3 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_0_cry_3_c_inv_LC_5_17_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_0_cry_3_c_inv_LC_5_17_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final5_0_cry_3_c_inv_LC_5_17_3  (
            .in0(_gnd_net_),
            .in1(N__11033),
            .in2(N__12676),
            .in3(N__10980),
            .lcout(\b2v_inst.reg_ancho_3_i_3 ),
            .ltout(),
            .carryin(\b2v_inst.valor_max_final5_0_cry_2 ),
            .carryout(\b2v_inst.valor_max_final5_0_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_0_cry_4_c_inv_LC_5_17_4 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_0_cry_4_c_inv_LC_5_17_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_0_cry_4_c_inv_LC_5_17_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final5_0_cry_4_c_inv_LC_5_17_4  (
            .in0(_gnd_net_),
            .in1(N__10958),
            .in2(N__12643),
            .in3(N__10909),
            .lcout(\b2v_inst.reg_ancho_3_i_4 ),
            .ltout(),
            .carryin(\b2v_inst.valor_max_final5_0_cry_3 ),
            .carryout(\b2v_inst.valor_max_final5_0_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_0_cry_5_c_inv_LC_5_17_5 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_0_cry_5_c_inv_LC_5_17_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_0_cry_5_c_inv_LC_5_17_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final5_0_cry_5_c_inv_LC_5_17_5  (
            .in0(_gnd_net_),
            .in1(N__10886),
            .in2(N__12613),
            .in3(N__12783),
            .lcout(\b2v_inst.reg_ancho_3_i_5 ),
            .ltout(),
            .carryin(\b2v_inst.valor_max_final5_0_cry_4 ),
            .carryout(\b2v_inst.valor_max_final5_0_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_0_cry_6_c_inv_LC_5_17_6 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_0_cry_6_c_inv_LC_5_17_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_0_cry_6_c_inv_LC_5_17_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final5_0_cry_6_c_inv_LC_5_17_6  (
            .in0(_gnd_net_),
            .in1(N__10846),
            .in2(N__12583),
            .in3(N__12807),
            .lcout(\b2v_inst.reg_ancho_3_i_6 ),
            .ltout(),
            .carryin(\b2v_inst.valor_max_final5_0_cry_5 ),
            .carryout(\b2v_inst.valor_max_final5_0_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_0_cry_7_c_inv_LC_5_17_7 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_0_cry_7_c_inv_LC_5_17_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_0_cry_7_c_inv_LC_5_17_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final5_0_cry_7_c_inv_LC_5_17_7  (
            .in0(_gnd_net_),
            .in1(N__10801),
            .in2(N__13267),
            .in3(N__10752),
            .lcout(\b2v_inst.reg_ancho_3_i_7 ),
            .ltout(),
            .carryin(\b2v_inst.valor_max_final5_0_cry_6 ),
            .carryout(\b2v_inst.valor_max_final50 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.valor_max_final50_THRU_LUT4_0_LC_5_18_0 .C_ON=1'b0;
    defparam \b2v_inst.valor_max_final50_THRU_LUT4_0_LC_5_18_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.valor_max_final50_THRU_LUT4_0_LC_5_18_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.valor_max_final50_THRU_LUT4_0_LC_5_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10730),
            .lcout(\b2v_inst.valor_max_final50_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir9_6_c_RNO_LC_5_18_1 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir9_6_c_RNO_LC_5_18_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir9_6_c_RNO_LC_5_18_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst.data_a_escribir9_6_c_RNO_LC_5_18_1  (
            .in0(N__12914),
            .in1(N__12986),
            .in2(N__12847),
            .in3(N__13058),
            .lcout(\b2v_inst.data_a_escribir9_6_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_2_cry_0_c_LC_5_19_0 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_2_cry_0_c_LC_5_19_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_2_cry_0_c_LC_5_19_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final5_2_cry_0_c_LC_5_19_0  (
            .in0(_gnd_net_),
            .in1(N__11512),
            .in2(N__12767),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_19_0_),
            .carryout(\b2v_inst.valor_max_final5_2_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_2_cry_1_c_LC_5_19_1 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_2_cry_1_c_LC_5_19_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_2_cry_1_c_LC_5_19_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final5_2_cry_1_c_LC_5_19_1  (
            .in0(_gnd_net_),
            .in1(N__11474),
            .in2(N__12737),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.valor_max_final5_2_cry_0 ),
            .carryout(\b2v_inst.valor_max_final5_2_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_2_cry_2_c_LC_5_19_2 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_2_cry_2_c_LC_5_19_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_2_cry_2_c_LC_5_19_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final5_2_cry_2_c_LC_5_19_2  (
            .in0(_gnd_net_),
            .in1(N__11428),
            .in2(N__12707),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.valor_max_final5_2_cry_1 ),
            .carryout(\b2v_inst.valor_max_final5_2_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_2_cry_3_c_LC_5_19_3 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_2_cry_3_c_LC_5_19_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_2_cry_3_c_LC_5_19_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final5_2_cry_3_c_LC_5_19_3  (
            .in0(_gnd_net_),
            .in1(N__11388),
            .in2(N__12677),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.valor_max_final5_2_cry_2 ),
            .carryout(\b2v_inst.valor_max_final5_2_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_2_cry_4_c_LC_5_19_4 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_2_cry_4_c_LC_5_19_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_2_cry_4_c_LC_5_19_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final5_2_cry_4_c_LC_5_19_4  (
            .in0(_gnd_net_),
            .in1(N__11344),
            .in2(N__12647),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.valor_max_final5_2_cry_3 ),
            .carryout(\b2v_inst.valor_max_final5_2_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_2_cry_5_c_LC_5_19_5 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_2_cry_5_c_LC_5_19_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_2_cry_5_c_LC_5_19_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final5_2_cry_5_c_LC_5_19_5  (
            .in0(_gnd_net_),
            .in1(N__11309),
            .in2(N__12617),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.valor_max_final5_2_cry_4 ),
            .carryout(\b2v_inst.valor_max_final5_2_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_2_cry_6_c_LC_5_19_6 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_2_cry_6_c_LC_5_19_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_2_cry_6_c_LC_5_19_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final5_2_cry_6_c_LC_5_19_6  (
            .in0(_gnd_net_),
            .in1(N__11262),
            .in2(N__12587),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.valor_max_final5_2_cry_5 ),
            .carryout(\b2v_inst.valor_max_final5_2_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_2_cry_7_c_LC_5_19_7 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_2_cry_7_c_LC_5_19_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_valor_max_final5_2_cry_7_c_LC_5_19_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.encontrar_maximo_valor_max_final5_2_cry_7_c_LC_5_19_7  (
            .in0(_gnd_net_),
            .in1(N__11221),
            .in2(N__13271),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.valor_max_final5_2_cry_6 ),
            .carryout(\b2v_inst.valor_max_final52 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.valor_max_final52_THRU_LUT4_0_LC_5_20_0 .C_ON=1'b0;
    defparam \b2v_inst.valor_max_final52_THRU_LUT4_0_LC_5_20_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.valor_max_final52_THRU_LUT4_0_LC_5_20_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.valor_max_final52_THRU_LUT4_0_LC_5_20_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11639),
            .lcout(\b2v_inst.valor_max_final52_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst3.bit_counter_2_LC_6_10_0 .C_ON=1'b0;
    defparam \b2v_inst3.bit_counter_2_LC_6_10_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst3.bit_counter_2_LC_6_10_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst3.bit_counter_2_LC_6_10_0  (
            .in0(N__13380),
            .in1(N__11589),
            .in2(_gnd_net_),
            .in3(N__11609),
            .lcout(\b2v_inst3.bit_counterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22419),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst3.bit_counter_1_LC_6_10_1 .C_ON=1'b0;
    defparam \b2v_inst3.bit_counter_1_LC_6_10_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst3.bit_counter_1_LC_6_10_1 .LUT_INIT=16'b0000011000001100;
    LogicCell40 \b2v_inst3.bit_counter_1_LC_6_10_1  (
            .in0(N__13356),
            .in1(N__11573),
            .in2(N__13382),
            .in3(N__13304),
            .lcout(\b2v_inst3.bit_counterZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22419),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst3.bit_counter_RNIHGA63_1_LC_6_10_2 .C_ON=1'b0;
    defparam \b2v_inst3.bit_counter_RNIHGA63_1_LC_6_10_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst3.bit_counter_RNIHGA63_1_LC_6_10_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \b2v_inst3.bit_counter_RNIHGA63_1_LC_6_10_2  (
            .in0(N__11572),
            .in1(N__13302),
            .in2(_gnd_net_),
            .in3(N__13355),
            .lcout(\b2v_inst3.un1_bit_counter_3_c2 ),
            .ltout(\b2v_inst3.un1_bit_counter_3_c2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst3.bit_counter_3_LC_6_10_3 .C_ON=1'b0;
    defparam \b2v_inst3.bit_counter_3_LC_6_10_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst3.bit_counter_3_LC_6_10_3 .LUT_INIT=16'b0001010101000000;
    LogicCell40 \b2v_inst3.bit_counter_3_LC_6_10_3  (
            .in0(N__13379),
            .in1(N__11591),
            .in2(N__11603),
            .in3(N__11551),
            .lcout(\b2v_inst3.bit_counterZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22419),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst3.bit_counter_RNIUR5G1_3_LC_6_10_4 .C_ON=1'b0;
    defparam \b2v_inst3.bit_counter_RNIUR5G1_3_LC_6_10_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst3.bit_counter_RNIUR5G1_3_LC_6_10_4 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \b2v_inst3.bit_counter_RNIUR5G1_3_LC_6_10_4  (
            .in0(N__11590),
            .in1(N__11571),
            .in2(N__11552),
            .in3(N__13300),
            .lcout(\b2v_inst3.N_258 ),
            .ltout(\b2v_inst3.N_258_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst3.fsm_state_RNIEPSN1_0_LC_6_10_5 .C_ON=1'b0;
    defparam \b2v_inst3.fsm_state_RNIEPSN1_0_LC_6_10_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst3.fsm_state_RNIEPSN1_0_LC_6_10_5 .LUT_INIT=16'b0111011101111111;
    LogicCell40 \b2v_inst3.fsm_state_RNIEPSN1_0_LC_6_10_5  (
            .in0(N__18841),
            .in1(N__12161),
            .in2(N__11594),
            .in3(N__12242),
            .lcout(\b2v_inst3.fsm_state_RNIEPSN1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst3.bit_counter_RNIVT2O_1_LC_6_10_6 .C_ON=1'b0;
    defparam \b2v_inst3.bit_counter_RNIVT2O_1_LC_6_10_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst3.bit_counter_RNIVT2O_1_LC_6_10_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \b2v_inst3.bit_counter_RNIVT2O_1_LC_6_10_6  (
            .in0(_gnd_net_),
            .in1(N__11588),
            .in2(_gnd_net_),
            .in3(N__11570),
            .lcout(),
            .ltout(\b2v_inst3.N_102_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst3.bit_counter_RNIL1PJ1_3_LC_6_10_7 .C_ON=1'b0;
    defparam \b2v_inst3.bit_counter_RNIL1PJ1_3_LC_6_10_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst3.bit_counter_RNIL1PJ1_3_LC_6_10_7 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \b2v_inst3.bit_counter_RNIL1PJ1_3_LC_6_10_7  (
            .in0(N__13301),
            .in1(N__12160),
            .in2(N__11555),
            .in3(N__11550),
            .lcout(\b2v_inst3.N_436 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst3.txd_reg_LC_6_11_0 .C_ON=1'b0;
    defparam \b2v_inst3.txd_reg_LC_6_11_0 .SEQ_MODE=4'b1001;
    defparam \b2v_inst3.txd_reg_LC_6_11_0 .LUT_INIT=16'b1100110010111011;
    LogicCell40 \b2v_inst3.txd_reg_LC_6_11_0  (
            .in0(N__13427),
            .in1(N__12165),
            .in2(_gnd_net_),
            .in3(N__12241),
            .lcout(uart_tx_o),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22263),
            .ce(),
            .sr(N__22885));
    defparam \b2v_inst.state_4_LC_6_11_1 .C_ON=1'b0;
    defparam \b2v_inst.state_4_LC_6_11_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.state_4_LC_6_11_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst.state_4_LC_6_11_1  (
            .in0(_gnd_net_),
            .in1(N__15902),
            .in2(_gnd_net_),
            .in3(N__15866),
            .lcout(SYNTHESIZED_WIRE_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22263),
            .ce(),
            .sr(N__22885));
    defparam \b2v_inst.state_fast_17_LC_6_11_2 .C_ON=1'b0;
    defparam \b2v_inst.state_fast_17_LC_6_11_2 .SEQ_MODE=4'b1011;
    defparam \b2v_inst.state_fast_17_LC_6_11_2 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \b2v_inst.state_fast_17_LC_6_11_2  (
            .in0(N__15867),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15903),
            .lcout(\b2v_inst.state_fastZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22263),
            .ce(),
            .sr(N__22885));
    defparam \b2v_inst.state_13_LC_6_11_3 .C_ON=1'b0;
    defparam \b2v_inst.state_13_LC_6_11_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.state_13_LC_6_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.state_13_LC_6_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15080),
            .lcout(\b2v_inst.stateZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22263),
            .ce(),
            .sr(N__22885));
    defparam \b2v_inst4.state_0_LC_6_11_4 .C_ON=1'b0;
    defparam \b2v_inst4.state_0_LC_6_11_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst4.state_0_LC_6_11_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \b2v_inst4.state_0_LC_6_11_4  (
            .in0(_gnd_net_),
            .in1(N__11706),
            .in2(_gnd_net_),
            .in3(N__15725),
            .lcout(\b2v_inst4.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22263),
            .ce(),
            .sr(N__22885));
    defparam \b2v_inst3.cycle_counter_0_LC_6_12_0 .C_ON=1'b0;
    defparam \b2v_inst3.cycle_counter_0_LC_6_12_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst3.cycle_counter_0_LC_6_12_0 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \b2v_inst3.cycle_counter_0_LC_6_12_0  (
            .in0(N__14342),
            .in1(N__13350),
            .in2(_gnd_net_),
            .in3(N__12117),
            .lcout(\b2v_inst3.cycle_counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22514),
            .ce(),
            .sr(N__22890));
    defparam \b2v_inst3.cycle_counter_1_LC_6_12_1 .C_ON=1'b0;
    defparam \b2v_inst3.cycle_counter_1_LC_6_12_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst3.cycle_counter_1_LC_6_12_1 .LUT_INIT=16'b0101101011110000;
    LogicCell40 \b2v_inst3.cycle_counter_1_LC_6_12_1  (
            .in0(N__12116),
            .in1(_gnd_net_),
            .in2(N__12200),
            .in3(N__14343),
            .lcout(\b2v_inst3.cycle_counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22514),
            .ce(),
            .sr(N__22890));
    defparam \b2v_inst3.cycle_counter_RNIVMHJ_1_LC_6_12_2 .C_ON=1'b0;
    defparam \b2v_inst3.cycle_counter_RNIVMHJ_1_LC_6_12_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst3.cycle_counter_RNIVMHJ_1_LC_6_12_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \b2v_inst3.cycle_counter_RNIVMHJ_1_LC_6_12_2  (
            .in0(_gnd_net_),
            .in1(N__12193),
            .in2(_gnd_net_),
            .in3(N__12114),
            .lcout(\b2v_inst3.next_bit_0_a3_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst3.cycle_counter_RNII2471_7_LC_6_12_3 .C_ON=1'b0;
    defparam \b2v_inst3.cycle_counter_RNII2471_7_LC_6_12_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst3.cycle_counter_RNII2471_7_LC_6_12_3 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \b2v_inst3.cycle_counter_RNII2471_7_LC_6_12_3  (
            .in0(N__11688),
            .in1(N__11669),
            .in2(N__11654),
            .in3(N__12033),
            .lcout(),
            .ltout(\b2v_inst3.next_bit_0_a3_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst3.cycle_counter_RNIKK7E2_3_LC_6_12_4 .C_ON=1'b0;
    defparam \b2v_inst3.cycle_counter_RNIKK7E2_3_LC_6_12_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst3.cycle_counter_RNIKK7E2_3_LC_6_12_4 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \b2v_inst3.cycle_counter_RNIKK7E2_3_LC_6_12_4  (
            .in0(N__12056),
            .in1(N__12079),
            .in2(N__12287),
            .in3(N__12284),
            .lcout(\b2v_inst3.N_105_7 ),
            .ltout(\b2v_inst3.N_105_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst3.fsm_state_RNI3QCR2_0_LC_6_12_5 .C_ON=1'b0;
    defparam \b2v_inst3.fsm_state_RNI3QCR2_0_LC_6_12_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst3.fsm_state_RNI3QCR2_0_LC_6_12_5 .LUT_INIT=16'b0000000011100010;
    LogicCell40 \b2v_inst3.fsm_state_RNI3QCR2_0_LC_6_12_5  (
            .in0(N__12264),
            .in1(N__12172),
            .in2(N__12245),
            .in3(N__12236),
            .lcout(\b2v_inst3.un2_n_fsm_state_0_sqmuxa_2_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst3.cycle_counter_RNIC1OQ_1_LC_6_12_6 .C_ON=1'b0;
    defparam \b2v_inst3.cycle_counter_RNIC1OQ_1_LC_6_12_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst3.cycle_counter_RNIC1OQ_1_LC_6_12_6 .LUT_INIT=16'b1100100000000000;
    LogicCell40 \b2v_inst3.cycle_counter_RNIC1OQ_1_LC_6_12_6  (
            .in0(N__12237),
            .in1(N__12194),
            .in2(N__12176),
            .in3(N__12115),
            .lcout(\b2v_inst3.un1_cycle_counter_5_c2 ),
            .ltout(\b2v_inst3.un1_cycle_counter_5_c2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst3.cycle_counter_4_LC_6_12_7 .C_ON=1'b0;
    defparam \b2v_inst3.cycle_counter_4_LC_6_12_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst3.cycle_counter_4_LC_6_12_7 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \b2v_inst3.cycle_counter_4_LC_6_12_7  (
            .in0(N__12080),
            .in1(N__12057),
            .in2(N__12038),
            .in3(N__12034),
            .lcout(\b2v_inst3.cycle_counterZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22514),
            .ce(),
            .sr(N__22890));
    defparam \b2v_inst4.pix_count_int_9_LC_6_13_0 .C_ON=1'b0;
    defparam \b2v_inst4.pix_count_int_9_LC_6_13_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst4.pix_count_int_9_LC_6_13_0 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \b2v_inst4.pix_count_int_9_LC_6_13_0  (
            .in0(N__12020),
            .in1(N__11984),
            .in2(N__11948),
            .in3(N__11882),
            .lcout(SYNTHESIZED_WIRE_2_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22230),
            .ce(),
            .sr(N__22894));
    defparam \b2v_inst.cuenta_RNIQI4F_2_LC_6_13_1 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_RNIQI4F_2_LC_6_13_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.cuenta_RNIQI4F_2_LC_6_13_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \b2v_inst.cuenta_RNIQI4F_2_LC_6_13_1  (
            .in0(N__13757),
            .in1(N__13670),
            .in2(_gnd_net_),
            .in3(N__13804),
            .lcout(\b2v_inst.cuenta_RNIQI4FZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.cuenta_RNIR03A_1_LC_6_13_2 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_RNIR03A_1_LC_6_13_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.cuenta_RNIR03A_1_LC_6_13_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \b2v_inst.cuenta_RNIR03A_1_LC_6_13_2  (
            .in0(_gnd_net_),
            .in1(N__13803),
            .in2(_gnd_net_),
            .in3(N__13758),
            .lcout(\b2v_inst.cuenta_RNIR03AZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.cuenta_pixel_RNI1NM11_6_LC_6_13_3 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_pixel_RNI1NM11_6_LC_6_13_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.cuenta_pixel_RNI1NM11_6_LC_6_13_3 .LUT_INIT=16'b1111010111111111;
    LogicCell40 \b2v_inst.cuenta_pixel_RNI1NM11_6_LC_6_13_3  (
            .in0(N__12500),
            .in1(_gnd_net_),
            .in2(N__12452),
            .in3(N__11844),
            .lcout(\b2v_inst.un11_cuenta_pixel_i_0_o2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.cuenta_pixel_RNO_0_6_LC_6_13_4 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_pixel_RNO_0_6_LC_6_13_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.cuenta_pixel_RNO_0_6_LC_6_13_4 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \b2v_inst.cuenta_pixel_RNO_0_6_LC_6_13_4  (
            .in0(N__11768),
            .in1(N__12499),
            .in2(_gnd_net_),
            .in3(N__12448),
            .lcout(\b2v_inst.cuenta_pixel_4_i_a2_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNI95JL_3_LC_6_13_5 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNI95JL_3_LC_6_13_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNI95JL_3_LC_6_13_5 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \b2v_inst.data_a_escribir_RNI95JL_3_LC_6_13_5  (
            .in0(N__14549),
            .in1(N__17666),
            .in2(_gnd_net_),
            .in3(N__17018),
            .lcout(N_213_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNIB7JL_5_LC_6_13_6 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNIB7JL_5_LC_6_13_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNIB7JL_5_LC_6_13_6 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \b2v_inst.data_a_escribir_RNIB7JL_5_LC_6_13_6  (
            .in0(N__17019),
            .in1(N__14489),
            .in2(_gnd_net_),
            .in3(N__17668),
            .lcout(N_209_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNIC8JL_6_LC_6_13_7 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNIC8JL_6_LC_6_13_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNIC8JL_6_LC_6_13_7 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \b2v_inst.data_a_escribir_RNIC8JL_6_LC_6_13_7  (
            .in0(N__14456),
            .in1(N__17667),
            .in2(_gnd_net_),
            .in3(N__17020),
            .lcout(N_207_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNIJV55_11_LC_6_14_0 .C_ON=1'b0;
    defparam \b2v_inst.state_RNIJV55_11_LC_6_14_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNIJV55_11_LC_6_14_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst.state_RNIJV55_11_LC_6_14_0  (
            .in0(_gnd_net_),
            .in1(N__18937),
            .in2(_gnd_net_),
            .in3(N__14094),
            .lcout(\b2v_inst.N_136_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_RX_Byte_2_LC_6_14_2 .C_ON=1'b0;
    defparam \b2v_inst1.r_RX_Byte_2_LC_6_14_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst1.r_RX_Byte_2_LC_6_14_2 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \b2v_inst1.r_RX_Byte_2_LC_6_14_2  (
            .in0(N__17189),
            .in1(N__12349),
            .in2(N__22746),
            .in3(N__17171),
            .lcout(SYNTHESIZED_WIRE_10_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22516),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_RX_Byte_3_LC_6_14_3 .C_ON=1'b0;
    defparam \b2v_inst1.r_RX_Byte_3_LC_6_14_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst1.r_RX_Byte_3_LC_6_14_3 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \b2v_inst1.r_RX_Byte_3_LC_6_14_3  (
            .in0(N__17172),
            .in1(N__12337),
            .in2(N__22748),
            .in3(N__14573),
            .lcout(SYNTHESIZED_WIRE_10_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22516),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_RX_Byte_4_LC_6_14_4 .C_ON=1'b0;
    defparam \b2v_inst1.r_RX_Byte_4_LC_6_14_4 .SEQ_MODE=4'b1000;
    defparam \b2v_inst1.r_RX_Byte_4_LC_6_14_4 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \b2v_inst1.r_RX_Byte_4_LC_6_14_4  (
            .in0(N__14561),
            .in1(N__12325),
            .in2(N__22747),
            .in3(N__17173),
            .lcout(SYNTHESIZED_WIRE_10_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22516),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_RX_Byte_5_LC_6_14_5 .C_ON=1'b0;
    defparam \b2v_inst1.r_RX_Byte_5_LC_6_14_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst1.r_RX_Byte_5_LC_6_14_5 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \b2v_inst1.r_RX_Byte_5_LC_6_14_5  (
            .in0(N__17174),
            .in1(N__12313),
            .in2(N__22749),
            .in3(N__15251),
            .lcout(SYNTHESIZED_WIRE_10_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22516),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_RX_Byte_6_LC_6_14_6 .C_ON=1'b0;
    defparam \b2v_inst1.r_RX_Byte_6_LC_6_14_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst1.r_RX_Byte_6_LC_6_14_6 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \b2v_inst1.r_RX_Byte_6_LC_6_14_6  (
            .in0(N__13115),
            .in1(N__22733),
            .in2(N__12302),
            .in3(N__17175),
            .lcout(SYNTHESIZED_WIRE_10_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22516),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_RX_Byte_7_LC_6_14_7 .C_ON=1'b0;
    defparam \b2v_inst1.r_RX_Byte_7_LC_6_14_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst1.r_RX_Byte_7_LC_6_14_7 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \b2v_inst1.r_RX_Byte_7_LC_6_14_7  (
            .in0(N__17176),
            .in1(N__12556),
            .in2(N__22750),
            .in3(N__18278),
            .lcout(SYNTHESIZED_WIRE_10_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22516),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_3_RNIGC1F1_5_LC_6_15_0 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_3_RNIGC1F1_5_LC_6_15_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_3_RNIGC1F1_5_LC_6_15_0 .LUT_INIT=16'b1111110111011101;
    LogicCell40 \b2v_inst.dir_mem_3_RNIGC1F1_5_LC_6_15_0  (
            .in0(N__15146),
            .in1(N__12509),
            .in2(N__14150),
            .in3(N__16951),
            .lcout(),
            .ltout(\b2v_inst.addr_ram_1_iv_i_2_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_RNIBUK83_5_LC_6_15_1 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_RNIBUK83_5_LC_6_15_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNIBUK83_5_LC_6_15_1 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \b2v_inst.dir_mem_RNIBUK83_5_LC_6_15_1  (
            .in0(N__16409),
            .in1(N__12515),
            .in2(N__12545),
            .in3(N__19264),
            .lcout(N_54),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_1_RNI1SAQ_5_LC_6_15_2 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_1_RNI1SAQ_5_LC_6_15_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_1_RNI1SAQ_5_LC_6_15_2 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \b2v_inst.dir_mem_1_RNI1SAQ_5_LC_6_15_2  (
            .in0(N__19979),
            .in1(N__16473),
            .in2(N__16697),
            .in3(N__15375),
            .lcout(\b2v_inst.addr_ram_1_iv_i_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNILLMH_6_LC_6_15_3 .C_ON=1'b0;
    defparam \b2v_inst.state_RNILLMH_6_LC_6_15_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNILLMH_6_LC_6_15_3 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \b2v_inst.state_RNILLMH_6_LC_6_15_3  (
            .in0(N__15181),
            .in1(N__15846),
            .in2(_gnd_net_),
            .in3(N__20478),
            .lcout(\b2v_inst.N_341 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_5_LC_6_15_4 .C_ON=1'b0;
    defparam \b2v_inst.state_5_LC_6_15_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.state_5_LC_6_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.state_5_LC_6_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15183),
            .lcout(\b2v_inst.stateZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22454),
            .ce(),
            .sr(N__22903));
    defparam \b2v_inst.state_RNI7PTB_6_LC_6_15_5 .C_ON=1'b0;
    defparam \b2v_inst.state_RNI7PTB_6_LC_6_15_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNI7PTB_6_LC_6_15_5 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \b2v_inst.state_RNI7PTB_6_LC_6_15_5  (
            .in0(N__15180),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15844),
            .lcout(\b2v_inst.N_238 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNIEG2F_6_LC_6_15_6 .C_ON=1'b0;
    defparam \b2v_inst.state_RNIEG2F_6_LC_6_15_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNIEG2F_6_LC_6_15_6 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \b2v_inst.state_RNIEG2F_6_LC_6_15_6  (
            .in0(N__15845),
            .in1(N__15182),
            .in2(_gnd_net_),
            .in3(N__17882),
            .lcout(),
            .ltout(\b2v_inst.N_404_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_3_RNI42DC1_0_LC_6_15_7 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_3_RNI42DC1_0_LC_6_15_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_3_RNI42DC1_0_LC_6_15_7 .LUT_INIT=16'b1111100011111111;
    LogicCell40 \b2v_inst.dir_mem_3_RNI42DC1_0_LC_6_15_7  (
            .in0(N__16950),
            .in1(N__14156),
            .in2(N__12503),
            .in3(N__15145),
            .lcout(\b2v_inst.addr_ram_1_iv_i_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.reg_ancho_3_6_LC_6_16_0 .C_ON=1'b0;
    defparam \b2v_inst.reg_ancho_3_6_LC_6_16_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_ancho_3_6_LC_6_16_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \b2v_inst.reg_ancho_3_6_LC_6_16_0  (
            .in0(N__15577),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14231),
            .lcout(\b2v_inst.reg_ancho_3Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22572),
            .ce(N__16046),
            .sr(N__22908));
    defparam \b2v_inst.reg_ancho_3_5_LC_6_16_1 .C_ON=1'b0;
    defparam \b2v_inst.reg_ancho_3_5_LC_6_16_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_ancho_3_5_LC_6_16_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \b2v_inst.reg_ancho_3_5_LC_6_16_1  (
            .in0(_gnd_net_),
            .in1(N__14694),
            .in2(_gnd_net_),
            .in3(N__15576),
            .lcout(\b2v_inst.reg_ancho_3Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22572),
            .ce(N__16046),
            .sr(N__22908));
    defparam \b2v_inst.encontrar_maximo_un3_valor_max2_cry_0_c_LC_6_17_0 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_un3_valor_max2_cry_0_c_LC_6_17_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_un3_valor_max2_cry_0_c_LC_6_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.encontrar_maximo_un3_valor_max2_cry_0_c_LC_6_17_0  (
            .in0(_gnd_net_),
            .in1(N__13060),
            .in2(N__12762),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_17_0_),
            .carryout(\b2v_inst.un3_valor_max2_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_un3_valor_max2_cry_1_c_LC_6_17_1 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_un3_valor_max2_cry_1_c_LC_6_17_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_un3_valor_max2_cry_1_c_LC_6_17_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.encontrar_maximo_un3_valor_max2_cry_1_c_LC_6_17_1  (
            .in0(_gnd_net_),
            .in1(N__12991),
            .in2(N__12735),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.un3_valor_max2_cry_0 ),
            .carryout(\b2v_inst.un3_valor_max2_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_un3_valor_max2_cry_2_c_LC_6_17_2 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_un3_valor_max2_cry_2_c_LC_6_17_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_un3_valor_max2_cry_2_c_LC_6_17_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.encontrar_maximo_un3_valor_max2_cry_2_c_LC_6_17_2  (
            .in0(_gnd_net_),
            .in1(N__12919),
            .in2(N__12702),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.un3_valor_max2_cry_1 ),
            .carryout(\b2v_inst.un3_valor_max2_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_un3_valor_max2_cry_3_c_LC_6_17_3 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_un3_valor_max2_cry_3_c_LC_6_17_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_un3_valor_max2_cry_3_c_LC_6_17_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.encontrar_maximo_un3_valor_max2_cry_3_c_LC_6_17_3  (
            .in0(_gnd_net_),
            .in1(N__12846),
            .in2(N__12675),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.un3_valor_max2_cry_2 ),
            .carryout(\b2v_inst.un3_valor_max2_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_un3_valor_max2_cry_4_c_LC_6_17_4 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_un3_valor_max2_cry_4_c_LC_6_17_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_un3_valor_max2_cry_4_c_LC_6_17_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.encontrar_maximo_un3_valor_max2_cry_4_c_LC_6_17_4  (
            .in0(_gnd_net_),
            .in1(N__13513),
            .in2(N__12642),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.un3_valor_max2_cry_3 ),
            .carryout(\b2v_inst.un3_valor_max2_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_un3_valor_max2_cry_5_c_LC_6_17_5 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_un3_valor_max2_cry_5_c_LC_6_17_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_un3_valor_max2_cry_5_c_LC_6_17_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.encontrar_maximo_un3_valor_max2_cry_5_c_LC_6_17_5  (
            .in0(_gnd_net_),
            .in1(N__14659),
            .in2(N__12612),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.un3_valor_max2_cry_4 ),
            .carryout(\b2v_inst.un3_valor_max2_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_un3_valor_max2_cry_6_c_LC_6_17_6 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_un3_valor_max2_cry_6_c_LC_6_17_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_un3_valor_max2_cry_6_c_LC_6_17_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.encontrar_maximo_un3_valor_max2_cry_6_c_LC_6_17_6  (
            .in0(_gnd_net_),
            .in1(N__14200),
            .in2(N__12582),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.un3_valor_max2_cry_5 ),
            .carryout(\b2v_inst.un3_valor_max2_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.encontrar_maximo_un3_valor_max2_cry_7_c_LC_6_17_7 .C_ON=1'b1;
    defparam \b2v_inst.encontrar_maximo_un3_valor_max2_cry_7_c_LC_6_17_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.encontrar_maximo_un3_valor_max2_cry_7_c_LC_6_17_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.encontrar_maximo_un3_valor_max2_cry_7_c_LC_6_17_7  (
            .in0(_gnd_net_),
            .in1(N__13601),
            .in2(N__13266),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst.un3_valor_max2_cry_6 ),
            .carryout(\b2v_inst.un3_valor_max2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.un3_valor_max2_THRU_LUT4_0_LC_6_18_0 .C_ON=1'b0;
    defparam \b2v_inst.un3_valor_max2_THRU_LUT4_0_LC_6_18_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.un3_valor_max2_THRU_LUT4_0_LC_6_18_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.un3_valor_max2_THRU_LUT4_0_LC_6_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13241),
            .lcout(\b2v_inst.un3_valor_max2_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst3.fsm_state_RNI6DTR2_0_LC_6_18_3 .C_ON=1'b0;
    defparam \b2v_inst3.fsm_state_RNI6DTR2_0_LC_6_18_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst3.fsm_state_RNI6DTR2_0_LC_6_18_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \b2v_inst3.fsm_state_RNI6DTR2_0_LC_6_18_3  (
            .in0(_gnd_net_),
            .in1(N__13141),
            .in2(_gnd_net_),
            .in3(N__13127),
            .lcout(\b2v_inst3.un2_n_fsm_state_0_sqmuxa_2_0_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_RX_Byte_RNO_0_6_LC_6_18_5 .C_ON=1'b0;
    defparam \b2v_inst1.r_RX_Byte_RNO_0_6_LC_6_18_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_RX_Byte_RNO_0_6_LC_6_18_5 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \b2v_inst1.r_RX_Byte_RNO_0_6_LC_6_18_5  (
            .in0(N__18260),
            .in1(N__18184),
            .in2(_gnd_net_),
            .in3(N__18125),
            .lcout(\b2v_inst1.r_RX_Bytece_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.reg_anterior_0_LC_6_19_1 .C_ON=1'b0;
    defparam \b2v_inst.reg_anterior_0_LC_6_19_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_anterior_0_LC_6_19_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \b2v_inst.reg_anterior_0_LC_6_19_1  (
            .in0(_gnd_net_),
            .in1(N__15559),
            .in2(_gnd_net_),
            .in3(N__13102),
            .lcout(\b2v_inst.reg_anteriorZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22244),
            .ce(N__15239),
            .sr(N__22914));
    defparam \b2v_inst.reg_anterior_1_LC_6_19_2 .C_ON=1'b0;
    defparam \b2v_inst.reg_anterior_1_LC_6_19_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_anterior_1_LC_6_19_2 .LUT_INIT=16'b0000101000001010;
    LogicCell40 \b2v_inst.reg_anterior_1_LC_6_19_2  (
            .in0(N__13027),
            .in1(_gnd_net_),
            .in2(N__15575),
            .in3(_gnd_net_),
            .lcout(\b2v_inst.reg_anteriorZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22244),
            .ce(N__15239),
            .sr(N__22914));
    defparam \b2v_inst.reg_anterior_2_LC_6_19_3 .C_ON=1'b0;
    defparam \b2v_inst.reg_anterior_2_LC_6_19_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_anterior_2_LC_6_19_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \b2v_inst.reg_anterior_2_LC_6_19_3  (
            .in0(_gnd_net_),
            .in1(N__15563),
            .in2(_gnd_net_),
            .in3(N__12958),
            .lcout(\b2v_inst.reg_anteriorZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22244),
            .ce(N__15239),
            .sr(N__22914));
    defparam \b2v_inst.reg_anterior_3_LC_6_19_4 .C_ON=1'b0;
    defparam \b2v_inst.reg_anterior_3_LC_6_19_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_anterior_3_LC_6_19_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \b2v_inst.reg_anterior_3_LC_6_19_4  (
            .in0(N__15564),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12886),
            .lcout(\b2v_inst.reg_anteriorZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22244),
            .ce(N__15239),
            .sr(N__22914));
    defparam \b2v_inst.reg_anterior_7_LC_6_19_5 .C_ON=1'b0;
    defparam \b2v_inst.reg_anterior_7_LC_6_19_5 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_anterior_7_LC_6_19_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \b2v_inst.reg_anterior_7_LC_6_19_5  (
            .in0(_gnd_net_),
            .in1(N__15566),
            .in2(_gnd_net_),
            .in3(N__13643),
            .lcout(\b2v_inst.reg_anteriorZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22244),
            .ce(N__15239),
            .sr(N__22914));
    defparam \b2v_inst.data_a_escribir9_7_c_RNO_LC_6_19_6 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir9_7_c_RNO_LC_6_19_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir9_7_c_RNO_LC_6_19_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst.data_a_escribir9_7_c_RNO_LC_6_19_6  (
            .in0(N__14198),
            .in1(N__14648),
            .in2(N__13603),
            .in3(N__13508),
            .lcout(\b2v_inst.data_a_escribir9_7_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.reg_anterior_4_LC_6_19_7 .C_ON=1'b0;
    defparam \b2v_inst.reg_anterior_4_LC_6_19_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_anterior_4_LC_6_19_7 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \b2v_inst.reg_anterior_4_LC_6_19_7  (
            .in0(N__13552),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15565),
            .lcout(\b2v_inst.reg_anteriorZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22244),
            .ce(N__15239),
            .sr(N__22914));
    defparam \b2v_inst3.data_to_send_esr_1_LC_6_20_2 .C_ON=1'b0;
    defparam \b2v_inst3.data_to_send_esr_1_LC_6_20_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst3.data_to_send_esr_1_LC_6_20_2 .LUT_INIT=16'b1111000000100010;
    LogicCell40 \b2v_inst3.data_to_send_esr_1_LC_6_20_2  (
            .in0(N__13481),
            .in1(N__14419),
            .in2(N__13391),
            .in3(N__14341),
            .lcout(\b2v_inst3.data_to_sendZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22571),
            .ce(N__14258),
            .sr(N__22918));
    defparam \b2v_inst3.data_to_send_esr_0_LC_6_20_4 .C_ON=1'b0;
    defparam \b2v_inst3.data_to_send_esr_0_LC_6_20_4 .SEQ_MODE=4'b1000;
    defparam \b2v_inst3.data_to_send_esr_0_LC_6_20_4 .LUT_INIT=16'b1111000000100010;
    LogicCell40 \b2v_inst3.data_to_send_esr_0_LC_6_20_4  (
            .in0(N__13460),
            .in1(N__14418),
            .in2(N__13436),
            .in3(N__14340),
            .lcout(\b2v_inst3.data_to_sendZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22571),
            .ce(N__14258),
            .sr(N__22918));
    defparam \b2v_inst3.data_to_send_esr_2_LC_6_20_5 .C_ON=1'b0;
    defparam \b2v_inst3.data_to_send_esr_2_LC_6_20_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst3.data_to_send_esr_2_LC_6_20_5 .LUT_INIT=16'b1000100011011000;
    LogicCell40 \b2v_inst3.data_to_send_esr_2_LC_6_20_5  (
            .in0(N__14339),
            .in1(N__14525),
            .in2(N__13415),
            .in3(N__14420),
            .lcout(\b2v_inst3.data_to_sendZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22571),
            .ce(N__14258),
            .sr(N__22918));
    defparam \b2v_inst3.bit_counter_0_LC_7_10_3 .C_ON=1'b0;
    defparam \b2v_inst3.bit_counter_0_LC_7_10_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst3.bit_counter_0_LC_7_10_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst3.bit_counter_0_LC_7_10_3  (
            .in0(N__13381),
            .in1(N__13303),
            .in2(_gnd_net_),
            .in3(N__13358),
            .lcout(\b2v_inst3.bit_counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22083),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.cuenta_RNIFIIS1_4_LC_7_11_0 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_RNIFIIS1_4_LC_7_11_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.cuenta_RNIFIIS1_4_LC_7_11_0 .LUT_INIT=16'b1011001111101100;
    LogicCell40 \b2v_inst.cuenta_RNIFIIS1_4_LC_7_11_0  (
            .in0(N__13852),
            .in1(N__15020),
            .in2(N__13280),
            .in3(N__14988),
            .lcout(\b2v_inst.state_ns_a2_0_o2_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.cuenta_RNIQI4F_0_2_LC_7_11_1 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_RNIQI4F_0_2_LC_7_11_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.cuenta_RNIQI4F_0_2_LC_7_11_1 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \b2v_inst.cuenta_RNIQI4F_0_2_LC_7_11_1  (
            .in0(N__13668),
            .in1(N__13801),
            .in2(_gnd_net_),
            .in3(N__13743),
            .lcout(\b2v_inst.state_ns_a2_0_a2_0_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.cuenta_RNIQ56K_0_3_LC_7_11_2 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_RNIQ56K_0_3_LC_7_11_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.cuenta_RNIQ56K_0_3_LC_7_11_2 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \b2v_inst.cuenta_RNIQ56K_0_3_LC_7_11_2  (
            .in0(N__13742),
            .in1(N__13666),
            .in2(N__13805),
            .in3(N__13686),
            .lcout(\b2v_inst.cuenta_RNIQ56K_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.cuenta_RNO_0_0_LC_7_11_3 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_RNO_0_0_LC_7_11_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.cuenta_RNO_0_0_LC_7_11_3 .LUT_INIT=16'b1011111100110011;
    LogicCell40 \b2v_inst.cuenta_RNO_0_0_LC_7_11_3  (
            .in0(N__18707),
            .in1(N__13745),
            .in2(N__17700),
            .in3(N__14606),
            .lcout(),
            .ltout(\b2v_inst.cuenta_5_i_a2_2_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.cuenta_0_LC_7_11_4 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_0_LC_7_11_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.cuenta_0_LC_7_11_4 .LUT_INIT=16'b1111101011111000;
    LogicCell40 \b2v_inst.cuenta_0_LC_7_11_4  (
            .in0(N__14859),
            .in1(N__16217),
            .in2(N__13694),
            .in3(N__16168),
            .lcout(\b2v_inst.cuentaZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21947),
            .ce(N__14905),
            .sr(N__22891));
    defparam \b2v_inst.cuenta_RNIQ56K_3_LC_7_11_5 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_RNIQ56K_3_LC_7_11_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.cuenta_RNIQ56K_3_LC_7_11_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst.cuenta_RNIQ56K_3_LC_7_11_5  (
            .in0(N__13665),
            .in1(N__13796),
            .in2(N__13688),
            .in3(N__13741),
            .lcout(\b2v_inst.un4_cuenta_c4 ),
            .ltout(\b2v_inst.un4_cuenta_c4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.cuenta_4_LC_7_11_6 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_4_LC_7_11_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.cuenta_4_LC_7_11_6 .LUT_INIT=16'b0000000000101000;
    LogicCell40 \b2v_inst.cuenta_4_LC_7_11_6  (
            .in0(N__17683),
            .in1(N__15021),
            .in2(N__13691),
            .in3(N__18708),
            .lcout(\b2v_inst.cuentaZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21947),
            .ce(N__14905),
            .sr(N__22891));
    defparam \b2v_inst.cuenta_RNO_1_3_LC_7_11_7 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_RNO_1_3_LC_7_11_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.cuenta_RNO_1_3_LC_7_11_7 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst.cuenta_RNO_1_3_LC_7_11_7  (
            .in0(N__13667),
            .in1(N__13800),
            .in2(_gnd_net_),
            .in3(N__13744),
            .lcout(\b2v_inst.cuenta_5_i_a2_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.cuenta_3_LC_7_12_0 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_3_LC_7_12_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.cuenta_3_LC_7_12_0 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \b2v_inst.cuenta_3_LC_7_12_0  (
            .in0(N__13853),
            .in1(N__13718),
            .in2(_gnd_net_),
            .in3(N__14585),
            .lcout(\b2v_inst.cuentaZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22084),
            .ce(N__14898),
            .sr(N__22895));
    defparam \b2v_inst.cuenta_2_LC_7_12_1 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_2_LC_7_12_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.cuenta_2_LC_7_12_1 .LUT_INIT=16'b0000010001000100;
    LogicCell40 \b2v_inst.cuenta_2_LC_7_12_1  (
            .in0(N__14584),
            .in1(N__13829),
            .in2(N__13820),
            .in3(N__13835),
            .lcout(\b2v_inst.cuentaZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22084),
            .ce(N__14898),
            .sr(N__22895));
    defparam \b2v_inst.cuenta_fast_RNIBDJQ_4_LC_7_12_2 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_fast_RNIBDJQ_4_LC_7_12_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.cuenta_fast_RNIBDJQ_4_LC_7_12_2 .LUT_INIT=16'b1010000010000000;
    LogicCell40 \b2v_inst.cuenta_fast_RNIBDJQ_4_LC_7_12_2  (
            .in0(N__13687),
            .in1(N__13669),
            .in2(N__13868),
            .in3(N__13802),
            .lcout(\b2v_inst.un2_cuentalto7_3 ),
            .ltout(\b2v_inst.un2_cuentalto7_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.cuenta_RNIKFO91_7_LC_7_12_3 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_RNIKFO91_7_LC_7_12_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.cuenta_RNIKFO91_7_LC_7_12_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst.cuenta_RNIKFO91_7_LC_7_12_3  (
            .in0(N__14925),
            .in1(N__14953),
            .in2(N__13874),
            .in3(N__15058),
            .lcout(\b2v_inst.N_351_0 ),
            .ltout(\b2v_inst.N_351_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.cuenta_fast_4_LC_7_12_4 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_fast_4_LC_7_12_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.cuenta_fast_4_LC_7_12_4 .LUT_INIT=16'b0000001000001000;
    LogicCell40 \b2v_inst.cuenta_fast_4_LC_7_12_4  (
            .in0(N__17669),
            .in1(N__13867),
            .in2(N__13871),
            .in3(N__14989),
            .lcout(\b2v_inst.cuenta_fastZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22084),
            .ce(N__14898),
            .sr(N__22895));
    defparam \b2v_inst.cuenta_RNI1OL72_0_LC_7_12_5 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_RNI1OL72_0_LC_7_12_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.cuenta_RNI1OL72_0_LC_7_12_5 .LUT_INIT=16'b0000000010001010;
    LogicCell40 \b2v_inst.cuenta_RNI1OL72_0_LC_7_12_5  (
            .in0(N__13851),
            .in1(N__18709),
            .in2(N__17701),
            .in3(N__13760),
            .lcout(\b2v_inst.N_376_1 ),
            .ltout(\b2v_inst.N_376_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.cuenta_1_LC_7_12_6 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_1_LC_7_12_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.cuenta_1_LC_7_12_6 .LUT_INIT=16'b0000000001001100;
    LogicCell40 \b2v_inst.cuenta_1_LC_7_12_6  (
            .in0(N__13828),
            .in1(N__13816),
            .in2(N__13808),
            .in3(N__14583),
            .lcout(\b2v_inst.cuentaZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22084),
            .ce(N__14898),
            .sr(N__22895));
    defparam \b2v_inst.cuenta_RNO_0_3_LC_7_13_0 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_RNO_0_3_LC_7_13_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.cuenta_RNO_0_3_LC_7_13_0 .LUT_INIT=16'b0000000010001010;
    LogicCell40 \b2v_inst.cuenta_RNO_0_3_LC_7_13_0  (
            .in0(N__13769),
            .in1(N__18703),
            .in2(N__17692),
            .in3(N__13759),
            .lcout(\b2v_inst.N_377 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNIP7VJ_10_LC_7_13_1 .C_ON=1'b0;
    defparam \b2v_inst.state_RNIP7VJ_10_LC_7_13_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNIP7VJ_10_LC_7_13_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst.state_RNIP7VJ_10_LC_7_13_1  (
            .in0(N__13892),
            .in1(N__15477),
            .in2(N__15224),
            .in3(N__16024),
            .lcout(\b2v_inst.N_491 ),
            .ltout(\b2v_inst.N_491_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNIFQKO_17_LC_7_13_2 .C_ON=1'b0;
    defparam \b2v_inst.state_RNIFQKO_17_LC_7_13_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNIFQKO_17_LC_7_13_2 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \b2v_inst.state_RNIFQKO_17_LC_7_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13712),
            .in3(N__17639),
            .lcout(\b2v_inst.state_RNIFQKOZ0Z_17 ),
            .ltout(\b2v_inst.state_RNIFQKOZ0Z_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNIFQKO_0_17_LC_7_13_3 .C_ON=1'b0;
    defparam \b2v_inst.state_RNIFQKO_0_17_LC_7_13_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNIFQKO_0_17_LC_7_13_3 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \b2v_inst.state_RNIFQKO_0_17_LC_7_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13697),
            .in3(_gnd_net_),
            .lcout(\b2v_inst.N_399_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNIDVTB_9_LC_7_13_4 .C_ON=1'b0;
    defparam \b2v_inst.state_RNIDVTB_9_LC_7_13_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNIDVTB_9_LC_7_13_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \b2v_inst.state_RNIDVTB_9_LC_7_13_4  (
            .in0(_gnd_net_),
            .in1(N__16023),
            .in2(_gnd_net_),
            .in3(N__13962),
            .lcout(\b2v_inst.N_236 ),
            .ltout(\b2v_inst.N_236_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_8_LC_7_13_5 .C_ON=1'b0;
    defparam \b2v_inst.state_8_LC_7_13_5 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.state_8_LC_7_13_5 .LUT_INIT=16'b1010000010110000;
    LogicCell40 \b2v_inst.state_8_LC_7_13_5  (
            .in0(N__13963),
            .in1(N__16077),
            .in2(N__13973),
            .in3(N__14824),
            .lcout(\b2v_inst.stateZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22554),
            .ce(),
            .sr(N__22899));
    defparam \b2v_inst.state_17_LC_7_13_6 .C_ON=1'b0;
    defparam \b2v_inst.state_17_LC_7_13_6 .SEQ_MODE=4'b1011;
    defparam \b2v_inst.state_17_LC_7_13_6 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \b2v_inst.state_17_LC_7_13_6  (
            .in0(N__15865),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15910),
            .lcout(\b2v_inst.stateZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22554),
            .ce(),
            .sr(N__22899));
    defparam \b2v_inst.state_9_LC_7_13_7 .C_ON=1'b0;
    defparam \b2v_inst.state_9_LC_7_13_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.state_9_LC_7_13_7 .LUT_INIT=16'b1010101010101000;
    LogicCell40 \b2v_inst.state_9_LC_7_13_7  (
            .in0(N__13893),
            .in1(N__16076),
            .in2(N__16229),
            .in3(N__16173),
            .lcout(\b2v_inst.stateZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22554),
            .ce(),
            .sr(N__22899));
    defparam \b2v_inst.dir_mem_1_RNI3UAQ_6_LC_7_14_0 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_1_RNI3UAQ_6_LC_7_14_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_1_RNI3UAQ_6_LC_7_14_0 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \b2v_inst.dir_mem_1_RNI3UAQ_6_LC_7_14_0  (
            .in0(N__16286),
            .in1(N__16465),
            .in2(N__14111),
            .in3(N__15369),
            .lcout(\b2v_inst.addr_ram_1_iv_i_1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNIMMMH_6_LC_7_14_1 .C_ON=1'b0;
    defparam \b2v_inst.state_RNIMMMH_6_LC_7_14_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNIMMMH_6_LC_7_14_1 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \b2v_inst.state_RNIMMMH_6_LC_7_14_1  (
            .in0(N__15184),
            .in1(N__15847),
            .in2(_gnd_net_),
            .in3(N__20631),
            .lcout(),
            .ltout(\b2v_inst.N_399_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_3_RNIIE1F1_6_LC_7_14_2 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_3_RNIIE1F1_6_LC_7_14_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_3_RNIIE1F1_6_LC_7_14_2 .LUT_INIT=16'b1111101111110011;
    LogicCell40 \b2v_inst.dir_mem_3_RNIIE1F1_6_LC_7_14_2  (
            .in0(N__14135),
            .in1(N__15139),
            .in2(N__13949),
            .in3(N__16936),
            .lcout(),
            .ltout(\b2v_inst.addr_ram_1_iv_i_2_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_RNIG3L83_6_LC_7_14_3 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_RNIG3L83_6_LC_7_14_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNIG3L83_6_LC_7_14_3 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \b2v_inst.dir_mem_RNIG3L83_6_LC_7_14_3  (
            .in0(N__16395),
            .in1(N__13946),
            .in2(N__13940),
            .in3(N__19127),
            .lcout(N_165),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_12_LC_7_14_4 .C_ON=1'b0;
    defparam \b2v_inst.state_12_LC_7_14_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.state_12_LC_7_14_4 .LUT_INIT=16'b1000100010001100;
    LogicCell40 \b2v_inst.state_12_LC_7_14_4  (
            .in0(N__15946),
            .in1(N__15370),
            .in2(N__16115),
            .in3(N__14820),
            .lcout(\b2v_inst.stateZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22589),
            .ce(),
            .sr(N__22904));
    defparam \b2v_inst.state_RNI3SA9_13_LC_7_14_5 .C_ON=1'b0;
    defparam \b2v_inst.state_RNI3SA9_13_LC_7_14_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNI3SA9_13_LC_7_14_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \b2v_inst.state_RNI3SA9_13_LC_7_14_5  (
            .in0(_gnd_net_),
            .in1(N__15945),
            .in2(_gnd_net_),
            .in3(N__13894),
            .lcout(\b2v_inst.N_235 ),
            .ltout(\b2v_inst.N_235_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_1_RNIKA1U_7_LC_7_14_6 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_1_RNIKA1U_7_LC_7_14_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_1_RNIKA1U_7_LC_7_14_6 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \b2v_inst.dir_mem_1_RNIKA1U_7_LC_7_14_6  (
            .in0(N__15287),
            .in1(N__18041),
            .in2(N__14099),
            .in3(N__16935),
            .lcout(\b2v_inst.addr_ram_1_0_iv_i_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_10_LC_7_15_0 .C_ON=1'b0;
    defparam \b2v_inst.state_10_LC_7_15_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.state_10_LC_7_15_0 .LUT_INIT=16'b1111000000010000;
    LogicCell40 \b2v_inst.state_10_LC_7_15_0  (
            .in0(N__14825),
            .in1(N__16111),
            .in2(N__16480),
            .in3(N__14096),
            .lcout(\b2v_inst.stateZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22352),
            .ce(),
            .sr(N__22909));
    defparam \b2v_inst.dir_mem_1_RNIPJAQ_1_LC_7_15_1 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_1_RNIPJAQ_1_LC_7_15_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_1_RNIPJAQ_1_LC_7_15_1 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \b2v_inst.dir_mem_1_RNIPJAQ_1_LC_7_15_1  (
            .in0(N__19949),
            .in1(N__16466),
            .in2(N__16526),
            .in3(N__15371),
            .lcout(\b2v_inst.addr_ram_1_0_iv_i_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNIVNA9_11_LC_7_15_2 .C_ON=1'b0;
    defparam \b2v_inst.state_RNIVNA9_11_LC_7_15_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNIVNA9_11_LC_7_15_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \b2v_inst.state_RNIVNA9_11_LC_7_15_2  (
            .in0(_gnd_net_),
            .in1(N__14095),
            .in2(_gnd_net_),
            .in3(N__15469),
            .lcout(\b2v_inst.N_237 ),
            .ltout(\b2v_inst.N_237_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_1_RNINHAQ_0_LC_7_15_3 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_1_RNINHAQ_0_LC_7_15_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_1_RNINHAQ_0_LC_7_15_3 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \b2v_inst.dir_mem_1_RNINHAQ_0_LC_7_15_3  (
            .in0(N__16493),
            .in1(N__20162),
            .in2(N__14072),
            .in3(N__15372),
            .lcout(),
            .ltout(\b2v_inst.addr_ram_1_iv_i_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_RNIG4063_0_LC_7_15_4 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_RNIG4063_0_LC_7_15_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNIG4063_0_LC_7_15_4 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \b2v_inst.dir_mem_RNIG4063_0_LC_7_15_4  (
            .in0(N__19895),
            .in1(N__14069),
            .in2(N__14063),
            .in3(N__16396),
            .lcout(N_167),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_RNIQQMS2_1_LC_7_15_5 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_RNIQQMS2_1_LC_7_15_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNIQQMS2_1_LC_7_15_5 .LUT_INIT=16'b1111111011101110;
    LogicCell40 \b2v_inst.dir_mem_RNIQQMS2_1_LC_7_15_5  (
            .in0(N__14162),
            .in1(N__14033),
            .in2(N__16405),
            .in3(N__19817),
            .lcout(N_60),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_1_RNIRLAQ_2_LC_7_15_6 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_1_RNIRLAQ_2_LC_7_15_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_1_RNIRLAQ_2_LC_7_15_6 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \b2v_inst.dir_mem_1_RNIRLAQ_2_LC_7_15_6  (
            .in0(N__15373),
            .in1(N__16508),
            .in2(N__16479),
            .in3(N__20000),
            .lcout(),
            .ltout(\b2v_inst.addr_ram_1_0_iv_i_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_RNIVVMS2_2_LC_7_15_7 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_RNIVVMS2_2_LC_7_15_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNIVVMS2_2_LC_7_15_7 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \b2v_inst.dir_mem_RNIVVMS2_2_LC_7_15_7  (
            .in0(N__16400),
            .in1(N__16880),
            .in2(N__14003),
            .in3(N__19217),
            .lcout(N_56),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_RNI88AO1_7_LC_7_16_0 .C_ON=1'b0;
    defparam \b2v_inst.indice_RNI88AO1_7_LC_7_16_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_RNI88AO1_7_LC_7_16_0 .LUT_INIT=16'b1111000111110101;
    LogicCell40 \b2v_inst.indice_RNI88AO1_7_LC_7_16_0  (
            .in0(N__20936),
            .in1(N__20632),
            .in2(N__17900),
            .in3(N__20503),
            .lcout(\b2v_inst.dir_mem_315_0 ),
            .ltout(\b2v_inst.dir_mem_315_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_3_1_LC_7_16_1 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_3_1_LC_7_16_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.dir_mem_3_1_LC_7_16_1 .LUT_INIT=16'b0101010110100101;
    LogicCell40 \b2v_inst.dir_mem_3_1_LC_7_16_1  (
            .in0(N__23027),
            .in1(_gnd_net_),
            .in2(N__14171),
            .in3(N__23211),
            .lcout(\b2v_inst.dir_mem_3Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22595),
            .ce(N__15274),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_3_2_LC_7_16_2 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_3_2_LC_7_16_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.dir_mem_3_2_LC_7_16_2 .LUT_INIT=16'b0110101010011001;
    LogicCell40 \b2v_inst.dir_mem_3_2_LC_7_16_2  (
            .in0(N__20147),
            .in1(N__23028),
            .in2(N__23219),
            .in3(N__15316),
            .lcout(\b2v_inst.dir_mem_3Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22595),
            .ce(N__15274),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_3_RNIBL331_1_LC_7_16_3 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_3_RNIBL331_1_LC_7_16_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_3_RNIBL331_1_LC_7_16_3 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \b2v_inst.dir_mem_3_RNIBL331_1_LC_7_16_3  (
            .in0(N__16952),
            .in1(N__14168),
            .in2(N__23054),
            .in3(N__17000),
            .lcout(\b2v_inst.addr_ram_1_0_iv_i_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_3_0_LC_7_16_4 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_3_0_LC_7_16_4 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.dir_mem_3_0_LC_7_16_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \b2v_inst.dir_mem_3_0_LC_7_16_4  (
            .in0(N__23210),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15315),
            .lcout(\b2v_inst.dir_mem_3Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22595),
            .ce(N__15274),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_3_5_LC_7_16_5 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_3_5_LC_7_16_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.dir_mem_3_5_LC_7_16_5 .LUT_INIT=16'b1001010110101001;
    LogicCell40 \b2v_inst.dir_mem_3_5_LC_7_16_5  (
            .in0(N__20504),
            .in1(N__16247),
            .in2(N__15325),
            .in3(N__18027),
            .lcout(\b2v_inst.dir_mem_3Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22595),
            .ce(N__15274),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_3_4_LC_7_16_6 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_3_4_LC_7_16_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.dir_mem_3_4_LC_7_16_6 .LUT_INIT=16'b0110011001011010;
    LogicCell40 \b2v_inst.dir_mem_3_4_LC_7_16_6  (
            .in0(N__18026),
            .in1(N__20825),
            .in2(N__15980),
            .in3(N__15317),
            .lcout(\b2v_inst.dir_mem_3Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22595),
            .ce(N__15274),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_3_6_LC_7_16_7 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_3_6_LC_7_16_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.dir_mem_3_6_LC_7_16_7 .LUT_INIT=16'b0101011010100110;
    LogicCell40 \b2v_inst.dir_mem_3_6_LC_7_16_7  (
            .in0(N__20633),
            .in1(N__16274),
            .in2(N__15326),
            .in3(N__16553),
            .lcout(\b2v_inst.dir_mem_3Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22595),
            .ce(N__15274),
            .sr(_gnd_net_));
    defparam \b2v_inst.data_a_escribir_RNID9JL_7_LC_7_17_0 .C_ON=1'b0;
    defparam \b2v_inst.data_a_escribir_RNID9JL_7_LC_7_17_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.data_a_escribir_RNID9JL_7_LC_7_17_0 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \b2v_inst.data_a_escribir_RNID9JL_7_LC_7_17_0  (
            .in0(N__17679),
            .in1(N__14371),
            .in2(_gnd_net_),
            .in3(N__17017),
            .lcout(N_205_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_2_6_LC_7_17_1 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_2_6_LC_7_17_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.dir_mem_2_6_LC_7_17_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \b2v_inst.dir_mem_2_6_LC_7_17_1  (
            .in0(N__20354),
            .in1(N__16732),
            .in2(_gnd_net_),
            .in3(N__15731),
            .lcout(\b2v_inst.dir_mem_2Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22354),
            .ce(N__16682),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_RX_Byte_RNO_0_3_LC_7_17_6 .C_ON=1'b0;
    defparam \b2v_inst1.r_RX_Byte_RNO_0_3_LC_7_17_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_RX_Byte_RNO_0_3_LC_7_17_6 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \b2v_inst1.r_RX_Byte_RNO_0_3_LC_7_17_6  (
            .in0(N__18163),
            .in1(N__18251),
            .in2(_gnd_net_),
            .in3(N__18123),
            .lcout(\b2v_inst1.r_RX_Bytece_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_RX_Byte_RNO_0_4_LC_7_17_7 .C_ON=1'b0;
    defparam \b2v_inst1.r_RX_Byte_RNO_0_4_LC_7_17_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_RX_Byte_RNO_0_4_LC_7_17_7 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \b2v_inst1.r_RX_Byte_RNO_0_4_LC_7_17_7  (
            .in0(N__18124),
            .in1(_gnd_net_),
            .in2(N__18259),
            .in3(N__18164),
            .lcout(\b2v_inst1.r_RX_Bytece_0_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst3.data_to_send_esr_3_LC_7_18_3 .C_ON=1'b0;
    defparam \b2v_inst3.data_to_send_esr_3_LC_7_18_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst3.data_to_send_esr_3_LC_7_18_3 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \b2v_inst3.data_to_send_esr_3_LC_7_18_3  (
            .in0(N__14413),
            .in1(N__14545),
            .in2(N__14498),
            .in3(N__14346),
            .lcout(\b2v_inst3.data_to_sendZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22242),
            .ce(N__14254),
            .sr(N__22915));
    defparam \b2v_inst3.data_to_send_esr_4_LC_7_18_4 .C_ON=1'b0;
    defparam \b2v_inst3.data_to_send_esr_4_LC_7_18_4 .SEQ_MODE=4'b1000;
    defparam \b2v_inst3.data_to_send_esr_4_LC_7_18_4 .LUT_INIT=16'b1010000011100100;
    LogicCell40 \b2v_inst3.data_to_send_esr_4_LC_7_18_4  (
            .in0(N__14344),
            .in1(N__14516),
            .in2(N__14465),
            .in3(N__14414),
            .lcout(\b2v_inst3.data_to_sendZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22242),
            .ce(N__14254),
            .sr(N__22915));
    defparam \b2v_inst3.data_to_send_esr_5_LC_7_18_5 .C_ON=1'b0;
    defparam \b2v_inst3.data_to_send_esr_5_LC_7_18_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst3.data_to_send_esr_5_LC_7_18_5 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \b2v_inst3.data_to_send_esr_5_LC_7_18_5  (
            .in0(N__14415),
            .in1(N__14485),
            .in2(N__14429),
            .in3(N__14347),
            .lcout(\b2v_inst3.data_to_sendZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22242),
            .ce(N__14254),
            .sr(N__22915));
    defparam \b2v_inst3.data_to_send_esr_6_LC_7_18_6 .C_ON=1'b0;
    defparam \b2v_inst3.data_to_send_esr_6_LC_7_18_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst3.data_to_send_esr_6_LC_7_18_6 .LUT_INIT=16'b1010000011100100;
    LogicCell40 \b2v_inst3.data_to_send_esr_6_LC_7_18_6  (
            .in0(N__14345),
            .in1(N__14455),
            .in2(N__14270),
            .in3(N__14416),
            .lcout(\b2v_inst3.data_to_sendZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22242),
            .ce(N__14254),
            .sr(N__22915));
    defparam \b2v_inst3.data_to_send_esr_7_LC_7_18_7 .C_ON=1'b0;
    defparam \b2v_inst3.data_to_send_esr_7_LC_7_18_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst3.data_to_send_esr_7_LC_7_18_7 .LUT_INIT=16'b1100110001010000;
    LogicCell40 \b2v_inst3.data_to_send_esr_7_LC_7_18_7  (
            .in0(N__14417),
            .in1(N__14269),
            .in2(N__14375),
            .in3(N__14348),
            .lcout(\b2v_inst3.data_to_sendZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22242),
            .ce(N__14254),
            .sr(N__22915));
    defparam \b2v_inst.reg_anterior_6_LC_7_19_0 .C_ON=1'b0;
    defparam \b2v_inst.reg_anterior_6_LC_7_19_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_anterior_6_LC_7_19_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \b2v_inst.reg_anterior_6_LC_7_19_0  (
            .in0(N__15535),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14242),
            .lcout(\b2v_inst.reg_anteriorZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22243),
            .ce(N__15235),
            .sr(N__22919));
    defparam \b2v_inst.reg_anterior_5_LC_7_19_1 .C_ON=1'b0;
    defparam \b2v_inst.reg_anterior_5_LC_7_19_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.reg_anterior_5_LC_7_19_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \b2v_inst.reg_anterior_5_LC_7_19_1  (
            .in0(_gnd_net_),
            .in1(N__15534),
            .in2(_gnd_net_),
            .in3(N__14705),
            .lcout(\b2v_inst.reg_anteriorZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22243),
            .ce(N__15235),
            .sr(N__22919));
    defparam \b2v_inst.cuenta_RNI5B3A_6_LC_8_11_0 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_RNI5B3A_6_LC_8_11_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.cuenta_RNI5B3A_6_LC_8_11_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst.cuenta_RNI5B3A_6_LC_8_11_0  (
            .in0(_gnd_net_),
            .in1(N__14952),
            .in2(_gnd_net_),
            .in3(N__15053),
            .lcout(),
            .ltout(\b2v_inst.un4_cuenta_ac0_11_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.cuenta_RNI4SC81_7_LC_8_11_1 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_RNI4SC81_7_LC_8_11_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.cuenta_RNI4SC81_7_LC_8_11_1 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \b2v_inst.cuenta_RNI4SC81_7_LC_8_11_1  (
            .in0(N__14985),
            .in1(N__14924),
            .in2(N__14624),
            .in3(N__15022),
            .lcout(\b2v_inst.cuenta_RNI4SC81Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.cuenta_RNIK17D1_4_LC_8_11_2 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_RNIK17D1_4_LC_8_11_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.cuenta_RNIK17D1_4_LC_8_11_2 .LUT_INIT=16'b1111111101100110;
    LogicCell40 \b2v_inst.cuenta_RNIK17D1_4_LC_8_11_2  (
            .in0(N__15026),
            .in1(N__14984),
            .in2(_gnd_net_),
            .in3(N__14621),
            .lcout(\b2v_inst.cuenta_5_i_o2_0_0_1 ),
            .ltout(\b2v_inst.cuenta_5_i_o2_0_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.cuenta_RNIO2VO3_4_LC_8_11_3 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_RNIO2VO3_4_LC_8_11_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.cuenta_RNIO2VO3_4_LC_8_11_3 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \b2v_inst.cuenta_RNIO2VO3_4_LC_8_11_3  (
            .in0(_gnd_net_),
            .in1(N__16202),
            .in2(N__14612),
            .in3(N__16150),
            .lcout(\b2v_inst.cuenta_RNIO2VO3Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.cuenta_RNI05B31_6_LC_8_11_4 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_RNI05B31_6_LC_8_11_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.cuenta_RNI05B31_6_LC_8_11_4 .LUT_INIT=16'b0111111011101110;
    LogicCell40 \b2v_inst.cuenta_RNI05B31_6_LC_8_11_4  (
            .in0(N__14957),
            .in1(N__15054),
            .in2(N__15029),
            .in3(N__14986),
            .lcout(\b2v_inst.state_ns_a2_0_o2_1_0_2 ),
            .ltout(\b2v_inst.state_ns_a2_0_o2_1_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_17_rep1_RNICDK34_LC_8_11_5 .C_ON=1'b0;
    defparam \b2v_inst.state_17_rep1_RNICDK34_LC_8_11_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_17_rep1_RNICDK34_LC_8_11_5 .LUT_INIT=16'b0101010101010100;
    LogicCell40 \b2v_inst.state_17_rep1_RNICDK34_LC_8_11_5  (
            .in0(N__19080),
            .in1(N__16151),
            .in2(N__14609),
            .in3(N__14605),
            .lcout(),
            .ltout(\b2v_inst.state_17_rep1_RNICDKZ0Z34_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_17_rep1_RNIOVB69_LC_8_11_6 .C_ON=1'b0;
    defparam \b2v_inst.state_17_rep1_RNIOVB69_LC_8_11_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_17_rep1_RNIOVB69_LC_8_11_6 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \b2v_inst.state_17_rep1_RNIOVB69_LC_8_11_6  (
            .in0(_gnd_net_),
            .in1(N__18749),
            .in2(N__14594),
            .in3(N__14591),
            .lcout(\b2v_inst.N_374 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.cuenta_5_LC_8_11_7 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_5_LC_8_11_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.cuenta_5_LC_8_11_7 .LUT_INIT=16'b0000000001111000;
    LogicCell40 \b2v_inst.cuenta_5_LC_8_11_7  (
            .in0(N__14987),
            .in1(N__15027),
            .in2(N__15062),
            .in3(N__14858),
            .lcout(\b2v_inst.cuentaZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21971),
            .ce(N__14906),
            .sr(N__22896));
    defparam \b2v_inst.dir_mem_RNO_3_0_LC_8_12_0 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_RNO_3_0_LC_8_12_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNO_3_0_LC_8_12_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst.dir_mem_RNO_3_0_LC_8_12_0  (
            .in0(N__14927),
            .in1(N__14955),
            .in2(N__17572),
            .in3(N__15060),
            .lcout(\b2v_inst.un2_indice_3_0_iv_0_a2_5_sx_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.cuenta_RNI925F_7_LC_8_12_2 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_RNI925F_7_LC_8_12_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.cuenta_RNI925F_7_LC_8_12_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \b2v_inst.cuenta_RNI925F_7_LC_8_12_2  (
            .in0(N__14926),
            .in1(N__14954),
            .in2(_gnd_net_),
            .in3(N__15059),
            .lcout(\b2v_inst.cuenta_RNI925FZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.cuenta_RNO_0_6_LC_8_12_3 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_RNO_0_6_LC_8_12_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.cuenta_RNO_0_6_LC_8_12_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \b2v_inst.cuenta_RNO_0_6_LC_8_12_3  (
            .in0(N__15061),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15028),
            .lcout(),
            .ltout(\b2v_inst.un4_cuenta_ac0_9_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.cuenta_6_LC_8_12_4 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_6_LC_8_12_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.cuenta_6_LC_8_12_4 .LUT_INIT=16'b0001010001000100;
    LogicCell40 \b2v_inst.cuenta_6_LC_8_12_4  (
            .in0(N__14856),
            .in1(N__14956),
            .in2(N__14993),
            .in3(N__14990),
            .lcout(\b2v_inst.cuentaZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22187),
            .ce(N__14897),
            .sr(N__22900));
    defparam \b2v_inst.cuenta_7_LC_8_12_5 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_7_LC_8_12_5 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.cuenta_7_LC_8_12_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \b2v_inst.cuenta_7_LC_8_12_5  (
            .in0(_gnd_net_),
            .in1(N__14857),
            .in2(_gnd_net_),
            .in3(N__16169),
            .lcout(\b2v_inst.cuentaZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22187),
            .ce(N__14897),
            .sr(N__22900));
    defparam \b2v_inst.state_17_rep1_RNI8QDK1_LC_8_12_6 .C_ON=1'b0;
    defparam \b2v_inst.state_17_rep1_RNI8QDK1_LC_8_12_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_17_rep1_RNI8QDK1_LC_8_12_6 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \b2v_inst.state_17_rep1_RNI8QDK1_LC_8_12_6  (
            .in0(_gnd_net_),
            .in1(N__19052),
            .in2(_gnd_net_),
            .in3(N__18699),
            .lcout(\b2v_inst.N_227 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.cuenta_RNI41OB2_6_LC_8_13_0 .C_ON=1'b0;
    defparam \b2v_inst.cuenta_RNI41OB2_6_LC_8_13_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.cuenta_RNI41OB2_6_LC_8_13_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \b2v_inst.cuenta_RNI41OB2_6_LC_8_13_0  (
            .in0(_gnd_net_),
            .in1(N__16221),
            .in2(_gnd_net_),
            .in3(N__16170),
            .lcout(\b2v_inst.N_232 ),
            .ltout(\b2v_inst.N_232_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_14_LC_8_13_1 .C_ON=1'b0;
    defparam \b2v_inst.state_14_LC_8_13_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.state_14_LC_8_13_1 .LUT_INIT=16'b1111111100000010;
    LogicCell40 \b2v_inst.state_14_LC_8_13_1  (
            .in0(N__15214),
            .in1(N__16101),
            .in2(N__14801),
            .in3(N__18985),
            .lcout(\b2v_inst.stateZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22468),
            .ce(),
            .sr(N__22905));
    defparam \b2v_inst.state_7_LC_8_13_2 .C_ON=1'b0;
    defparam \b2v_inst.state_7_LC_8_13_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.state_7_LC_8_13_2 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \b2v_inst.state_7_LC_8_13_2  (
            .in0(N__16222),
            .in1(N__15215),
            .in2(N__16112),
            .in3(N__16171),
            .lcout(\b2v_inst.stateZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22468),
            .ce(),
            .sr(N__22905));
    defparam \b2v_inst.state_fast_15_LC_8_13_3 .C_ON=1'b0;
    defparam \b2v_inst.state_fast_15_LC_8_13_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.state_fast_15_LC_8_13_3 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \b2v_inst.state_fast_15_LC_8_13_3  (
            .in0(N__16172),
            .in1(N__16223),
            .in2(N__16044),
            .in3(N__16100),
            .lcout(\b2v_inst.state_fastZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22468),
            .ce(),
            .sr(N__22905));
    defparam \b2v_inst.state_RNIRA0K_15_LC_8_13_4 .C_ON=1'b0;
    defparam \b2v_inst.state_RNIRA0K_15_LC_8_13_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNIRA0K_15_LC_8_13_4 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \b2v_inst.state_RNIRA0K_15_LC_8_13_4  (
            .in0(N__18984),
            .in1(N__19062),
            .in2(_gnd_net_),
            .in3(N__15213),
            .lcout(\b2v_inst.N_239 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_RNO_2_6_LC_8_13_5 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_RNO_2_6_LC_8_13_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNO_2_6_LC_8_13_5 .LUT_INIT=16'b1101110111111111;
    LogicCell40 \b2v_inst.dir_mem_RNO_2_6_LC_8_13_5  (
            .in0(N__18918),
            .in1(N__19076),
            .in2(_gnd_net_),
            .in3(N__18983),
            .lcout(\b2v_inst.N_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNITETB_0_LC_8_14_0 .C_ON=1'b0;
    defparam \b2v_inst.state_RNITETB_0_LC_8_14_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNITETB_0_LC_8_14_0 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \b2v_inst.state_RNITETB_0_LC_8_14_0  (
            .in0(N__15073),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15439),
            .lcout(\b2v_inst.state_RNITETBZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_1_RNITNAQ_3_LC_8_14_1 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_1_RNITNAQ_3_LC_8_14_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_1_RNITNAQ_3_LC_8_14_1 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \b2v_inst.dir_mem_1_RNITNAQ_3_LC_8_14_1  (
            .in0(N__15374),
            .in1(N__15989),
            .in2(N__20210),
            .in3(N__16458),
            .lcout(\b2v_inst.addr_ram_1_iv_i_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNIHV0E_6_LC_8_14_2 .C_ON=1'b0;
    defparam \b2v_inst.state_RNIHV0E_6_LC_8_14_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNIHV0E_6_LC_8_14_2 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \b2v_inst.state_RNIHV0E_6_LC_8_14_2  (
            .in0(N__15185),
            .in1(N__15871),
            .in2(_gnd_net_),
            .in3(N__17115),
            .lcout(),
            .ltout(\b2v_inst.N_351_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_3_RNIAKBB1_3_LC_8_14_3 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_3_RNIAKBB1_3_LC_8_14_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_3_RNIAKBB1_3_LC_8_14_3 .LUT_INIT=16'b1111101111110011;
    LogicCell40 \b2v_inst.dir_mem_3_RNIAKBB1_3_LC_8_14_3  (
            .in0(N__15296),
            .in1(N__15138),
            .in2(N__15119),
            .in3(N__16946),
            .lcout(),
            .ltout(\b2v_inst.addr_ram_1_iv_i_2_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_RNIVVU43_3_LC_8_14_4 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_RNIVVU43_3_LC_8_14_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNIVVU43_3_LC_8_14_4 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \b2v_inst.dir_mem_RNIVVU43_3_LC_8_14_4  (
            .in0(N__16374),
            .in1(N__15116),
            .in2(N__15110),
            .in3(N__19322),
            .lcout(N_58),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_0_LC_8_14_5 .C_ON=1'b0;
    defparam \b2v_inst.state_0_LC_8_14_5 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.state_0_LC_8_14_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst.state_0_LC_8_14_5  (
            .in0(N__15440),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22355),
            .ce(),
            .sr(N__22910));
    defparam \b2v_inst.state_1_LC_8_14_6 .C_ON=1'b0;
    defparam \b2v_inst.state_1_LC_8_14_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.state_1_LC_8_14_6 .LUT_INIT=16'b1111111000000000;
    LogicCell40 \b2v_inst.state_1_LC_8_14_6  (
            .in0(N__16224),
            .in1(N__16174),
            .in2(N__16114),
            .in3(N__15470),
            .lcout(\b2v_inst.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22355),
            .ce(),
            .sr(N__22910));
    defparam \b2v_inst.dir_mem_3_RNIHR331_4_LC_8_15_0 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_3_RNIHR331_4_LC_8_15_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_3_RNIHR331_4_LC_8_15_0 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \b2v_inst.dir_mem_3_RNIHR331_4_LC_8_15_0  (
            .in0(N__17012),
            .in1(N__16953),
            .in2(N__15431),
            .in3(N__18005),
            .lcout(),
            .ltout(\b2v_inst.addr_ram_1_0_iv_i_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_RNI9ANS2_4_LC_8_15_1 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_RNI9ANS2_4_LC_8_15_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNI9ANS2_4_LC_8_15_1 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \b2v_inst.dir_mem_RNI9ANS2_4_LC_8_15_1  (
            .in0(N__16394),
            .in1(N__15332),
            .in2(N__15419),
            .in3(N__19373),
            .lcout(N_163),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_1_RNO_1_4_LC_8_15_2 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_1_RNO_1_4_LC_8_15_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_1_RNO_1_4_LC_8_15_2 .LUT_INIT=16'b0111011100010001;
    LogicCell40 \b2v_inst.dir_mem_1_RNO_1_4_LC_8_15_2  (
            .in0(N__20492),
            .in1(N__20687),
            .in2(_gnd_net_),
            .in3(N__18006),
            .lcout(),
            .ltout(\b2v_inst.g0_11_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_1_4_LC_8_15_3 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_1_4_LC_8_15_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.dir_mem_1_4_LC_8_15_3 .LUT_INIT=16'b1001101010011001;
    LogicCell40 \b2v_inst.dir_mem_1_4_LC_8_15_3  (
            .in0(N__18007),
            .in1(N__17912),
            .in2(N__15389),
            .in3(N__20610),
            .lcout(\b2v_inst.dir_mem_1Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22351),
            .ce(N__19920),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_1_RNIVPAQ_4_LC_8_15_4 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_1_RNIVPAQ_4_LC_8_15_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_1_RNIVPAQ_4_LC_8_15_4 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \b2v_inst.dir_mem_1_RNIVPAQ_4_LC_8_15_4  (
            .in0(N__16474),
            .in1(N__15386),
            .in2(N__16541),
            .in3(N__15376),
            .lcout(\b2v_inst.addr_ram_1_0_iv_i_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_3_3_LC_8_16_0 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_3_3_LC_8_16_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.dir_mem_3_3_LC_8_16_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst.dir_mem_3_3_LC_8_16_0  (
            .in0(N__15761),
            .in1(N__17045),
            .in2(_gnd_net_),
            .in3(N__15324),
            .lcout(\b2v_inst.dir_mem_3Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22594),
            .ce(N__15275),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_3_7_LC_8_16_1 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_3_7_LC_8_16_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.dir_mem_3_7_LC_8_16_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \b2v_inst.dir_mem_3_7_LC_8_16_1  (
            .in0(N__20639),
            .in1(N__16270),
            .in2(_gnd_net_),
            .in3(N__20934),
            .lcout(\b2v_inst.dir_mem_3Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22594),
            .ce(N__15275),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_RX_Byte_RNO_0_5_LC_8_16_2 .C_ON=1'b0;
    defparam \b2v_inst1.r_RX_Byte_RNO_0_5_LC_8_16_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_RX_Byte_RNO_0_5_LC_8_16_2 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \b2v_inst1.r_RX_Byte_RNO_0_5_LC_8_16_2  (
            .in0(N__18191),
            .in1(N__18104),
            .in2(_gnd_net_),
            .in3(N__18239),
            .lcout(\b2v_inst1.r_RX_Bytece_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_SM_Main_RNIC98H_2_LC_8_16_4 .C_ON=1'b0;
    defparam \b2v_inst1.r_SM_Main_RNIC98H_2_LC_8_16_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_SM_Main_RNIC98H_2_LC_8_16_4 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \b2v_inst1.r_SM_Main_RNIC98H_2_LC_8_16_4  (
            .in0(N__23483),
            .in1(N__23753),
            .in2(_gnd_net_),
            .in3(N__23629),
            .lcout(\b2v_inst1.r_SM_Main_d_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_3_RNO_0_3_LC_8_17_0 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_3_RNO_0_3_LC_8_17_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_3_RNO_0_3_LC_8_17_0 .LUT_INIT=16'b1100110010011001;
    LogicCell40 \b2v_inst.dir_mem_3_RNO_0_3_LC_8_17_0  (
            .in0(N__23081),
            .in1(N__20332),
            .in2(_gnd_net_),
            .in3(N__20140),
            .lcout(\b2v_inst.dir_mem_3_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_RX_Byte_RNO_0_1_LC_8_17_3 .C_ON=1'b0;
    defparam \b2v_inst1.r_RX_Byte_RNO_0_1_LC_8_17_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_RX_Byte_RNO_0_1_LC_8_17_3 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \b2v_inst1.r_RX_Byte_RNO_0_1_LC_8_17_3  (
            .in0(N__18119),
            .in1(N__18165),
            .in2(_gnd_net_),
            .in3(N__18255),
            .lcout(),
            .ltout(\b2v_inst1.r_RX_Bytece_0_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_RX_Byte_1_LC_8_17_4 .C_ON=1'b0;
    defparam \b2v_inst1.r_RX_Byte_1_LC_8_17_4 .SEQ_MODE=4'b1000;
    defparam \b2v_inst1.r_RX_Byte_1_LC_8_17_4 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \b2v_inst1.r_RX_Byte_1_LC_8_17_4  (
            .in0(N__15742),
            .in1(N__22708),
            .in2(N__15752),
            .in3(N__17170),
            .lcout(SYNTHESIZED_WIRE_10_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22353),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_2_RNO_0_6_LC_8_17_7 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_2_RNO_0_6_LC_8_17_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_2_RNO_0_6_LC_8_17_7 .LUT_INIT=16'b0011011011001100;
    LogicCell40 \b2v_inst.dir_mem_2_RNO_0_6_LC_8_17_7  (
            .in0(N__18028),
            .in1(N__20636),
            .in2(N__17060),
            .in3(N__20501),
            .lcout(\b2v_inst.dir_mem_2_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_Bit_Index_0_LC_8_18_0 .C_ON=1'b0;
    defparam \b2v_inst1.r_Bit_Index_0_LC_8_18_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst1.r_Bit_Index_0_LC_8_18_0 .LUT_INIT=16'b1111000011010010;
    LogicCell40 \b2v_inst1.r_Bit_Index_0_LC_8_18_0  (
            .in0(N__16633),
            .in1(N__23494),
            .in2(N__18185),
            .in3(N__23754),
            .lcout(\b2v_inst1.r_Bit_IndexZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22593),
            .ce(),
            .sr(N__24063));
    defparam \b2v_inst1.r_RX_DV_LC_8_18_1 .C_ON=1'b0;
    defparam \b2v_inst1.r_RX_DV_LC_8_18_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst1.r_RX_DV_LC_8_18_1 .LUT_INIT=16'b1110100011100000;
    LogicCell40 \b2v_inst1.r_RX_DV_LC_8_18_1  (
            .in0(N__23755),
            .in1(N__23630),
            .in2(N__15719),
            .in3(N__16634),
            .lcout(SYNTHESIZED_WIRE_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22593),
            .ce(),
            .sr(N__24063));
    defparam \b2v_inst.ignorar_anterior_LC_8_20_0 .C_ON=1'b0;
    defparam \b2v_inst.ignorar_anterior_LC_8_20_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.ignorar_anterior_LC_8_20_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst.ignorar_anterior_LC_8_20_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15684),
            .lcout(\b2v_inst.ignorar_anteriorZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22480),
            .ce(N__15521),
            .sr(N__22921));
    defparam \b2v_inst.dir_mem_RNO_0_6_LC_9_10_0 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_RNO_0_6_LC_9_10_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNO_0_6_LC_9_10_0 .LUT_INIT=16'b0000000011001010;
    LogicCell40 \b2v_inst.dir_mem_RNO_0_6_LC_9_10_0  (
            .in0(N__15797),
            .in1(N__15803),
            .in2(N__15506),
            .in3(N__18775),
            .lcout(),
            .ltout(\b2v_inst.N_7_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_6_LC_9_10_1 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_6_LC_9_10_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.dir_mem_6_LC_9_10_1 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \b2v_inst.dir_mem_6_LC_9_10_1  (
            .in0(N__17828),
            .in1(N__16808),
            .in2(N__15809),
            .in3(N__16574),
            .lcout(\b2v_inst.dir_memZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22392),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_RNO_5_6_LC_9_10_2 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_RNO_5_6_LC_9_10_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNO_5_6_LC_9_10_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst.dir_mem_RNO_5_6_LC_9_10_2  (
            .in0(_gnd_net_),
            .in1(N__19320),
            .in2(_gnd_net_),
            .in3(N__19213),
            .lcout(),
            .ltout(\b2v_inst.g2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_RNO_3_6_LC_9_10_3 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_RNO_3_6_LC_9_10_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNO_3_6_LC_9_10_3 .LUT_INIT=16'b1010101001101010;
    LogicCell40 \b2v_inst.dir_mem_RNO_3_6_LC_9_10_3  (
            .in0(N__19112),
            .in1(N__15926),
            .in2(N__15806),
            .in3(N__19727),
            .lcout(\b2v_inst.g1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_RNO_4_6_LC_9_10_4 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_RNO_4_6_LC_9_10_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNO_4_6_LC_9_10_4 .LUT_INIT=16'b1010101010011010;
    LogicCell40 \b2v_inst.dir_mem_RNO_4_6_LC_9_10_4  (
            .in0(N__20635),
            .in1(N__21145),
            .in2(N__16829),
            .in3(N__21059),
            .lcout(\b2v_inst.un2_indice_21_s0_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_RNITB3H1_6_LC_9_10_5 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_RNITB3H1_6_LC_9_10_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNITB3H1_6_LC_9_10_5 .LUT_INIT=16'b0011110010011001;
    LogicCell40 \b2v_inst.dir_mem_RNITB3H1_6_LC_9_10_5  (
            .in0(N__20634),
            .in1(N__17782),
            .in2(N__19119),
            .in3(N__19726),
            .lcout(\b2v_inst.dir_mem_RNITB3H1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_3_LC_9_11_1 .C_ON=1'b0;
    defparam \b2v_inst.indice_3_LC_9_11_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.indice_3_LC_9_11_1 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \b2v_inst.indice_3_LC_9_11_1  (
            .in0(N__20139),
            .in1(N__23134),
            .in2(N__20276),
            .in3(N__23084),
            .lcout(\b2v_inst.indiceZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22114),
            .ce(N__22952),
            .sr(N__22901));
    defparam \b2v_inst.state_fast_RNI711G_0_15_LC_9_11_2 .C_ON=1'b0;
    defparam \b2v_inst.state_fast_RNI711G_0_15_LC_9_11_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_fast_RNI711G_0_15_LC_9_11_2 .LUT_INIT=16'b0101010101110111;
    LogicCell40 \b2v_inst.state_fast_RNI711G_0_15_LC_9_11_2  (
            .in0(N__18916),
            .in1(N__15776),
            .in2(_gnd_net_),
            .in3(N__15787),
            .lcout(\b2v_inst.N_253 ),
            .ltout(\b2v_inst.N_253_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_RNIGVEE1_0_LC_9_11_3 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_RNIGVEE1_0_LC_9_11_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNIGVEE1_0_LC_9_11_3 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \b2v_inst.dir_mem_RNIGVEE1_0_LC_9_11_3  (
            .in0(N__19862),
            .in1(N__21038),
            .in2(N__15791),
            .in3(N__17768),
            .lcout(\b2v_inst.dir_mem_RNIGVEE1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_fast_RNI711G_15_LC_9_11_4 .C_ON=1'b0;
    defparam \b2v_inst.state_fast_RNI711G_15_LC_9_11_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_fast_RNI711G_15_LC_9_11_4 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \b2v_inst.state_fast_RNI711G_15_LC_9_11_4  (
            .in0(N__18917),
            .in1(N__15788),
            .in2(_gnd_net_),
            .in3(N__15775),
            .lcout(\b2v_inst.N_253_i ),
            .ltout(\b2v_inst.N_253_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_RNII5PO1_1_LC_9_11_5 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_RNII5PO1_1_LC_9_11_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNII5PO1_1_LC_9_11_5 .LUT_INIT=16'b0011110010100101;
    LogicCell40 \b2v_inst.dir_mem_RNII5PO1_1_LC_9_11_5  (
            .in0(N__21146),
            .in1(N__19816),
            .in2(N__15764),
            .in3(N__19721),
            .lcout(\b2v_inst.dir_mem_RNII5PO1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_RNIN53H1_3_LC_9_11_6 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_RNIN53H1_3_LC_9_11_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNIN53H1_3_LC_9_11_6 .LUT_INIT=16'b0100101111100001;
    LogicCell40 \b2v_inst.dir_mem_RNIN53H1_3_LC_9_11_6  (
            .in0(N__19723),
            .in1(N__20242),
            .in2(N__17790),
            .in3(N__19319),
            .lcout(\b2v_inst.dir_mem_RNIN53H1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_RNIL33H1_2_LC_9_11_7 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_RNIL33H1_2_LC_9_11_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNIL33H1_2_LC_9_11_7 .LUT_INIT=16'b0110011011000011;
    LogicCell40 \b2v_inst.dir_mem_RNIL33H1_2_LC_9_11_7  (
            .in0(N__19205),
            .in1(N__17764),
            .in2(N__20146),
            .in3(N__19722),
            .lcout(\b2v_inst.dir_mem_RNIL33H1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_17_rep1_RNIBDUK1_LC_9_12_0 .C_ON=1'b0;
    defparam \b2v_inst.state_17_rep1_RNIBDUK1_LC_9_12_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_17_rep1_RNIBDUK1_LC_9_12_0 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \b2v_inst.state_17_rep1_RNIBDUK1_LC_9_12_0  (
            .in0(N__18922),
            .in1(N__19066),
            .in2(_gnd_net_),
            .in3(N__18745),
            .lcout(\b2v_inst.N_467 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_RNO_0_0_LC_9_12_1 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_RNO_0_0_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNO_0_0_LC_9_12_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \b2v_inst.dir_mem_RNO_0_0_LC_9_12_1  (
            .in0(_gnd_net_),
            .in1(N__15959),
            .in2(_gnd_net_),
            .in3(N__17391),
            .lcout(),
            .ltout(\b2v_inst.N_452_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_0_LC_9_12_2 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_0_LC_9_12_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.dir_mem_0_LC_9_12_2 .LUT_INIT=16'b0000000001001100;
    LogicCell40 \b2v_inst.dir_mem_0_LC_9_12_2  (
            .in0(N__23152),
            .in1(N__16235),
            .in2(N__15953),
            .in3(N__17585),
            .lcout(\b2v_inst.dir_memZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22501),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNIL165_13_LC_9_12_3 .C_ON=1'b0;
    defparam \b2v_inst.state_RNIL165_13_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNIL165_13_LC_9_12_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst.state_RNIL165_13_LC_9_12_3  (
            .in0(_gnd_net_),
            .in1(N__18923),
            .in2(_gnd_net_),
            .in3(N__15950),
            .lcout(\b2v_inst.N_134_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_RNO_6_6_LC_9_12_5 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_RNO_6_6_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNO_6_6_LC_9_12_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst.dir_mem_RNO_6_6_LC_9_12_5  (
            .in0(N__19372),
            .in1(N__19815),
            .in2(N__19260),
            .in3(N__19869),
            .lcout(\b2v_inst.g2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_17_rep1_LC_9_13_0 .C_ON=1'b0;
    defparam \b2v_inst.state_17_rep1_LC_9_13_0 .SEQ_MODE=4'b1011;
    defparam \b2v_inst.state_17_rep1_LC_9_13_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \b2v_inst.state_17_rep1_LC_9_13_0  (
            .in0(_gnd_net_),
            .in1(N__15914),
            .in2(_gnd_net_),
            .in3(N__15872),
            .lcout(\b2v_inst.state_17_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22318),
            .ce(),
            .sr(N__22911));
    defparam \b2v_inst.dir_mem_RNO_7_0_LC_9_13_1 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_RNO_7_0_LC_9_13_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNO_7_0_LC_9_13_1 .LUT_INIT=16'b0101111111100000;
    LogicCell40 \b2v_inst.dir_mem_RNO_7_0_LC_9_13_1  (
            .in0(N__19070),
            .in1(N__18982),
            .in2(N__18939),
            .in3(N__19873),
            .lcout(),
            .ltout(\b2v_inst.g4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_RNO_2_0_LC_9_13_2 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_RNO_2_0_LC_9_13_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNO_2_0_LC_9_13_2 .LUT_INIT=16'b0011001011111010;
    LogicCell40 \b2v_inst.dir_mem_RNO_2_0_LC_9_13_2  (
            .in0(N__18773),
            .in1(N__16814),
            .in2(N__16238),
            .in3(N__16301),
            .lcout(\b2v_inst.g0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNIBERF_15_LC_9_13_3 .C_ON=1'b0;
    defparam \b2v_inst.state_RNIBERF_15_LC_9_13_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNIBERF_15_LC_9_13_3 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \b2v_inst.state_RNIBERF_15_LC_9_13_3  (
            .in0(N__18927),
            .in1(N__19048),
            .in2(_gnd_net_),
            .in3(N__18981),
            .lcout(\b2v_inst.N_451 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_15_LC_9_13_4 .C_ON=1'b0;
    defparam \b2v_inst.state_15_LC_9_13_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.state_15_LC_9_13_4 .LUT_INIT=16'b1111111000000000;
    LogicCell40 \b2v_inst.state_15_LC_9_13_4  (
            .in0(N__16228),
            .in1(N__16175),
            .in2(N__16113),
            .in3(N__16037),
            .lcout(\b2v_inst.stateZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22318),
            .ce(),
            .sr(N__22911));
    defparam \b2v_inst.indice_0_rep1_RNI3OC22_LC_9_14_0 .C_ON=1'b0;
    defparam \b2v_inst.indice_0_rep1_RNI3OC22_LC_9_14_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_0_rep1_RNI3OC22_LC_9_14_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst.indice_0_rep1_RNI3OC22_LC_9_14_0  (
            .in0(N__19667),
            .in1(N__17486),
            .in2(N__17398),
            .in3(N__17507),
            .lcout(\b2v_inst.N_410 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_2_RNO_0_3_LC_9_14_1 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_2_RNO_0_3_LC_9_14_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_2_RNO_0_3_LC_9_14_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \b2v_inst.dir_mem_2_RNO_0_3_LC_9_14_1  (
            .in0(N__23083),
            .in1(N__20298),
            .in2(_gnd_net_),
            .in3(N__20117),
            .lcout(),
            .ltout(\b2v_inst.dir_mem_2_RNO_0Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_2_3_LC_9_14_2 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_2_3_LC_9_14_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.dir_mem_2_3_LC_9_14_2 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst.dir_mem_2_3_LC_9_14_2  (
            .in0(_gnd_net_),
            .in1(N__17341),
            .in2(N__15992),
            .in3(N__16733),
            .lcout(\b2v_inst.dir_mem_2Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22502),
            .ce(N__16673),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_3_RNO_0_4_LC_9_14_5 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_3_RNO_0_4_LC_9_14_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_3_RNO_0_4_LC_9_14_5 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \b2v_inst.dir_mem_3_RNO_0_4_LC_9_14_5  (
            .in0(N__23082),
            .in1(N__20297),
            .in2(_gnd_net_),
            .in3(N__20116),
            .lcout(\b2v_inst.un1_dir_mem_3_ns_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_2_7_LC_9_15_0 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_2_7_LC_9_15_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.dir_mem_2_7_LC_9_15_0 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \b2v_inst.dir_mem_2_7_LC_9_15_0  (
            .in0(N__20604),
            .in1(N__20914),
            .in2(N__20500),
            .in3(N__15965),
            .lcout(\b2v_inst.dir_mem_2Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22319),
            .ce(N__16677),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_2_RNO_0_7_LC_9_15_1 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_2_RNO_0_7_LC_9_15_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_2_RNO_0_7_LC_9_15_1 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \b2v_inst.dir_mem_2_RNO_0_7_LC_9_15_1  (
            .in0(N__18391),
            .in1(N__17872),
            .in2(N__20768),
            .in3(N__19673),
            .lcout(\b2v_inst.dir_mem_2_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_2_RNI8NDV_7_LC_9_15_2 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_2_RNI8NDV_7_LC_9_15_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_2_RNI8NDV_7_LC_9_15_2 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \b2v_inst.dir_mem_2_RNI8NDV_7_LC_9_15_2  (
            .in0(N__17013),
            .in1(N__16478),
            .in2(N__16418),
            .in3(N__20913),
            .lcout(),
            .ltout(\b2v_inst.addr_ram_1_0_iv_i_1_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_RNIOPNS2_7_LC_9_15_3 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_RNIOPNS2_7_LC_9_15_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNIOPNS2_7_LC_9_15_3 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \b2v_inst.dir_mem_RNIOPNS2_7_LC_9_15_3  (
            .in0(N__16401),
            .in1(N__19160),
            .in2(N__16349),
            .in3(N__16346),
            .lcout(N_50),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_RNO_8_0_LC_9_15_4 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_RNO_8_0_LC_9_15_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNO_8_0_LC_9_15_4 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \b2v_inst.dir_mem_RNO_8_0_LC_9_15_4  (
            .in0(N__17871),
            .in1(N__20912),
            .in2(N__18395),
            .in3(N__18336),
            .lcout(),
            .ltout(\b2v_inst.g0_2_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_RNO_6_0_LC_9_15_5 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_RNO_6_0_LC_9_15_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNO_6_0_LC_9_15_5 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \b2v_inst.dir_mem_RNO_6_0_LC_9_15_5  (
            .in0(N__18938),
            .in1(N__19082),
            .in2(N__16304),
            .in3(N__20603),
            .lcout(\b2v_inst.g0_2_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_1_RNO_0_6_LC_9_16_0 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_1_RNO_0_6_LC_9_16_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_1_RNO_0_6_LC_9_16_0 .LUT_INIT=16'b0001000000001000;
    LogicCell40 \b2v_inst.dir_mem_1_RNO_0_6_LC_9_16_0  (
            .in0(N__20296),
            .in1(N__18004),
            .in2(N__16565),
            .in3(N__20637),
            .lcout(),
            .ltout(\b2v_inst.i4_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_1_6_LC_9_16_1 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_1_6_LC_9_16_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.dir_mem_1_6_LC_9_16_1 .LUT_INIT=16'b0110011011100100;
    LogicCell40 \b2v_inst.dir_mem_1_6_LC_9_16_1  (
            .in0(N__20494),
            .in1(N__20638),
            .in2(N__16289),
            .in3(N__20933),
            .lcout(\b2v_inst.dir_mem_1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22569),
            .ce(N__19926),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_RNI3ML81_3_LC_9_16_2 .C_ON=1'b0;
    defparam \b2v_inst.indice_RNI3ML81_3_LC_9_16_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_RNI3ML81_3_LC_9_16_2 .LUT_INIT=16'b1111111000000000;
    LogicCell40 \b2v_inst.indice_RNI3ML81_3_LC_9_16_2  (
            .in0(N__20294),
            .in1(N__18002),
            .in2(N__16259),
            .in3(N__20493),
            .lcout(\b2v_inst.un2_dir_mem_3_c5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_3_rep1_RNIS3BN_LC_9_16_3 .C_ON=1'b0;
    defparam \b2v_inst.indice_3_rep1_RNIS3BN_LC_9_16_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_3_rep1_RNIS3BN_LC_9_16_3 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \b2v_inst.indice_3_rep1_RNIS3BN_LC_9_16_3  (
            .in0(N__17116),
            .in1(N__19514),
            .in2(_gnd_net_),
            .in3(N__21174),
            .lcout(\b2v_inst.un2_dir_mem_3_ac0_3 ),
            .ltout(\b2v_inst.un2_dir_mem_3_ac0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_3_RNO_0_5_LC_9_16_4 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_3_RNO_0_5_LC_9_16_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_3_RNO_0_5_LC_9_16_4 .LUT_INIT=16'b0011001100000101;
    LogicCell40 \b2v_inst.dir_mem_3_RNO_0_5_LC_9_16_4  (
            .in0(N__20295),
            .in1(N__20797),
            .in2(N__16250),
            .in3(N__18003),
            .lcout(\b2v_inst.un1_dir_mem_3_ns_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_1_RNO_1_6_LC_9_16_5 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_1_RNO_1_6_LC_9_16_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_1_RNO_1_6_LC_9_16_5 .LUT_INIT=16'b0011000001110001;
    LogicCell40 \b2v_inst.dir_mem_1_RNO_1_6_LC_9_16_5  (
            .in0(N__21092),
            .in1(N__20115),
            .in2(N__18019),
            .in3(N__21176),
            .lcout(\b2v_inst.m7_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_0_rep2_RNI875S_LC_9_16_6 .C_ON=1'b0;
    defparam \b2v_inst.indice_0_rep2_RNI875S_LC_9_16_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_0_rep2_RNI875S_LC_9_16_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst.indice_0_rep2_RNI875S_LC_9_16_6  (
            .in0(N__21175),
            .in1(N__20093),
            .in2(N__20324),
            .in3(N__21091),
            .lcout(\b2v_inst.un8_dir_mem_3_c4 ),
            .ltout(\b2v_inst.un8_dir_mem_3_c4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_3_RNO_0_6_LC_9_16_7 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_3_RNO_0_6_LC_9_16_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_3_RNO_0_6_LC_9_16_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \b2v_inst.dir_mem_3_RNO_0_6_LC_9_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16556),
            .in3(N__20957),
            .lcout(\b2v_inst.un8_dir_mem_3_c6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_2_RNO_0_4_LC_9_17_0 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_2_RNO_0_4_LC_9_17_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_2_RNO_0_4_LC_9_17_0 .LUT_INIT=16'b0100110001001101;
    LogicCell40 \b2v_inst.dir_mem_2_RNO_0_4_LC_9_17_0  (
            .in0(N__20123),
            .in1(N__20330),
            .in2(N__23077),
            .in3(N__21094),
            .lcout(),
            .ltout(\b2v_inst.un2_indice_1_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_2_4_LC_9_17_1 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_2_4_LC_9_17_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.dir_mem_2_4_LC_9_17_1 .LUT_INIT=16'b1110011100011000;
    LogicCell40 \b2v_inst.dir_mem_2_4_LC_9_17_1  (
            .in0(N__20331),
            .in1(N__16725),
            .in2(N__16544),
            .in3(N__18029),
            .lcout(\b2v_inst.dir_mem_2Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22412),
            .ce(N__16678),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_2_1_LC_9_17_2 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_2_1_LC_9_17_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.dir_mem_2_1_LC_9_17_2 .LUT_INIT=16'b0101010110011001;
    LogicCell40 \b2v_inst.dir_mem_2_1_LC_9_17_2  (
            .in0(N__23063),
            .in1(N__23202),
            .in2(_gnd_net_),
            .in3(N__16724),
            .lcout(\b2v_inst.dir_mem_2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22412),
            .ce(N__16678),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_2_2_LC_9_17_3 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_2_2_LC_9_17_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.dir_mem_2_2_LC_9_17_3 .LUT_INIT=16'b0111001011011000;
    LogicCell40 \b2v_inst.dir_mem_2_2_LC_9_17_3  (
            .in0(N__16722),
            .in1(N__20124),
            .in2(N__17471),
            .in3(N__23064),
            .lcout(\b2v_inst.dir_mem_2Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22412),
            .ce(N__16678),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_RNI6V1O2_7_LC_9_17_4 .C_ON=1'b0;
    defparam \b2v_inst.indice_RNI6V1O2_7_LC_9_17_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_RNI6V1O2_7_LC_9_17_4 .LUT_INIT=16'b0000000000010011;
    LogicCell40 \b2v_inst.indice_RNI6V1O2_7_LC_9_17_4  (
            .in0(N__19615),
            .in1(N__18299),
            .in2(N__20666),
            .in3(N__20932),
            .lcout(\b2v_inst.dir_mem_215_0 ),
            .ltout(\b2v_inst.dir_mem_215_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_2_0_LC_9_17_5 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_2_0_LC_9_17_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.dir_mem_2_0_LC_9_17_5 .LUT_INIT=16'b1010010110100101;
    LogicCell40 \b2v_inst.dir_mem_2_0_LC_9_17_5  (
            .in0(N__23201),
            .in1(_gnd_net_),
            .in2(N__16496),
            .in3(_gnd_net_),
            .lcout(\b2v_inst.dir_mem_2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22412),
            .ce(N__16678),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_2_5_LC_9_17_6 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_2_5_LC_9_17_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.dir_mem_2_5_LC_9_17_6 .LUT_INIT=16'b0100011110111000;
    LogicCell40 \b2v_inst.dir_mem_2_5_LC_9_17_6  (
            .in0(N__20664),
            .in1(N__16723),
            .in2(N__17930),
            .in3(N__20502),
            .lcout(\b2v_inst.dir_mem_2Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22412),
            .ce(N__16678),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_SM_Main_ns_2_0__m13_LC_9_18_0 .C_ON=1'b0;
    defparam \b2v_inst1.r_SM_Main_ns_2_0__m13_LC_9_18_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_SM_Main_ns_2_0__m13_LC_9_18_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \b2v_inst1.r_SM_Main_ns_2_0__m13_LC_9_18_0  (
            .in0(_gnd_net_),
            .in1(N__21359),
            .in2(_gnd_net_),
            .in3(N__24020),
            .lcout(\b2v_inst1.N_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_RNIN0GU1_0_LC_10_10_0 .C_ON=1'b1;
    defparam \b2v_inst.dir_mem_RNIN0GU1_0_LC_10_10_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNIN0GU1_0_LC_10_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst.dir_mem_RNIN0GU1_0_LC_10_10_0  (
            .in0(_gnd_net_),
            .in1(N__17773),
            .in2(N__16625),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_10_10_0_),
            .carryout(\b2v_inst.un2_indice_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_RNO_4_1_LC_10_10_1 .C_ON=1'b1;
    defparam \b2v_inst.dir_mem_RNO_4_1_LC_10_10_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNO_4_1_LC_10_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst.dir_mem_RNO_4_1_LC_10_10_1  (
            .in0(_gnd_net_),
            .in1(N__16616),
            .in2(N__17792),
            .in3(N__16610),
            .lcout(\b2v_inst.un2_indice_20_1 ),
            .ltout(),
            .carryin(\b2v_inst.un2_indice_cry_0 ),
            .carryout(\b2v_inst.un2_indice_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_RNO_2_2_LC_10_10_2 .C_ON=1'b1;
    defparam \b2v_inst.dir_mem_RNO_2_2_LC_10_10_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNO_2_2_LC_10_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst.dir_mem_RNO_2_2_LC_10_10_2  (
            .in0(_gnd_net_),
            .in1(N__16607),
            .in2(N__17794),
            .in3(N__16601),
            .lcout(\b2v_inst.un2_indice_20_2 ),
            .ltout(),
            .carryin(\b2v_inst.un2_indice_cry_1 ),
            .carryout(\b2v_inst.un2_indice_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_RNO_2_3_LC_10_10_3 .C_ON=1'b1;
    defparam \b2v_inst.dir_mem_RNO_2_3_LC_10_10_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNO_2_3_LC_10_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst.dir_mem_RNO_2_3_LC_10_10_3  (
            .in0(_gnd_net_),
            .in1(N__16598),
            .in2(N__17793),
            .in3(N__16592),
            .lcout(\b2v_inst.un2_indice_20_3 ),
            .ltout(),
            .carryin(\b2v_inst.un2_indice_cry_2 ),
            .carryout(\b2v_inst.un2_indice_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_RNO_1_4_LC_10_10_4 .C_ON=1'b1;
    defparam \b2v_inst.dir_mem_RNO_1_4_LC_10_10_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNO_1_4_LC_10_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst.dir_mem_RNO_1_4_LC_10_10_4  (
            .in0(_gnd_net_),
            .in1(N__17780),
            .in2(N__16745),
            .in3(N__16589),
            .lcout(\b2v_inst.un2_indice_20_4 ),
            .ltout(),
            .carryin(\b2v_inst.un2_indice_cry_3 ),
            .carryout(\b2v_inst.un2_indice_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_RNO_2_5_LC_10_10_5 .C_ON=1'b1;
    defparam \b2v_inst.dir_mem_RNO_2_5_LC_10_10_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNO_2_5_LC_10_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst.dir_mem_RNO_2_5_LC_10_10_5  (
            .in0(_gnd_net_),
            .in1(N__17786),
            .in2(N__16841),
            .in3(N__16586),
            .lcout(\b2v_inst.un2_indice_20_5 ),
            .ltout(),
            .carryin(\b2v_inst.un2_indice_cry_4 ),
            .carryout(\b2v_inst.un2_indice_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_RNO_1_6_LC_10_10_6 .C_ON=1'b1;
    defparam \b2v_inst.dir_mem_RNO_1_6_LC_10_10_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNO_1_6_LC_10_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst.dir_mem_RNO_1_6_LC_10_10_6  (
            .in0(_gnd_net_),
            .in1(N__17781),
            .in2(N__16583),
            .in3(N__16568),
            .lcout(\b2v_inst.un2_indice_20_6 ),
            .ltout(),
            .carryin(\b2v_inst.un2_indice_cry_5 ),
            .carryout(\b2v_inst.un2_indice_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_RNO_3_7_LC_10_10_7 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_RNO_3_7_LC_10_10_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNO_3_7_LC_10_10_7 .LUT_INIT=16'b0010111011010001;
    LogicCell40 \b2v_inst.dir_mem_RNO_3_7_LC_10_10_7  (
            .in0(N__20935),
            .in1(N__19740),
            .in2(N__19159),
            .in3(N__16775),
            .lcout(\b2v_inst.un2_indice_20_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_1_rep2_LC_10_11_1 .C_ON=1'b0;
    defparam \b2v_inst.indice_1_rep2_LC_10_11_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.indice_1_rep2_LC_10_11_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \b2v_inst.indice_1_rep2_LC_10_11_1  (
            .in0(N__21134),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23166),
            .lcout(\b2v_inst.indice_1_repZ0Z2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21964),
            .ce(N__22951),
            .sr(N__22906));
    defparam \b2v_inst.indice_0_rep2_RNIHJJG_LC_10_11_2 .C_ON=1'b0;
    defparam \b2v_inst.indice_0_rep2_RNIHJJG_LC_10_11_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_0_rep2_RNIHJJG_LC_10_11_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \b2v_inst.indice_0_rep2_RNIHJJG_LC_10_11_2  (
            .in0(_gnd_net_),
            .in1(N__21133),
            .in2(_gnd_net_),
            .in3(N__21058),
            .lcout(\b2v_inst.un2_indice_21_s0_1 ),
            .ltout(\b2v_inst.un2_indice_21_s0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_RNO_2_1_LC_10_11_3 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_RNO_2_1_LC_10_11_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNO_2_1_LC_10_11_3 .LUT_INIT=16'b0011000000000000;
    LogicCell40 \b2v_inst.dir_mem_RNO_2_1_LC_10_11_3  (
            .in0(_gnd_net_),
            .in1(N__18766),
            .in2(N__16772),
            .in3(N__17399),
            .lcout(\b2v_inst.dir_mem_RNO_2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_0_rep2_LC_10_11_4 .C_ON=1'b0;
    defparam \b2v_inst.indice_0_rep2_LC_10_11_4 .SEQ_MODE=4'b1011;
    defparam \b2v_inst.indice_0_rep2_LC_10_11_4 .LUT_INIT=16'b1000111100001111;
    LogicCell40 \b2v_inst.indice_0_rep2_LC_10_11_4  (
            .in0(N__19671),
            .in1(N__21005),
            .in2(N__21085),
            .in3(N__19613),
            .lcout(\b2v_inst.indice_0_repZ0Z2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21964),
            .ce(N__22951),
            .sr(N__22906));
    defparam \b2v_inst.dir_mem_RNO_3_1_LC_10_11_5 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_RNO_3_1_LC_10_11_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNO_3_1_LC_10_11_5 .LUT_INIT=16'b1111111100100000;
    LogicCell40 \b2v_inst.dir_mem_RNO_3_1_LC_10_11_5  (
            .in0(N__17400),
            .in1(N__18767),
            .in2(N__16769),
            .in3(N__16760),
            .lcout(),
            .ltout(\b2v_inst.dir_mem_RNO_3Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_RNO_0_1_LC_10_11_6 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_RNO_0_1_LC_10_11_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNO_0_1_LC_10_11_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst.dir_mem_RNO_0_1_LC_10_11_6  (
            .in0(_gnd_net_),
            .in1(N__16754),
            .in2(N__16748),
            .in3(N__16803),
            .lcout(\b2v_inst.un2_indice_3_iv_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_0_LC_10_11_7 .C_ON=1'b0;
    defparam \b2v_inst.indice_0_LC_10_11_7 .SEQ_MODE=4'b1011;
    defparam \b2v_inst.indice_0_LC_10_11_7 .LUT_INIT=16'b1000000011111111;
    LogicCell40 \b2v_inst.indice_0_LC_10_11_7  (
            .in0(N__21004),
            .in1(N__19672),
            .in2(N__19616),
            .in3(N__23167),
            .lcout(\b2v_inst.indiceZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21964),
            .ce(N__22951),
            .sr(N__22906));
    defparam \b2v_inst.dir_mem_RNIP73H1_4_LC_10_12_0 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_RNIP73H1_4_LC_10_12_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNIP73H1_4_LC_10_12_0 .LUT_INIT=16'b0110011011000011;
    LogicCell40 \b2v_inst.dir_mem_RNIP73H1_4_LC_10_12_0  (
            .in0(N__19357),
            .in1(N__17769),
            .in2(N__17973),
            .in3(N__19724),
            .lcout(\b2v_inst.dir_mem_RNIP73H1Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_4_LC_10_12_1 .C_ON=1'b0;
    defparam \b2v_inst.indice_4_LC_10_12_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.indice_4_LC_10_12_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \b2v_inst.indice_4_LC_10_12_1  (
            .in0(_gnd_net_),
            .in1(N__20822),
            .in2(_gnd_net_),
            .in3(N__17958),
            .lcout(\b2v_inst.indiceZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22280),
            .ce(N__22950),
            .sr(N__22912));
    defparam \b2v_inst.indice_5_LC_10_12_2 .C_ON=1'b0;
    defparam \b2v_inst.indice_5_LC_10_12_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.indice_5_LC_10_12_2 .LUT_INIT=16'b0000000001101010;
    LogicCell40 \b2v_inst.indice_5_LC_10_12_2  (
            .in0(N__20407),
            .in1(N__20824),
            .in2(N__17974),
            .in3(N__21265),
            .lcout(\b2v_inst.indiceZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22280),
            .ce(N__22950),
            .sr(N__22912));
    defparam \b2v_inst.indice_4_rep1_LC_10_12_4 .C_ON=1'b0;
    defparam \b2v_inst.indice_4_rep1_LC_10_12_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.indice_4_rep1_LC_10_12_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \b2v_inst.indice_4_rep1_LC_10_12_4  (
            .in0(N__20823),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21222),
            .lcout(\b2v_inst.indice_4_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22280),
            .ce(N__22950),
            .sr(N__22912));
    defparam \b2v_inst.dir_mem_RNIR93H1_5_LC_10_12_5 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_RNIR93H1_5_LC_10_12_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNIR93H1_5_LC_10_12_5 .LUT_INIT=16'b0111100000101101;
    LogicCell40 \b2v_inst.dir_mem_RNIR93H1_5_LC_10_12_5  (
            .in0(N__19725),
            .in1(N__19256),
            .in2(N__17791),
            .in3(N__20404),
            .lcout(\b2v_inst.dir_mem_RNIR93H1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_RNO_7_6_LC_10_12_6 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_RNO_7_6_LC_10_12_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNO_7_6_LC_10_12_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst.dir_mem_RNO_7_6_LC_10_12_6  (
            .in0(N__20405),
            .in1(N__17108),
            .in2(N__19519),
            .in3(N__21220),
            .lcout(\b2v_inst.g1_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_RNO_5_0_LC_10_12_7 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_RNO_5_0_LC_10_12_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNO_5_0_LC_10_12_7 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \b2v_inst.dir_mem_RNO_5_0_LC_10_12_7  (
            .in0(N__21221),
            .in1(N__18986),
            .in2(N__17117),
            .in3(N__20406),
            .lcout(\b2v_inst.g0_2_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_RNO_0_5_LC_10_13_0 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_RNO_0_5_LC_10_13_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNO_0_5_LC_10_13_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \b2v_inst.dir_mem_RNO_0_5_LC_10_13_0  (
            .in0(_gnd_net_),
            .in1(N__16868),
            .in2(_gnd_net_),
            .in3(N__18764),
            .lcout(),
            .ltout(\b2v_inst.N_411_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_5_LC_10_13_1 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_5_LC_10_13_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.dir_mem_5_LC_10_13_1 .LUT_INIT=16'b1111110111110101;
    LogicCell40 \b2v_inst.dir_mem_5_LC_10_13_1  (
            .in0(N__17303),
            .in1(N__16804),
            .in2(N__16787),
            .in3(N__16784),
            .lcout(\b2v_inst.dir_memZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21945),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_4_rep1_RNI93E71_LC_10_13_2 .C_ON=1'b0;
    defparam \b2v_inst.indice_4_rep1_RNI93E71_LC_10_13_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_4_rep1_RNI93E71_LC_10_13_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst.indice_4_rep1_RNI93E71_LC_10_13_2  (
            .in0(N__20277),
            .in1(N__21206),
            .in2(N__19517),
            .in3(N__21155),
            .lcout(\b2v_inst.un8_dir_mem_2_c4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_3_rep1_RNI4RFQ_LC_10_13_3 .C_ON=1'b0;
    defparam \b2v_inst.indice_3_rep1_RNI4RFQ_LC_10_13_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_3_rep1_RNI4RFQ_LC_10_13_3 .LUT_INIT=16'b1111111000000001;
    LogicCell40 \b2v_inst.indice_3_rep1_RNI4RFQ_LC_10_13_3  (
            .in0(N__21157),
            .in1(N__21084),
            .in2(N__19518),
            .in3(N__17088),
            .lcout(\b2v_inst.un2_indice_21_s0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_RNO_3_5_LC_10_13_4 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_RNO_3_5_LC_10_13_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNO_3_5_LC_10_13_4 .LUT_INIT=16'b0101011011111111;
    LogicCell40 \b2v_inst.dir_mem_RNO_3_5_LC_10_13_4  (
            .in0(N__20403),
            .in1(N__17962),
            .in2(N__16862),
            .in3(N__17380),
            .lcout(\b2v_inst.un2_indice_3_iv_0_a2_2_sx_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_2_rep1_RNIQKCO_LC_10_13_5 .C_ON=1'b0;
    defparam \b2v_inst.indice_2_rep1_RNIQKCO_LC_10_13_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_2_rep1_RNIQKCO_LC_10_13_5 .LUT_INIT=16'b1110111000010001;
    LogicCell40 \b2v_inst.indice_2_rep1_RNIQKCO_LC_10_13_5  (
            .in0(N__21156),
            .in1(N__21083),
            .in2(_gnd_net_),
            .in3(N__19504),
            .lcout(\b2v_inst.un2_indice_21_s0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_4_rep1_RNIP76I_0_LC_10_13_6 .C_ON=1'b0;
    defparam \b2v_inst.indice_4_rep1_RNIP76I_0_LC_10_13_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_4_rep1_RNIP76I_0_LC_10_13_6 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \b2v_inst.indice_4_rep1_RNIP76I_0_LC_10_13_6  (
            .in0(N__20402),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21204),
            .lcout(\b2v_inst.un2_indice_3_0_iv_0_a2_0_8_2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_fast_RNIDAJG_2_LC_10_13_7 .C_ON=1'b0;
    defparam \b2v_inst.indice_fast_RNIDAJG_2_LC_10_13_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_fast_RNIDAJG_2_LC_10_13_7 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \b2v_inst.indice_fast_RNIDAJG_2_LC_10_13_7  (
            .in0(N__21205),
            .in1(N__17087),
            .in2(_gnd_net_),
            .in3(N__18338),
            .lcout(\b2v_inst.indice_fast_RNIDAJGZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_3_rep1_RNI2RFQ_LC_10_14_0 .C_ON=1'b0;
    defparam \b2v_inst.indice_3_rep1_RNI2RFQ_LC_10_14_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_3_rep1_RNI2RFQ_LC_10_14_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \b2v_inst.indice_3_rep1_RNI2RFQ_LC_10_14_0  (
            .in0(N__17112),
            .in1(N__18389),
            .in2(N__19515),
            .in3(N__17873),
            .lcout(\b2v_inst.un2_indice_0_d0_c4_d ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_RNO_5_7_LC_10_14_1 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_RNO_5_7_LC_10_14_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNO_5_7_LC_10_14_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \b2v_inst.dir_mem_RNO_5_7_LC_10_14_1  (
            .in0(_gnd_net_),
            .in1(N__20630),
            .in2(_gnd_net_),
            .in3(N__20441),
            .lcout(),
            .ltout(\b2v_inst.un2_m1_e_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_RNO_2_7_LC_10_14_2 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_RNO_2_7_LC_10_14_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNO_2_7_LC_10_14_2 .LUT_INIT=16'b1110111100010000;
    LogicCell40 \b2v_inst.dir_mem_RNO_2_7_LC_10_14_2  (
            .in0(N__21225),
            .in1(N__16855),
            .in2(N__16844),
            .in3(N__20928),
            .lcout(\b2v_inst.dir_mem_RNO_2Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_0_rep1_LC_10_14_3 .C_ON=1'b0;
    defparam \b2v_inst.indice_0_rep1_LC_10_14_3 .SEQ_MODE=4'b1011;
    defparam \b2v_inst.indice_0_rep1_LC_10_14_3 .LUT_INIT=16'b1101010101010101;
    LogicCell40 \b2v_inst.indice_0_rep1_LC_10_14_3  (
            .in0(N__17875),
            .in1(N__21003),
            .in2(N__19614),
            .in3(N__19665),
            .lcout(\b2v_inst.indice_0_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22281),
            .ce(N__22949),
            .sr(N__22913));
    defparam \b2v_inst.dir_mem_RNO_4_4_LC_10_14_4 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_RNO_4_4_LC_10_14_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNO_4_4_LC_10_14_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst.dir_mem_RNO_4_4_LC_10_14_4  (
            .in0(N__17113),
            .in1(N__18390),
            .in2(N__19516),
            .in3(N__17874),
            .lcout(),
            .ltout(\b2v_inst.dir_mem_RNO_4Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_RNO_2_4_LC_10_14_5 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_RNO_2_4_LC_10_14_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNO_2_4_LC_10_14_5 .LUT_INIT=16'b0011111111110011;
    LogicCell40 \b2v_inst.dir_mem_RNO_2_4_LC_10_14_5  (
            .in0(_gnd_net_),
            .in1(N__17390),
            .in2(N__17048),
            .in3(N__21224),
            .lcout(\b2v_inst.dir_mem_RNO_2Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_3_rep1_LC_10_14_6 .C_ON=1'b0;
    defparam \b2v_inst.indice_3_rep1_LC_10_14_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.indice_3_rep1_LC_10_14_6 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \b2v_inst.indice_3_rep1_LC_10_14_6  (
            .in0(N__20113),
            .in1(N__23036),
            .in2(N__20333),
            .in3(N__23195),
            .lcout(\b2v_inst.indice_3_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22281),
            .ce(N__22949),
            .sr(N__22913));
    defparam \b2v_inst.indice_RNIA33N_1_LC_10_14_7 .C_ON=1'b0;
    defparam \b2v_inst.indice_RNIA33N_1_LC_10_14_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_RNIA33N_1_LC_10_14_7 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \b2v_inst.indice_RNIA33N_1_LC_10_14_7  (
            .in0(N__23037),
            .in1(N__20323),
            .in2(N__23215),
            .in3(N__20114),
            .lcout(\b2v_inst.indice_RNIA33NZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_3_RNIDN331_2_LC_10_15_0 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_3_RNIDN331_2_LC_10_15_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_3_RNIDN331_2_LC_10_15_0 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \b2v_inst.dir_mem_3_RNIDN331_2_LC_10_15_0  (
            .in0(N__17011),
            .in1(N__16957),
            .in2(N__16895),
            .in3(N__20094),
            .lcout(\b2v_inst.addr_ram_1_0_iv_i_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_2_LC_10_15_1 .C_ON=1'b0;
    defparam \b2v_inst.indice_2_LC_10_15_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.indice_2_LC_10_15_1 .LUT_INIT=16'b0000000001101010;
    LogicCell40 \b2v_inst.indice_2_LC_10_15_1  (
            .in0(N__20095),
            .in1(N__23174),
            .in2(N__23076),
            .in3(N__21251),
            .lcout(\b2v_inst.indiceZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21946),
            .ce(N__22947),
            .sr(N__22916));
    defparam \b2v_inst.indice_4_rep1_RNIQ9HI1_LC_10_15_2 .C_ON=1'b0;
    defparam \b2v_inst.indice_4_rep1_RNIQ9HI1_LC_10_15_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_4_rep1_RNIQ9HI1_LC_10_15_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \b2v_inst.indice_4_rep1_RNIQ9HI1_LC_10_15_2  (
            .in0(N__20990),
            .in1(N__19603),
            .in2(_gnd_net_),
            .in3(N__19656),
            .lcout(\b2v_inst.un10_indice ),
            .ltout(\b2v_inst.un10_indice_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_fast_2_LC_10_15_3 .C_ON=1'b0;
    defparam \b2v_inst.indice_fast_2_LC_10_15_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.indice_fast_2_LC_10_15_3 .LUT_INIT=16'b0000011000001100;
    LogicCell40 \b2v_inst.indice_fast_2_LC_10_15_3  (
            .in0(N__23058),
            .in1(N__18337),
            .in2(N__16871),
            .in3(N__23175),
            .lcout(\b2v_inst.indice_fastZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21946),
            .ce(N__22947),
            .sr(N__22916));
    defparam \b2v_inst.indice_fast_3_LC_10_15_5 .C_ON=1'b0;
    defparam \b2v_inst.indice_fast_3_LC_10_15_5 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.indice_fast_3_LC_10_15_5 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \b2v_inst.indice_fast_3_LC_10_15_5  (
            .in0(N__23059),
            .in1(N__20106),
            .in2(N__20329),
            .in3(N__23176),
            .lcout(\b2v_inst.indice_fastZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21946),
            .ce(N__22947),
            .sr(N__22916));
    defparam \b2v_inst.indice_1_rep1_LC_10_15_6 .C_ON=1'b0;
    defparam \b2v_inst.indice_1_rep1_LC_10_15_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.indice_1_rep1_LC_10_15_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \b2v_inst.indice_1_rep1_LC_10_15_6  (
            .in0(N__23173),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18392),
            .lcout(\b2v_inst.indice_1_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21946),
            .ce(N__22947),
            .sr(N__22916));
    defparam \b2v_inst1.r_RX_Byte_RNO_0_2_LC_10_16_1 .C_ON=1'b0;
    defparam \b2v_inst1.r_RX_Byte_RNO_0_2_LC_10_16_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_RX_Byte_RNO_0_2_LC_10_16_1 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \b2v_inst1.r_RX_Byte_RNO_0_2_LC_10_16_1  (
            .in0(N__18090),
            .in1(N__18227),
            .in2(_gnd_net_),
            .in3(N__18193),
            .lcout(\b2v_inst1.r_RX_Bytece_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_Clk_Count_RNO_10_5_LC_10_16_3 .C_ON=1'b0;
    defparam \b2v_inst1.r_Clk_Count_RNO_10_5_LC_10_16_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_Clk_Count_RNO_10_5_LC_10_16_3 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \b2v_inst1.r_Clk_Count_RNO_10_5_LC_10_16_3  (
            .in0(N__23591),
            .in1(N__21467),
            .in2(N__23474),
            .in3(N__21563),
            .lcout(\b2v_inst1.g0_0_i_a6_3_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_Clk_Count_RNI9O3K3_6_LC_10_16_4 .C_ON=1'b0;
    defparam \b2v_inst1.r_Clk_Count_RNI9O3K3_6_LC_10_16_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_Clk_Count_RNI9O3K3_6_LC_10_16_4 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \b2v_inst1.r_Clk_Count_RNI9O3K3_6_LC_10_16_4  (
            .in0(N__24018),
            .in1(N__23749),
            .in2(N__21354),
            .in3(N__23593),
            .lcout(\b2v_inst1.r_RX_Byte_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_Clk_Count_RNO_1_6_LC_10_16_5 .C_ON=1'b0;
    defparam \b2v_inst1.r_Clk_Count_RNO_1_6_LC_10_16_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_Clk_Count_RNO_1_6_LC_10_16_5 .LUT_INIT=16'b0010001100000101;
    LogicCell40 \b2v_inst1.r_Clk_Count_RNO_1_6_LC_10_16_5  (
            .in0(N__23592),
            .in1(N__23445),
            .in2(N__23756),
            .in3(N__24019),
            .lcout(\b2v_inst1.g0_7_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_RX_Byte_RNO_0_0_LC_10_16_7 .C_ON=1'b0;
    defparam \b2v_inst1.r_RX_Byte_RNO_0_0_LC_10_16_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_RX_Byte_RNO_0_0_LC_10_16_7 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \b2v_inst1.r_RX_Byte_RNO_0_0_LC_10_16_7  (
            .in0(N__18089),
            .in1(N__18226),
            .in2(_gnd_net_),
            .in3(N__18192),
            .lcout(\b2v_inst1.r_RX_Bytece_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_SM_Main_2_LC_10_17_0 .C_ON=1'b0;
    defparam \b2v_inst1.r_SM_Main_2_LC_10_17_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst1.r_SM_Main_2_LC_10_17_0 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \b2v_inst1.r_SM_Main_2_LC_10_17_0  (
            .in0(N__23989),
            .in1(N__23738),
            .in2(N__23623),
            .in3(N__21353),
            .lcout(\b2v_inst1.r_SM_MainZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22411),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_Clk_Count_RNO_6_4_LC_10_17_1 .C_ON=1'b0;
    defparam \b2v_inst1.r_Clk_Count_RNO_6_4_LC_10_17_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_Clk_Count_RNO_6_4_LC_10_17_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \b2v_inst1.r_Clk_Count_RNO_6_4_LC_10_17_1  (
            .in0(N__23910),
            .in1(N__23594),
            .in2(_gnd_net_),
            .in3(N__23988),
            .lcout(\b2v_inst1.g0_0_i_a6_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_2_RNO_2_6_LC_10_17_2 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_2_RNO_2_6_LC_10_17_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_2_RNO_2_6_LC_10_17_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \b2v_inst.dir_mem_2_RNO_2_6_LC_10_17_2  (
            .in0(N__17114),
            .in1(N__21158),
            .in2(N__19520),
            .in3(N__21093),
            .lcout(\b2v_inst.un2_dir_mem_2_c4_d ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_Clk_Count_RNO_11_5_LC_10_17_4 .C_ON=1'b0;
    defparam \b2v_inst1.r_Clk_Count_RNO_11_5_LC_10_17_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_Clk_Count_RNO_11_5_LC_10_17_4 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \b2v_inst1.r_Clk_Count_RNO_11_5_LC_10_17_4  (
            .in0(N__23987),
            .in1(N__23603),
            .in2(N__23475),
            .in3(N__23911),
            .lcout(\b2v_inst1.g0_0_i_a6_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_Clk_Count_RNO_3_5_LC_10_17_7 .C_ON=1'b0;
    defparam \b2v_inst1.r_Clk_Count_RNO_3_5_LC_10_17_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_Clk_Count_RNO_3_5_LC_10_17_7 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \b2v_inst1.r_Clk_Count_RNO_3_5_LC_10_17_7  (
            .in0(N__19411),
            .in1(N__22694),
            .in2(N__23625),
            .in3(N__21725),
            .lcout(\b2v_inst1.N_11_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_Clk_Count_1_LC_10_18_0 .C_ON=1'b0;
    defparam \b2v_inst1.r_Clk_Count_1_LC_10_18_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst1.r_Clk_Count_1_LC_10_18_0 .LUT_INIT=16'b1110110011101110;
    LogicCell40 \b2v_inst1.r_Clk_Count_1_LC_10_18_0  (
            .in0(N__21395),
            .in1(N__17204),
            .in2(N__23496),
            .in3(N__18461),
            .lcout(\b2v_inst1.r_Clk_CountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22453),
            .ce(),
            .sr(N__24082));
    defparam \b2v_inst1.r_Clk_Count_RNO_3_6_LC_10_18_1 .C_ON=1'b0;
    defparam \b2v_inst1.r_Clk_Count_RNO_3_6_LC_10_18_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_Clk_Count_RNO_3_6_LC_10_18_1 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \b2v_inst1.r_Clk_Count_RNO_3_6_LC_10_18_1  (
            .in0(N__23837),
            .in1(N__21456),
            .in2(N__21562),
            .in3(N__23918),
            .lcout(),
            .ltout(\b2v_inst1.N_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_Clk_Count_RNO_0_6_LC_10_18_2 .C_ON=1'b0;
    defparam \b2v_inst1.r_Clk_Count_RNO_0_6_LC_10_18_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_Clk_Count_RNO_0_6_LC_10_18_2 .LUT_INIT=16'b1100111110001111;
    LogicCell40 \b2v_inst1.r_Clk_Count_RNO_0_6_LC_10_18_2  (
            .in0(N__21694),
            .in1(N__23919),
            .in2(N__17237),
            .in3(N__23343),
            .lcout(\b2v_inst1.N_11_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_Clk_Count_RNO_7_5_LC_10_18_3 .C_ON=1'b0;
    defparam \b2v_inst1.r_Clk_Count_RNO_7_5_LC_10_18_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_Clk_Count_RNO_7_5_LC_10_18_3 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \b2v_inst1.r_Clk_Count_RNO_7_5_LC_10_18_3  (
            .in0(N__19418),
            .in1(N__22690),
            .in2(_gnd_net_),
            .in3(N__21724),
            .lcout(\b2v_inst1.N_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_Clk_Count_RNI64771_1_LC_10_18_4 .C_ON=1'b0;
    defparam \b2v_inst1.r_Clk_Count_RNI64771_1_LC_10_18_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_Clk_Count_RNI64771_1_LC_10_18_4 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \b2v_inst1.r_Clk_Count_RNI64771_1_LC_10_18_4  (
            .in0(N__21455),
            .in1(N__21552),
            .in2(_gnd_net_),
            .in3(N__23836),
            .lcout(\b2v_inst1.N_9 ),
            .ltout(\b2v_inst1.N_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_Clk_Count_RNO_8_5_LC_10_18_5 .C_ON=1'b0;
    defparam \b2v_inst1.r_Clk_Count_RNO_8_5_LC_10_18_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_Clk_Count_RNO_8_5_LC_10_18_5 .LUT_INIT=16'b1010101010001010;
    LogicCell40 \b2v_inst1.r_Clk_Count_RNO_8_5_LC_10_18_5  (
            .in0(N__17234),
            .in1(N__23342),
            .in2(N__17228),
            .in3(N__21693),
            .lcout(),
            .ltout(\b2v_inst1.N_19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_Clk_Count_RNO_2_5_LC_10_18_6 .C_ON=1'b0;
    defparam \b2v_inst1.r_Clk_Count_RNO_2_5_LC_10_18_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_Clk_Count_RNO_2_5_LC_10_18_6 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \b2v_inst1.r_Clk_Count_RNO_2_5_LC_10_18_6  (
            .in0(N__18287),
            .in1(N__17225),
            .in2(N__17216),
            .in3(N__17213),
            .lcout(\b2v_inst1.g0_0_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_Clk_Count_RNO_2_1_LC_10_19_0 .C_ON=1'b0;
    defparam \b2v_inst1.r_Clk_Count_RNO_2_1_LC_10_19_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_Clk_Count_RNO_2_1_LC_10_19_0 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \b2v_inst1.r_Clk_Count_RNO_2_1_LC_10_19_0  (
            .in0(N__21734),
            .in1(N__23729),
            .in2(N__17198),
            .in3(N__23620),
            .lcout(\b2v_inst1.r_SM_Main_1_sqmuxa_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_Clk_Count_RNO_5_1_LC_10_19_1 .C_ON=1'b0;
    defparam \b2v_inst1.r_Clk_Count_RNO_5_1_LC_10_19_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_Clk_Count_RNO_5_1_LC_10_19_1 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \b2v_inst1.r_Clk_Count_RNO_5_1_LC_10_19_1  (
            .in0(N__19416),
            .in1(N__23316),
            .in2(N__22698),
            .in3(N__21689),
            .lcout(\b2v_inst1.g0_3_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_Clk_Count_RNO_6_5_LC_10_19_2 .C_ON=1'b0;
    defparam \b2v_inst1.r_Clk_Count_RNO_6_5_LC_10_19_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_Clk_Count_RNO_6_5_LC_10_19_2 .LUT_INIT=16'b1010000010000000;
    LogicCell40 \b2v_inst1.r_Clk_Count_RNO_6_5_LC_10_19_2  (
            .in0(N__21690),
            .in1(N__23728),
            .in2(N__23341),
            .in3(N__23619),
            .lcout(),
            .ltout(\b2v_inst1.g0_0_i_a6_2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_Clk_Count_RNO_1_5_LC_10_19_3 .C_ON=1'b0;
    defparam \b2v_inst1.r_Clk_Count_RNO_1_5_LC_10_19_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_Clk_Count_RNO_1_5_LC_10_19_3 .LUT_INIT=16'b1100110011101100;
    LogicCell40 \b2v_inst1.r_Clk_Count_RNO_1_5_LC_10_19_3  (
            .in0(N__17294),
            .in1(N__17288),
            .in2(N__17297),
            .in3(N__18449),
            .lcout(\b2v_inst1.g0_0_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_Clk_Count_RNO_5_5_LC_10_19_4 .C_ON=1'b0;
    defparam \b2v_inst1.r_Clk_Count_RNO_5_5_LC_10_19_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_Clk_Count_RNO_5_5_LC_10_19_4 .LUT_INIT=16'b0010001010101010;
    LogicCell40 \b2v_inst1.r_Clk_Count_RNO_5_5_LC_10_19_4  (
            .in0(N__23915),
            .in1(N__23618),
            .in2(_gnd_net_),
            .in3(N__24003),
            .lcout(\b2v_inst1.g0_0_i_a6_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_Clk_Count_RNO_4_5_LC_10_19_5 .C_ON=1'b0;
    defparam \b2v_inst1.r_Clk_Count_RNO_4_5_LC_10_19_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_Clk_Count_RNO_4_5_LC_10_19_5 .LUT_INIT=16'b0000000100010001;
    LogicCell40 \b2v_inst1.r_Clk_Count_RNO_4_5_LC_10_19_5  (
            .in0(N__23617),
            .in1(N__23705),
            .in2(N__23495),
            .in3(N__23916),
            .lcout(\b2v_inst1.N_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_RNO_0_4_LC_11_11_0 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_RNO_0_4_LC_11_11_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNO_0_4_LC_11_11_0 .LUT_INIT=16'b0101111101001100;
    LogicCell40 \b2v_inst.dir_mem_RNO_0_4_LC_11_11_0  (
            .in0(N__17535),
            .in1(N__17282),
            .in2(N__17429),
            .in3(N__18770),
            .lcout(),
            .ltout(\b2v_inst.un2_indice_3_0_i_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_4_LC_11_11_1 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_4_LC_11_11_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.dir_mem_4_LC_11_11_1 .LUT_INIT=16'b0101000000010000;
    LogicCell40 \b2v_inst.dir_mem_4_LC_11_11_1  (
            .in0(N__18530),
            .in1(N__18771),
            .in2(N__17270),
            .in3(N__17267),
            .lcout(\b2v_inst.dir_memZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21874),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_RNO_1_2_LC_11_11_2 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_RNO_1_2_LC_11_11_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNO_1_2_LC_11_11_2 .LUT_INIT=16'b1011010011110000;
    LogicCell40 \b2v_inst.dir_mem_RNO_1_2_LC_11_11_2  (
            .in0(N__19755),
            .in1(N__19808),
            .in2(N__19212),
            .in3(N__19890),
            .lcout(\b2v_inst.un2_indice_21_s1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_RNO_0_7_LC_11_11_3 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_RNO_0_7_LC_11_11_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNO_0_7_LC_11_11_3 .LUT_INIT=16'b0000010010101110;
    LogicCell40 \b2v_inst.dir_mem_RNO_0_7_LC_11_11_3  (
            .in0(N__18769),
            .in1(N__17411),
            .in2(N__17258),
            .in3(N__17246),
            .lcout(),
            .ltout(\b2v_inst.un2_indice_3_0_iv_0_0_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_7_LC_11_11_4 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_7_LC_11_11_4 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.dir_mem_7_LC_11_11_4 .LUT_INIT=16'b0000000000001101;
    LogicCell40 \b2v_inst.dir_mem_7_LC_11_11_4  (
            .in0(N__17537),
            .in1(N__19091),
            .in2(N__17240),
            .in3(N__18529),
            .lcout(\b2v_inst.dir_memZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21874),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_RNO_0_2_LC_11_11_5 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_RNO_0_2_LC_11_11_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNO_0_2_LC_11_11_5 .LUT_INIT=16'b0000010010101110;
    LogicCell40 \b2v_inst.dir_mem_RNO_0_2_LC_11_11_5  (
            .in0(N__18768),
            .in1(N__17410),
            .in2(N__17467),
            .in3(N__17444),
            .lcout(),
            .ltout(\b2v_inst.un2_indice_3_0_iv_0_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_2_LC_11_11_6 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_2_LC_11_11_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.dir_mem_2_LC_11_11_6 .LUT_INIT=16'b0000000000001101;
    LogicCell40 \b2v_inst.dir_mem_2_LC_11_11_6  (
            .in0(N__17536),
            .in1(N__17438),
            .in2(N__17432),
            .in3(N__18528),
            .lcout(\b2v_inst.dir_memZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21874),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_RNO_3_4_LC_11_11_7 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_RNO_3_4_LC_11_11_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNO_3_4_LC_11_11_7 .LUT_INIT=16'b0011001101100110;
    LogicCell40 \b2v_inst.dir_mem_RNO_3_4_LC_11_11_7  (
            .in0(N__17309),
            .in1(N__19362),
            .in2(_gnd_net_),
            .in3(N__19754),
            .lcout(\b2v_inst.dir_mem_RNO_3Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_RNO_1_3_LC_11_12_0 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_RNO_1_3_LC_11_12_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNO_1_3_LC_11_12_0 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \b2v_inst.dir_mem_RNO_1_3_LC_11_12_0  (
            .in0(N__19315),
            .in1(N__17417),
            .in2(_gnd_net_),
            .in3(N__19199),
            .lcout(\b2v_inst.un2_indice_21_s1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_RNO_3_3_LC_11_12_1 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_RNO_3_3_LC_11_12_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNO_3_3_LC_11_12_1 .LUT_INIT=16'b0100000001000000;
    LogicCell40 \b2v_inst.dir_mem_RNO_3_3_LC_11_12_1  (
            .in0(N__19760),
            .in1(N__19805),
            .in2(N__19889),
            .in3(_gnd_net_),
            .lcout(\b2v_inst.un2_indice_0_d1_c2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_RNO_0_3_LC_11_12_2 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_RNO_0_3_LC_11_12_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNO_0_3_LC_11_12_2 .LUT_INIT=16'b0000001011001110;
    LogicCell40 \b2v_inst.dir_mem_RNO_0_3_LC_11_12_2  (
            .in0(N__17409),
            .in1(N__18772),
            .in2(N__17342),
            .in3(N__17327),
            .lcout(),
            .ltout(\b2v_inst.un2_indice_3_0_iv_0_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_3_LC_11_12_3 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_3_LC_11_12_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.dir_mem_3_LC_11_12_3 .LUT_INIT=16'b0000010000000101;
    LogicCell40 \b2v_inst.dir_mem_3_LC_11_12_3  (
            .in0(N__18527),
            .in1(N__17318),
            .in2(N__17312),
            .in3(N__17534),
            .lcout(\b2v_inst.dir_memZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22081),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_RNO_5_4_LC_11_12_4 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_RNO_5_4_LC_11_12_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNO_5_4_LC_11_12_4 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \b2v_inst.dir_mem_RNO_5_4_LC_11_12_4  (
            .in0(N__19804),
            .in1(N__19198),
            .in2(N__19321),
            .in3(N__19876),
            .lcout(\b2v_inst.dir_mem_RNO_5Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_RNO_1_5_LC_11_12_6 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_RNO_1_5_LC_11_12_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNO_1_5_LC_11_12_6 .LUT_INIT=16'b0101000100010101;
    LogicCell40 \b2v_inst.dir_mem_RNO_1_5_LC_11_12_6  (
            .in0(N__17823),
            .in1(N__17525),
            .in2(N__19385),
            .in3(N__19255),
            .lcout(\b2v_inst.un2_indice_3_iv_0_1_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_1_LC_11_12_7 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_1_LC_11_12_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.dir_mem_1_LC_11_12_7 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \b2v_inst.dir_mem_1_LC_11_12_7  (
            .in0(N__17526),
            .in1(N__17824),
            .in2(N__19685),
            .in3(N__17804),
            .lcout(\b2v_inst.dir_memZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22081),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_RNO_4_0_LC_11_13_0 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_RNO_4_0_LC_11_13_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNO_4_0_LC_11_13_0 .LUT_INIT=16'b0110011000111100;
    LogicCell40 \b2v_inst.dir_mem_RNO_4_0_LC_11_13_0  (
            .in0(N__19894),
            .in1(N__17798),
            .in2(N__21095),
            .in3(N__19756),
            .lcout(),
            .ltout(\b2v_inst.un2_indice_20_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_RNO_1_0_LC_11_13_1 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_RNO_1_0_LC_11_13_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNO_1_0_LC_11_13_1 .LUT_INIT=16'b0000011100000000;
    LogicCell40 \b2v_inst.dir_mem_RNO_1_0_LC_11_13_1  (
            .in0(N__18931),
            .in1(N__17699),
            .in2(N__17588),
            .in3(N__18763),
            .lcout(\b2v_inst.N_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNIN365_15_LC_11_13_2 .C_ON=1'b0;
    defparam \b2v_inst.state_RNIN365_15_LC_11_13_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNIN365_15_LC_11_13_2 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \b2v_inst.state_RNIN365_15_LC_11_13_2  (
            .in0(_gnd_net_),
            .in1(N__18932),
            .in2(_gnd_net_),
            .in3(N__18990),
            .lcout(\b2v_inst.N_228 ),
            .ltout(\b2v_inst.N_228_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_17_rep1_RNIVTJP1_LC_11_13_3 .C_ON=1'b0;
    defparam \b2v_inst.state_17_rep1_RNIVTJP1_LC_11_13_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_17_rep1_RNIVTJP1_LC_11_13_3 .LUT_INIT=16'b0101010011111100;
    LogicCell40 \b2v_inst.state_17_rep1_RNIVTJP1_LC_11_13_3  (
            .in0(N__17573),
            .in1(N__19075),
            .in2(N__17552),
            .in3(N__17549),
            .lcout(\b2v_inst.N_234 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_0_rep1_RNIO9HI1_LC_11_13_4 .C_ON=1'b0;
    defparam \b2v_inst.indice_0_rep1_RNIO9HI1_LC_11_13_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_0_rep1_RNIO9HI1_LC_11_13_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \b2v_inst.indice_0_rep1_RNIO9HI1_LC_11_13_4  (
            .in0(N__19655),
            .in1(N__17482),
            .in2(_gnd_net_),
            .in3(N__17506),
            .lcout(),
            .ltout(\b2v_inst.N_383_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_17_rep1_RNIN75C3_LC_11_13_5 .C_ON=1'b0;
    defparam \b2v_inst.state_17_rep1_RNIN75C3_LC_11_13_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_17_rep1_RNIN75C3_LC_11_13_5 .LUT_INIT=16'b0011000000010000;
    LogicCell40 \b2v_inst.state_17_rep1_RNIN75C3_LC_11_13_5  (
            .in0(N__19071),
            .in1(N__17495),
            .in2(N__17489),
            .in3(N__18762),
            .lcout(\b2v_inst.state_17_rep1_RNIN75CZ0Z3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_0_rep1_RNIEF5S_LC_11_14_0 .C_ON=1'b0;
    defparam \b2v_inst.indice_0_rep1_RNIEF5S_LC_11_14_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_0_rep1_RNIEF5S_LC_11_14_0 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \b2v_inst.indice_0_rep1_RNIEF5S_LC_11_14_0  (
            .in0(N__20867),
            .in1(N__17868),
            .in2(N__18393),
            .in3(N__20557),
            .lcout(\b2v_inst.un2_indice_3_0_iv_0_a2_0_8_3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_fast_RNIHI54_3_LC_11_14_2 .C_ON=1'b0;
    defparam \b2v_inst.indice_fast_RNIHI54_3_LC_11_14_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_fast_RNIHI54_3_LC_11_14_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \b2v_inst.indice_fast_RNIHI54_3_LC_11_14_2  (
            .in0(_gnd_net_),
            .in1(N__20710),
            .in2(_gnd_net_),
            .in3(N__18330),
            .lcout(\b2v_inst.un10_indice_2 ),
            .ltout(\b2v_inst.un10_indice_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_fast_RNI7BF71_4_LC_11_14_3 .C_ON=1'b0;
    defparam \b2v_inst.indice_fast_RNI7BF71_4_LC_11_14_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_fast_RNI7BF71_4_LC_11_14_3 .LUT_INIT=16'b1011111110001100;
    LogicCell40 \b2v_inst.indice_fast_RNI7BF71_4_LC_11_14_3  (
            .in0(N__20756),
            .in1(N__17834),
            .in2(N__18056),
            .in3(N__18053),
            .lcout(\b2v_inst.dir_mem_115lto6_1 ),
            .ltout(\b2v_inst.dir_mem_115lto6_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_1_RNO_0_7_LC_11_14_4 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_1_RNO_0_7_LC_11_14_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_1_RNO_0_7_LC_11_14_4 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \b2v_inst.dir_mem_1_RNO_0_7_LC_11_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18047),
            .in3(N__20192),
            .lcout(),
            .ltout(\b2v_inst.un1_dir_mem_1_mb_1_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_1_7_LC_11_14_5 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_1_7_LC_11_14_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.dir_mem_1_7_LC_11_14_5 .LUT_INIT=16'b1010101001010100;
    LogicCell40 \b2v_inst.dir_mem_1_7_LC_11_14_5  (
            .in0(N__19588),
            .in1(N__20180),
            .in2(N__18044),
            .in3(N__20868),
            .lcout(\b2v_inst.dir_mem_1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22082),
            .ce(N__19933),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_2_RNO_0_5_LC_11_15_0 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_2_RNO_0_5_LC_11_15_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_2_RNO_0_5_LC_11_15_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \b2v_inst.dir_mem_2_RNO_0_5_LC_11_15_0  (
            .in0(N__18018),
            .in1(N__20096),
            .in2(N__20027),
            .in3(N__20325),
            .lcout(\b2v_inst.un2_dir_mem_2_c5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_1_RNO_2_4_LC_11_15_1 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_1_RNO_2_4_LC_11_15_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_1_RNO_2_4_LC_11_15_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \b2v_inst.dir_mem_1_RNO_2_4_LC_11_15_1  (
            .in0(_gnd_net_),
            .in1(N__21172),
            .in2(_gnd_net_),
            .in3(N__21090),
            .lcout(),
            .ltout(\b2v_inst.N_4_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_1_RNO_0_4_LC_11_15_2 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_1_RNO_0_4_LC_11_15_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_1_RNO_0_4_LC_11_15_2 .LUT_INIT=16'b1011111111111111;
    LogicCell40 \b2v_inst.dir_mem_1_RNO_0_4_LC_11_15_2  (
            .in0(N__20898),
            .in1(N__20097),
            .in2(N__17915),
            .in3(N__20326),
            .lcout(\b2v_inst.N_8_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_0_rep1_RNIATP21_LC_11_15_3 .C_ON=1'b0;
    defparam \b2v_inst.indice_0_rep1_RNIATP21_LC_11_15_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_0_rep1_RNIATP21_LC_11_15_3 .LUT_INIT=16'b0000000000010011;
    LogicCell40 \b2v_inst.indice_0_rep1_RNIATP21_LC_11_15_3  (
            .in0(N__17870),
            .in1(N__20897),
            .in2(N__18394),
            .in3(N__21223),
            .lcout(),
            .ltout(\b2v_inst.dir_mem_315lto8_a0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_fast_RNIRFV61_3_LC_11_15_4 .C_ON=1'b0;
    defparam \b2v_inst.indice_fast_RNIRFV61_3_LC_11_15_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_fast_RNIRFV61_3_LC_11_15_4 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \b2v_inst.indice_fast_RNIRFV61_3_LC_11_15_4  (
            .in0(_gnd_net_),
            .in1(N__20712),
            .in2(N__17903),
            .in3(N__18332),
            .lcout(\b2v_inst.indice_fast_RNIRFV61Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_0_rep1_RNIFJJG_LC_11_15_5 .C_ON=1'b0;
    defparam \b2v_inst.indice_0_rep1_RNIFJJG_LC_11_15_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_0_rep1_RNIFJJG_LC_11_15_5 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \b2v_inst.indice_0_rep1_RNIFJJG_LC_11_15_5  (
            .in0(N__17869),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18381),
            .lcout(\b2v_inst.indice_0_rep1_RNIFJJGZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_fast_RNIJ9NJ_3_LC_11_15_6 .C_ON=1'b0;
    defparam \b2v_inst.indice_fast_RNIJ9NJ_3_LC_11_15_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_fast_RNIJ9NJ_3_LC_11_15_6 .LUT_INIT=16'b1000000000000001;
    LogicCell40 \b2v_inst.indice_fast_RNIJ9NJ_3_LC_11_15_6  (
            .in0(N__18382),
            .in1(N__20711),
            .in2(N__20763),
            .in3(N__18331),
            .lcout(),
            .ltout(\b2v_inst.dir_mem_215lt6_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_RNIG39V_6_LC_11_15_7 .C_ON=1'b0;
    defparam \b2v_inst.indice_RNIG39V_6_LC_11_15_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_RNIG39V_6_LC_11_15_7 .LUT_INIT=16'b0000110000000000;
    LogicCell40 \b2v_inst.indice_RNIG39V_6_LC_11_15_7  (
            .in0(_gnd_net_),
            .in1(N__20453),
            .in2(N__18302),
            .in3(N__20561),
            .lcout(\b2v_inst.dir_mem_215lt8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_Clk_Count_RNO_9_5_LC_11_16_0 .C_ON=1'b0;
    defparam \b2v_inst1.r_Clk_Count_RNO_9_5_LC_11_16_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_Clk_Count_RNO_9_5_LC_11_16_0 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \b2v_inst1.r_Clk_Count_RNO_9_5_LC_11_16_0  (
            .in0(N__21657),
            .in1(N__24016),
            .in2(N__23344),
            .in3(N__23832),
            .lcout(\b2v_inst1.g0_0_i_a6_3_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_Clk_Count_RNO_0_3_LC_11_16_2 .C_ON=1'b0;
    defparam \b2v_inst1.r_Clk_Count_RNO_0_3_LC_11_16_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_Clk_Count_RNO_0_3_LC_11_16_2 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \b2v_inst1.r_Clk_Count_RNO_0_3_LC_11_16_2  (
            .in0(N__21560),
            .in1(_gnd_net_),
            .in2(N__21476),
            .in3(N__23833),
            .lcout(\b2v_inst1.un1_r_Clk_Count_ac0_3_out ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_SM_Main_ns_2_0__m16_e_LC_11_16_3 .C_ON=1'b0;
    defparam \b2v_inst1.r_SM_Main_ns_2_0__m16_e_LC_11_16_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_SM_Main_ns_2_0__m16_e_LC_11_16_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \b2v_inst1.r_SM_Main_ns_2_0__m16_e_LC_11_16_3  (
            .in0(N__18224),
            .in1(N__18088),
            .in2(_gnd_net_),
            .in3(N__18186),
            .lcout(\b2v_inst1.r_rx_byteZ0Z_7 ),
            .ltout(\b2v_inst1.r_rx_byteZ0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_SM_Main_ns_2_0__m17_LC_11_16_4 .C_ON=1'b0;
    defparam \b2v_inst1.r_SM_Main_ns_2_0__m17_LC_11_16_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_SM_Main_ns_2_0__m17_LC_11_16_4 .LUT_INIT=16'b1001100011001100;
    LogicCell40 \b2v_inst1.r_SM_Main_ns_2_0__m17_LC_11_16_4  (
            .in0(N__21351),
            .in1(N__23741),
            .in2(N__18263),
            .in3(N__24017),
            .lcout(\b2v_inst1.N_32_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_Clk_Count_RNO_4_6_LC_11_16_5 .C_ON=1'b0;
    defparam \b2v_inst1.r_Clk_Count_RNO_4_6_LC_11_16_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_Clk_Count_RNO_4_6_LC_11_16_5 .LUT_INIT=16'b1011101111111111;
    LogicCell40 \b2v_inst1.r_Clk_Count_RNO_4_6_LC_11_16_5  (
            .in0(N__20339),
            .in1(N__21463),
            .in2(_gnd_net_),
            .in3(N__21559),
            .lcout(\b2v_inst1.N_10_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_Bit_Index_2_LC_11_16_6 .C_ON=1'b0;
    defparam \b2v_inst1.r_Bit_Index_2_LC_11_16_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst1.r_Bit_Index_2_LC_11_16_6 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \b2v_inst1.r_Bit_Index_2_LC_11_16_6  (
            .in0(N__21311),
            .in1(N__18225),
            .in2(N__18194),
            .in3(N__18103),
            .lcout(\b2v_inst1.r_Bit_IndexZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22455),
            .ce(),
            .sr(N__24081));
    defparam \b2v_inst1.r_Bit_Index_1_LC_11_16_7 .C_ON=1'b0;
    defparam \b2v_inst1.r_Bit_Index_1_LC_11_16_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst1.r_Bit_Index_1_LC_11_16_7 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \b2v_inst1.r_Bit_Index_1_LC_11_16_7  (
            .in0(N__18102),
            .in1(N__18187),
            .in2(_gnd_net_),
            .in3(N__21310),
            .lcout(\b2v_inst1.r_Bit_IndexZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22455),
            .ce(),
            .sr(N__24081));
    defparam \b2v_inst1.r_Clk_Count_RNO_0_5_LC_11_17_0 .C_ON=1'b0;
    defparam \b2v_inst1.r_Clk_Count_RNO_0_5_LC_11_17_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_Clk_Count_RNO_0_5_LC_11_17_0 .LUT_INIT=16'b1110111101001111;
    LogicCell40 \b2v_inst1.r_Clk_Count_RNO_0_5_LC_11_17_0  (
            .in0(N__21661),
            .in1(N__18455),
            .in2(N__23351),
            .in3(N__18448),
            .lcout(\b2v_inst1.N_14_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_SM_Main_ns_2_0__m22_ns_1_LC_11_17_1 .C_ON=1'b0;
    defparam \b2v_inst1.r_SM_Main_ns_2_0__m22_ns_1_LC_11_17_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_SM_Main_ns_2_0__m22_ns_1_LC_11_17_1 .LUT_INIT=16'b0111011100001100;
    LogicCell40 \b2v_inst1.r_SM_Main_ns_2_0__m22_ns_1_LC_11_17_1  (
            .in0(N__23992),
            .in1(N__23727),
            .in2(N__22709),
            .in3(N__23589),
            .lcout(\b2v_inst1.m22_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_Clk_Count_RNO_9_4_LC_11_17_2 .C_ON=1'b0;
    defparam \b2v_inst1.r_Clk_Count_RNO_9_4_LC_11_17_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_Clk_Count_RNO_9_4_LC_11_17_2 .LUT_INIT=16'b0111001011111010;
    LogicCell40 \b2v_inst1.r_Clk_Count_RNO_9_4_LC_11_17_2  (
            .in0(N__23588),
            .in1(N__23903),
            .in2(N__23748),
            .in3(N__23991),
            .lcout(\b2v_inst1.N_9_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_SM_Main_ns_2_0__m2_0_LC_11_17_3 .C_ON=1'b0;
    defparam \b2v_inst1.r_SM_Main_ns_2_0__m2_0_LC_11_17_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_SM_Main_ns_2_0__m2_0_LC_11_17_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst1.r_SM_Main_ns_2_0__m2_0_LC_11_17_3  (
            .in0(_gnd_net_),
            .in1(N__21439),
            .in2(_gnd_net_),
            .in3(N__21527),
            .lcout(\b2v_inst1.un1_r_Clk_Count_ac0_1_out ),
            .ltout(\b2v_inst1.un1_r_Clk_Count_ac0_1_out_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_SM_Main_ns_2_0__m6_LC_11_17_4 .C_ON=1'b0;
    defparam \b2v_inst1.r_SM_Main_ns_2_0__m6_LC_11_17_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_SM_Main_ns_2_0__m6_LC_11_17_4 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \b2v_inst1.r_SM_Main_ns_2_0__m6_LC_11_17_4  (
            .in0(N__21660),
            .in1(N__19415),
            .in2(N__18437),
            .in3(N__23315),
            .lcout(\b2v_inst1.N_29_mux ),
            .ltout(\b2v_inst1.N_29_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_SM_Main_1_LC_11_17_5 .C_ON=1'b0;
    defparam \b2v_inst1.r_SM_Main_1_LC_11_17_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst1.r_SM_Main_1_LC_11_17_5 .LUT_INIT=16'b1110111010100000;
    LogicCell40 \b2v_inst1.r_SM_Main_1_LC_11_17_5  (
            .in0(N__18434),
            .in1(N__21352),
            .in2(N__18428),
            .in3(N__23590),
            .lcout(\b2v_inst1.r_SM_MainZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22561),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_SM_Main_ns_2_0__m10_LC_11_17_6 .C_ON=1'b0;
    defparam \b2v_inst1.r_SM_Main_ns_2_0__m10_LC_11_17_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_SM_Main_ns_2_0__m10_LC_11_17_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst1.r_SM_Main_ns_2_0__m10_LC_11_17_6  (
            .in0(N__21528),
            .in1(N__23902),
            .in2(N__21462),
            .in3(N__23820),
            .lcout(),
            .ltout(\b2v_inst1.N_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_SM_Main_ns_2_0__m12_LC_11_17_7 .C_ON=1'b0;
    defparam \b2v_inst1.r_SM_Main_ns_2_0__m12_LC_11_17_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_SM_Main_ns_2_0__m12_LC_11_17_7 .LUT_INIT=16'b0101010101000111;
    LogicCell40 \b2v_inst1.r_SM_Main_ns_2_0__m12_LC_11_17_7  (
            .in0(N__23904),
            .in1(N__23347),
            .in2(N__18425),
            .in3(N__21659),
            .lcout(\b2v_inst1.N_28_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_Clk_Count_5_LC_11_18_1 .C_ON=1'b0;
    defparam \b2v_inst1.r_Clk_Count_5_LC_11_18_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst1.r_Clk_Count_5_LC_11_18_1 .LUT_INIT=16'b0000010100000001;
    LogicCell40 \b2v_inst1.r_Clk_Count_5_LC_11_18_1  (
            .in0(N__18422),
            .in1(N__18413),
            .in2(N__18407),
            .in3(N__23901),
            .lcout(\b2v_inst1.r_Clk_CountZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22550),
            .ce(),
            .sr(N__24093));
    defparam \b2v_inst1.r_SM_Main_ns_2_0__m6_2_LC_11_18_3 .C_ON=1'b0;
    defparam \b2v_inst1.r_SM_Main_ns_2_0__m6_2_LC_11_18_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_SM_Main_ns_2_0__m6_2_LC_11_18_3 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \b2v_inst1.r_SM_Main_ns_2_0__m6_2_LC_11_18_3  (
            .in0(N__23984),
            .in1(N__23900),
            .in2(_gnd_net_),
            .in3(N__23809),
            .lcout(\b2v_inst1.m6_2 ),
            .ltout(\b2v_inst1.m6_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_SM_Main_ns_2_0__g0_6_LC_11_18_4 .C_ON=1'b0;
    defparam \b2v_inst1.r_SM_Main_ns_2_0__g0_6_LC_11_18_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_SM_Main_ns_2_0__g0_6_LC_11_18_4 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \b2v_inst1.r_SM_Main_ns_2_0__g0_6_LC_11_18_4  (
            .in0(N__21656),
            .in1(N__23285),
            .in2(N__18512),
            .in3(N__21723),
            .lcout(\b2v_inst1.N_29_mux_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_Clk_Count_RNO_2_6_LC_11_18_5 .C_ON=1'b0;
    defparam \b2v_inst1.r_Clk_Count_RNO_2_6_LC_11_18_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_Clk_Count_RNO_2_6_LC_11_18_5 .LUT_INIT=16'b0101010100100000;
    LogicCell40 \b2v_inst1.r_Clk_Count_RNO_2_6_LC_11_18_5  (
            .in0(N__23985),
            .in1(N__23612),
            .in2(N__23742),
            .in3(N__18509),
            .lcout(),
            .ltout(\b2v_inst1.g0_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_Clk_Count_6_LC_11_18_6 .C_ON=1'b0;
    defparam \b2v_inst1.r_Clk_Count_6_LC_11_18_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst1.r_Clk_Count_6_LC_11_18_6 .LUT_INIT=16'b0000001100001011;
    LogicCell40 \b2v_inst1.r_Clk_Count_6_LC_11_18_6  (
            .in0(N__23613),
            .in1(N__18500),
            .in2(N__18488),
            .in3(N__18485),
            .lcout(\b2v_inst1.r_Clk_CountZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22550),
            .ce(),
            .sr(N__24093));
    defparam \b2v_inst1.r_SM_Main_ns_2_0__m9_LC_11_19_1 .C_ON=1'b0;
    defparam \b2v_inst1.r_SM_Main_ns_2_0__m9_LC_11_19_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_SM_Main_ns_2_0__m9_LC_11_19_1 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \b2v_inst1.r_SM_Main_ns_2_0__m9_LC_11_19_1  (
            .in0(N__23708),
            .in1(_gnd_net_),
            .in2(N__22699),
            .in3(N__21767),
            .lcout(),
            .ltout(\b2v_inst1.N_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_SM_Main_0_LC_11_19_2 .C_ON=1'b0;
    defparam \b2v_inst1.r_SM_Main_0_LC_11_19_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst1.r_SM_Main_0_LC_11_19_2 .LUT_INIT=16'b0100010000000101;
    LogicCell40 \b2v_inst1.r_SM_Main_0_LC_11_19_2  (
            .in0(N__23482),
            .in1(N__18476),
            .in2(N__18467),
            .in3(N__23622),
            .lcout(\b2v_inst1.r_SM_MainZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22510),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_Clk_Count_RNIAI9K1_1_LC_11_19_4 .C_ON=1'b0;
    defparam \b2v_inst1.r_Clk_Count_RNIAI9K1_1_LC_11_19_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_Clk_Count_RNIAI9K1_1_LC_11_19_4 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \b2v_inst1.r_Clk_Count_RNIAI9K1_1_LC_11_19_4  (
            .in0(N__21443),
            .in1(N__21532),
            .in2(N__21695),
            .in3(N__23821),
            .lcout(\b2v_inst1.N_11_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_Clk_Count_RNO_3_1_LC_11_19_5 .C_ON=1'b0;
    defparam \b2v_inst1.r_Clk_Count_RNO_3_1_LC_11_19_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_Clk_Count_RNO_3_1_LC_11_19_5 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \b2v_inst1.r_Clk_Count_RNO_3_1_LC_11_19_5  (
            .in0(N__21533),
            .in1(N__23762),
            .in2(N__21692),
            .in3(N__21444),
            .lcout(),
            .ltout(\b2v_inst1.g2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_Clk_Count_RNO_0_1_LC_11_19_6 .C_ON=1'b0;
    defparam \b2v_inst1.r_Clk_Count_RNO_0_1_LC_11_19_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_Clk_Count_RNO_0_1_LC_11_19_6 .LUT_INIT=16'b1010101011110011;
    LogicCell40 \b2v_inst1.r_Clk_Count_RNO_0_1_LC_11_19_6  (
            .in0(N__21578),
            .in1(N__23707),
            .in2(N__18464),
            .in3(N__23621),
            .lcout(\b2v_inst1.g2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_Clk_Count_RNO_0_4_LC_11_19_7 .C_ON=1'b0;
    defparam \b2v_inst1.r_Clk_Count_RNO_0_4_LC_11_19_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_Clk_Count_RNO_0_4_LC_11_19_7 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \b2v_inst1.r_Clk_Count_RNO_0_4_LC_11_19_7  (
            .in0(N__22679),
            .in1(N__19417),
            .in2(_gnd_net_),
            .in3(N__21733),
            .lcout(\b2v_inst1.N_7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_12_11_0.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_12_11_0.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_12_11_0.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_12_11_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_RNO_4_5_LC_12_12_1 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_RNO_4_5_LC_12_12_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNO_4_5_LC_12_12_1 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \b2v_inst.dir_mem_RNO_4_5_LC_12_12_1  (
            .in0(N__19301),
            .in1(N__19200),
            .in2(N__19331),
            .in3(N__19757),
            .lcout(\b2v_inst.un2_indice_0_d1_c5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_RNIJMO11_4_LC_12_12_2 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_RNIJMO11_4_LC_12_12_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNIJMO11_4_LC_12_12_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \b2v_inst.dir_mem_RNIJMO11_4_LC_12_12_2  (
            .in0(N__19361),
            .in1(N__19806),
            .in2(_gnd_net_),
            .in3(N__19874),
            .lcout(\b2v_inst.un2_indice_0_d1_ac0_7_s_0_0 ),
            .ltout(\b2v_inst.un2_indice_0_d1_ac0_7_s_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_RNO_4_7_LC_12_12_3 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_RNO_4_7_LC_12_12_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNO_4_7_LC_12_12_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst.dir_mem_RNO_4_7_LC_12_12_3  (
            .in0(N__19302),
            .in1(N__19265),
            .in2(N__19220),
            .in3(N__19201),
            .lcout(),
            .ltout(\b2v_inst.un2_indice_0_d1_ac0_9_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_RNO_1_7_LC_12_12_4 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_RNO_1_7_LC_12_12_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNO_1_7_LC_12_12_4 .LUT_INIT=16'b1001110011001100;
    LogicCell40 \b2v_inst.dir_mem_RNO_1_7_LC_12_12_4  (
            .in0(N__19759),
            .in1(N__19149),
            .in2(N__19130),
            .in3(N__19126),
            .lcout(\b2v_inst.un2_indice_21_s1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNIVTJP1_15_LC_12_12_5 .C_ON=1'b0;
    defparam \b2v_inst.state_RNIVTJP1_15_LC_12_12_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNIVTJP1_15_LC_12_12_5 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \b2v_inst.state_RNIVTJP1_15_LC_12_12_5  (
            .in0(N__19081),
            .in1(N__18997),
            .in2(N__18940),
            .in3(N__18765),
            .lcout(),
            .ltout(\b2v_inst.N_384_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.state_RNIM5P55_15_LC_12_12_6 .C_ON=1'b0;
    defparam \b2v_inst.state_RNIM5P55_15_LC_12_12_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.state_RNIM5P55_15_LC_12_12_6 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \b2v_inst.state_RNIM5P55_15_LC_12_12_6  (
            .in0(_gnd_net_),
            .in1(N__18552),
            .in2(N__18539),
            .in3(N__18536),
            .lcout(\b2v_inst.un2_indice_3_0_iv_0_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_RNO_1_1_LC_12_12_7 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_RNO_1_1_LC_12_12_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_RNO_1_1_LC_12_12_7 .LUT_INIT=16'b1100110001100110;
    LogicCell40 \b2v_inst.dir_mem_RNO_1_1_LC_12_12_7  (
            .in0(N__19875),
            .in1(N__19807),
            .in2(_gnd_net_),
            .in3(N__19758),
            .lcout(\b2v_inst.un2_indice_21_s1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_fast_0_LC_12_13_0 .C_ON=1'b0;
    defparam \b2v_inst.indice_fast_0_LC_12_13_0 .SEQ_MODE=4'b1011;
    defparam \b2v_inst.indice_fast_0_LC_12_13_0 .LUT_INIT=16'b1011001100110011;
    LogicCell40 \b2v_inst.indice_fast_0_LC_12_13_0  (
            .in0(N__19587),
            .in1(N__19550),
            .in2(N__21002),
            .in3(N__19666),
            .lcout(\b2v_inst.indice_fastZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22102),
            .ce(N__22948),
            .sr(N__22917));
    defparam \b2v_inst.indice_RNITPHB_6_LC_12_13_1 .C_ON=1'b0;
    defparam \b2v_inst.indice_RNITPHB_6_LC_12_13_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_RNITPHB_6_LC_12_13_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst.indice_RNITPHB_6_LC_12_13_1  (
            .in0(_gnd_net_),
            .in1(N__20617),
            .in2(_gnd_net_),
            .in3(N__20476),
            .lcout(\b2v_inst.CO1 ),
            .ltout(\b2v_inst.CO1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_2_rep1_RNI6ULR_LC_12_13_2 .C_ON=1'b0;
    defparam \b2v_inst.indice_2_rep1_RNI6ULR_LC_12_13_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_2_rep1_RNI6ULR_LC_12_13_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst.indice_2_rep1_RNI6ULR_LC_12_13_2  (
            .in0(N__19467),
            .in1(N__20685),
            .in2(N__19556),
            .in3(N__20019),
            .lcout(\b2v_inst.un8_dir_mem_1_c7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_fast_RNIDE54_0_LC_12_13_3 .C_ON=1'b0;
    defparam \b2v_inst.indice_fast_RNIDE54_0_LC_12_13_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_fast_RNIDE54_0_LC_12_13_3 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \b2v_inst.indice_fast_RNIDE54_0_LC_12_13_3  (
            .in0(N__19549),
            .in1(_gnd_net_),
            .in2(N__19538),
            .in3(_gnd_net_),
            .lcout(\b2v_inst.un2_dir_mem_2_c2 ),
            .ltout(\b2v_inst.un2_dir_mem_2_c2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_1_RNO_0_5_LC_12_13_4 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_1_RNO_0_5_LC_12_13_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_1_RNO_0_5_LC_12_13_4 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \b2v_inst.dir_mem_1_RNO_0_5_LC_12_13_4  (
            .in0(N__20477),
            .in1(N__19472),
            .in2(N__19553),
            .in3(N__20686),
            .lcout(\b2v_inst.dir_mem_1_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_fast_RNIF91E_0_LC_12_13_5 .C_ON=1'b0;
    defparam \b2v_inst.indice_fast_RNIF91E_0_LC_12_13_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_fast_RNIF91E_0_LC_12_13_5 .LUT_INIT=16'b0011011111111111;
    LogicCell40 \b2v_inst.indice_fast_RNIF91E_0_LC_12_13_5  (
            .in0(N__19548),
            .in1(N__19466),
            .in2(N__19537),
            .in3(N__20723),
            .lcout(\b2v_inst.indice_fast_RNIF91EZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_fast_1_LC_12_13_6 .C_ON=1'b0;
    defparam \b2v_inst.indice_fast_1_LC_12_13_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.indice_fast_1_LC_12_13_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \b2v_inst.indice_fast_1_LC_12_13_6  (
            .in0(_gnd_net_),
            .in1(N__23206),
            .in2(_gnd_net_),
            .in3(N__19536),
            .lcout(\b2v_inst.indice_fastZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22102),
            .ce(N__22948),
            .sr(N__22917));
    defparam \b2v_inst.indice_2_rep1_LC_12_13_7 .C_ON=1'b0;
    defparam \b2v_inst.indice_2_rep1_LC_12_13_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.indice_2_rep1_LC_12_13_7 .LUT_INIT=16'b0001001100100000;
    LogicCell40 \b2v_inst.indice_2_rep1_LC_12_13_7  (
            .in0(N__23021),
            .in1(N__21266),
            .in2(N__23217),
            .in3(N__19468),
            .lcout(\b2v_inst.indice_2_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22102),
            .ce(N__22948),
            .sr(N__22917));
    defparam \b2v_inst.dir_mem_1_RNO_0_3_LC_12_14_0 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_1_RNO_0_3_LC_12_14_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_1_RNO_0_3_LC_12_14_0 .LUT_INIT=16'b0011011011001100;
    LogicCell40 \b2v_inst.dir_mem_1_RNO_0_3_LC_12_14_0  (
            .in0(N__23022),
            .in1(N__20327),
            .in2(N__23216),
            .in3(N__20141),
            .lcout(),
            .ltout(\b2v_inst.dir_mem_1_RNO_0Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_1_3_LC_12_14_1 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_1_3_LC_12_14_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.dir_mem_1_3_LC_12_14_1 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \b2v_inst.dir_mem_1_3_LC_12_14_1  (
            .in0(N__20328),
            .in1(_gnd_net_),
            .in2(N__20213),
            .in3(N__19963),
            .lcout(\b2v_inst.dir_mem_1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22388),
            .ce(N__19934),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_fast_RNI6ULR_4_LC_12_14_2 .C_ON=1'b0;
    defparam \b2v_inst.indice_fast_RNI6ULR_4_LC_12_14_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_fast_RNI6ULR_4_LC_12_14_2 .LUT_INIT=16'b0111001110111111;
    LogicCell40 \b2v_inst.indice_fast_RNI6ULR_4_LC_12_14_2  (
            .in0(N__20198),
            .in1(N__20579),
            .in2(N__20764),
            .in3(N__20484),
            .lcout(\b2v_inst.dir_mem_115lto8_1 ),
            .ltout(\b2v_inst.dir_mem_115lto8_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_RNI36K43_7_LC_12_14_3 .C_ON=1'b0;
    defparam \b2v_inst.indice_RNI36K43_7_LC_12_14_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_RNI36K43_7_LC_12_14_3 .LUT_INIT=16'b0000000000110001;
    LogicCell40 \b2v_inst.indice_RNI36K43_7_LC_12_14_3  (
            .in0(N__20186),
            .in1(N__20179),
            .in2(N__20168),
            .in3(N__20927),
            .lcout(\b2v_inst.dir_mem_115_0 ),
            .ltout(\b2v_inst.dir_mem_115_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_1_0_LC_12_14_4 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_1_0_LC_12_14_4 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.dir_mem_1_0_LC_12_14_4 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \b2v_inst.dir_mem_1_0_LC_12_14_4  (
            .in0(N__23199),
            .in1(_gnd_net_),
            .in2(N__20165),
            .in3(_gnd_net_),
            .lcout(\b2v_inst.dir_mem_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22388),
            .ce(N__19934),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_1_2_LC_12_14_5 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_1_2_LC_12_14_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.dir_mem_1_2_LC_12_14_5 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \b2v_inst.dir_mem_1_2_LC_12_14_5  (
            .in0(N__20142),
            .in1(N__20020),
            .in2(_gnd_net_),
            .in3(N__19962),
            .lcout(\b2v_inst.dir_mem_1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22388),
            .ce(N__19934),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_1_5_LC_12_14_6 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_1_5_LC_12_14_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.dir_mem_1_5_LC_12_14_6 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \b2v_inst.dir_mem_1_5_LC_12_14_6  (
            .in0(N__19964),
            .in1(N__19985),
            .in2(_gnd_net_),
            .in3(N__20485),
            .lcout(\b2v_inst.dir_mem_1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22388),
            .ce(N__19934),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_1_1_LC_12_14_7 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_1_1_LC_12_14_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst.dir_mem_1_1_LC_12_14_7 .LUT_INIT=16'b1001100111001100;
    LogicCell40 \b2v_inst.dir_mem_1_1_LC_12_14_7  (
            .in0(N__23200),
            .in1(N__23023),
            .in2(_gnd_net_),
            .in3(N__19961),
            .lcout(\b2v_inst.dir_mem_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22388),
            .ce(N__19934),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_4_rep1_RNIP76I_LC_12_15_0 .C_ON=1'b0;
    defparam \b2v_inst.indice_4_rep1_RNIP76I_LC_12_15_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_4_rep1_RNIP76I_LC_12_15_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst.indice_4_rep1_RNIP76I_LC_12_15_0  (
            .in0(_gnd_net_),
            .in1(N__21232),
            .in2(_gnd_net_),
            .in3(N__20482),
            .lcout(\b2v_inst.un8_dir_mem_3_ac0_9_0 ),
            .ltout(\b2v_inst.un8_dir_mem_3_ac0_9_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_6_LC_12_15_1 .C_ON=1'b0;
    defparam \b2v_inst.indice_6_LC_12_15_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.indice_6_LC_12_15_1 .LUT_INIT=16'b0000000001101010;
    LogicCell40 \b2v_inst.indice_6_LC_12_15_1  (
            .in0(N__20577),
            .in1(N__20826),
            .in2(N__21269),
            .in3(N__21261),
            .lcout(\b2v_inst.indiceZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21884),
            .ce(N__22946),
            .sr(N__22920));
    defparam \b2v_inst.indice_4_rep1_RNICTP21_LC_12_15_2 .C_ON=1'b0;
    defparam \b2v_inst.indice_4_rep1_RNICTP21_LC_12_15_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_4_rep1_RNICTP21_LC_12_15_2 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \b2v_inst.indice_4_rep1_RNICTP21_LC_12_15_2  (
            .in0(N__21233),
            .in1(N__21173),
            .in2(N__20899),
            .in3(N__21086),
            .lcout(\b2v_inst.un10_indice_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_7_LC_12_15_3 .C_ON=1'b0;
    defparam \b2v_inst.indice_7_LC_12_15_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.indice_7_LC_12_15_3 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \b2v_inst.indice_7_LC_12_15_3  (
            .in0(N__20578),
            .in1(N__20872),
            .in2(N__20953),
            .in3(N__20827),
            .lcout(\b2v_inst.indiceZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21884),
            .ce(N__22946),
            .sr(N__22920));
    defparam \b2v_inst.indice_fast_4_LC_12_15_4 .C_ON=1'b0;
    defparam \b2v_inst.indice_fast_4_LC_12_15_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.indice_fast_4_LC_12_15_4 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \b2v_inst.indice_fast_4_LC_12_15_4  (
            .in0(N__20755),
            .in1(_gnd_net_),
            .in2(N__20831),
            .in3(_gnd_net_),
            .lcout(\b2v_inst.indice_fastZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21884),
            .ce(N__22946),
            .sr(N__22920));
    defparam \b2v_inst.indice_fast_RNIJK54_3_LC_12_15_5 .C_ON=1'b0;
    defparam \b2v_inst.indice_fast_RNIJK54_3_LC_12_15_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.indice_fast_RNIJK54_3_LC_12_15_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst.indice_fast_RNIJK54_3_LC_12_15_5  (
            .in0(_gnd_net_),
            .in1(N__20754),
            .in2(_gnd_net_),
            .in3(N__20722),
            .lcout(\b2v_inst.un8_dir_mem_1_ac0_7_out ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.dir_mem_2_RNO_1_6_LC_12_15_6 .C_ON=1'b0;
    defparam \b2v_inst.dir_mem_2_RNO_1_6_LC_12_15_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst.dir_mem_2_RNO_1_6_LC_12_15_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \b2v_inst.dir_mem_2_RNO_1_6_LC_12_15_6  (
            .in0(N__20665),
            .in1(N__20576),
            .in2(_gnd_net_),
            .in3(N__20483),
            .lcout(\b2v_inst.dir_mem_2_RNO_1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_Clk_Count_RNO_5_6_LC_12_16_1 .C_ON=1'b0;
    defparam \b2v_inst1.r_Clk_Count_RNO_5_6_LC_12_16_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_Clk_Count_RNO_5_6_LC_12_16_1 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \b2v_inst1.r_Clk_Count_RNO_5_6_LC_12_16_1  (
            .in0(N__21658),
            .in1(N__23921),
            .in2(N__23346),
            .in3(N__23835),
            .lcout(\b2v_inst1.g0_i_o5_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_SM_Main_ns_2_0__g0_1_4_LC_12_16_3 .C_ON=1'b0;
    defparam \b2v_inst1.r_SM_Main_ns_2_0__g0_1_4_LC_12_16_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_SM_Main_ns_2_0__g0_1_4_LC_12_16_3 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \b2v_inst1.r_SM_Main_ns_2_0__g0_1_4_LC_12_16_3  (
            .in0(N__24014),
            .in1(N__23920),
            .in2(N__23345),
            .in3(N__23834),
            .lcout(),
            .ltout(\b2v_inst1.g0_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_SM_Main_ns_2_0__g0_0_LC_12_16_4 .C_ON=1'b0;
    defparam \b2v_inst1.r_SM_Main_ns_2_0__g0_0_LC_12_16_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_SM_Main_ns_2_0__g0_0_LC_12_16_4 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \b2v_inst1.r_SM_Main_ns_2_0__g0_0_LC_12_16_4  (
            .in0(N__21662),
            .in1(N__21479),
            .in2(N__21362),
            .in3(N__21561),
            .lcout(\b2v_inst1.N_29_mux_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_SM_Main_RNIAP3K3_2_LC_12_16_6 .C_ON=1'b0;
    defparam \b2v_inst1.r_SM_Main_RNIAP3K3_2_LC_12_16_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_SM_Main_RNIAP3K3_2_LC_12_16_6 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \b2v_inst1.r_SM_Main_RNIAP3K3_2_LC_12_16_6  (
            .in0(N__23497),
            .in1(N__23739),
            .in2(N__21355),
            .in3(N__24015),
            .lcout(\b2v_inst1.un1_r_SM_Main_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_SM_Main_ns_2_0__g0_1_0_LC_12_17_0 .C_ON=1'b0;
    defparam \b2v_inst1.r_SM_Main_ns_2_0__g0_1_0_LC_12_17_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_SM_Main_ns_2_0__g0_1_0_LC_12_17_0 .LUT_INIT=16'b0000011100001111;
    LogicCell40 \b2v_inst1.r_SM_Main_ns_2_0__g0_1_0_LC_12_17_0  (
            .in0(N__21477),
            .in1(N__21542),
            .in2(N__21666),
            .in3(N__23831),
            .lcout(),
            .ltout(\b2v_inst1.g0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_SM_Main_ns_2_0__g0_LC_12_17_1 .C_ON=1'b0;
    defparam \b2v_inst1.r_SM_Main_ns_2_0__g0_LC_12_17_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_SM_Main_ns_2_0__g0_LC_12_17_1 .LUT_INIT=16'b1000110000000000;
    LogicCell40 \b2v_inst1.r_SM_Main_ns_2_0__g0_LC_12_17_1  (
            .in0(N__23314),
            .in1(N__24005),
            .in2(N__21299),
            .in3(N__23913),
            .lcout(),
            .ltout(\b2v_inst1.N_14_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_SM_Main_RNIVAI26_0_LC_12_17_2 .C_ON=1'b0;
    defparam \b2v_inst1.r_SM_Main_RNIVAI26_0_LC_12_17_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_SM_Main_RNIVAI26_0_LC_12_17_2 .LUT_INIT=16'b1110010011110101;
    LogicCell40 \b2v_inst1.r_SM_Main_RNIVAI26_0_LC_12_17_2  (
            .in0(N__23599),
            .in1(N__21296),
            .in2(N__21290),
            .in3(N__23740),
            .lcout(\b2v_inst1.un1_r_SM_Main_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_Clk_Count_RNO_8_4_LC_12_17_3 .C_ON=1'b0;
    defparam \b2v_inst1.r_Clk_Count_RNO_8_4_LC_12_17_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_Clk_Count_RNO_8_4_LC_12_17_3 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \b2v_inst1.r_Clk_Count_RNO_8_4_LC_12_17_3  (
            .in0(N__21543),
            .in1(N__23598),
            .in2(N__23484),
            .in3(N__21478),
            .lcout(),
            .ltout(\b2v_inst1.g0_0_i_a6_1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_Clk_Count_RNO_3_4_LC_12_17_4 .C_ON=1'b0;
    defparam \b2v_inst1.r_Clk_Count_RNO_3_4_LC_12_17_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_Clk_Count_RNO_3_4_LC_12_17_4 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \b2v_inst1.r_Clk_Count_RNO_3_4_LC_12_17_4  (
            .in0(N__23912),
            .in1(N__21284),
            .in2(N__21287),
            .in3(N__23830),
            .lcout(\b2v_inst1.g0_0_i_a6_1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_Clk_Count_RNO_7_4_LC_12_17_5 .C_ON=1'b0;
    defparam \b2v_inst1.r_Clk_Count_RNO_7_4_LC_12_17_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_Clk_Count_RNO_7_4_LC_12_17_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \b2v_inst1.r_Clk_Count_RNO_7_4_LC_12_17_5  (
            .in0(_gnd_net_),
            .in1(N__21639),
            .in2(_gnd_net_),
            .in3(N__24004),
            .lcout(\b2v_inst1.g0_0_i_a6_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_Clk_Count_3_LC_12_17_6 .C_ON=1'b0;
    defparam \b2v_inst1.r_Clk_Count_3_LC_12_17_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst1.r_Clk_Count_3_LC_12_17_6 .LUT_INIT=16'b1001101000010010;
    LogicCell40 \b2v_inst1.r_Clk_Count_3_LC_12_17_6  (
            .in0(N__21643),
            .in1(N__21747),
            .in2(N__21278),
            .in3(N__23455),
            .lcout(\b2v_inst1.r_Clk_CountZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22251),
            .ce(),
            .sr(N__24094));
    defparam \b2v_inst1.r_Clk_Count_RNO_0_0_LC_12_18_0 .C_ON=1'b0;
    defparam \b2v_inst1.r_Clk_Count_RNO_0_0_LC_12_18_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_Clk_Count_RNO_0_0_LC_12_18_0 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \b2v_inst1.r_Clk_Count_RNO_0_0_LC_12_18_0  (
            .in0(N__23704),
            .in1(N__21766),
            .in2(N__22689),
            .in3(N__23608),
            .lcout(),
            .ltout(\b2v_inst1.r_SM_Main_1_sqmuxa_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_Clk_Count_0_LC_12_18_1 .C_ON=1'b0;
    defparam \b2v_inst1.r_Clk_Count_0_LC_12_18_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst1.r_Clk_Count_0_LC_12_18_1 .LUT_INIT=16'b1111100111110001;
    LogicCell40 \b2v_inst1.r_Clk_Count_0_LC_12_18_1  (
            .in0(N__21531),
            .in1(N__21748),
            .in2(N__21752),
            .in3(N__23490),
            .lcout(\b2v_inst1.r_Clk_CountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22461),
            .ce(),
            .sr(N__24092));
    defparam \b2v_inst1.r_Clk_Count_2_LC_12_18_3 .C_ON=1'b0;
    defparam \b2v_inst1.r_Clk_Count_2_LC_12_18_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst1.r_Clk_Count_2_LC_12_18_3 .LUT_INIT=16'b1001000110100010;
    LogicCell40 \b2v_inst1.r_Clk_Count_2_LC_12_18_3  (
            .in0(N__23823),
            .in1(N__21749),
            .in2(N__23498),
            .in3(N__21732),
            .lcout(\b2v_inst1.r_Clk_CountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22461),
            .ce(),
            .sr(N__24092));
    defparam \b2v_inst1.r_SM_Main_ns_2_0__g0_3_1_LC_12_18_4 .C_ON=1'b0;
    defparam \b2v_inst1.r_SM_Main_ns_2_0__g0_3_1_LC_12_18_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_SM_Main_ns_2_0__g0_3_1_LC_12_18_4 .LUT_INIT=16'b0000011100001111;
    LogicCell40 \b2v_inst1.r_SM_Main_ns_2_0__g0_3_1_LC_12_18_4  (
            .in0(N__21453),
            .in1(N__21529),
            .in2(N__21691),
            .in3(N__23822),
            .lcout(),
            .ltout(\b2v_inst1.g0_3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_SM_Main_ns_2_0__g0_3_LC_12_18_5 .C_ON=1'b0;
    defparam \b2v_inst1.r_SM_Main_ns_2_0__g0_3_LC_12_18_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_SM_Main_ns_2_0__g0_3_LC_12_18_5 .LUT_INIT=16'b1000110000000000;
    LogicCell40 \b2v_inst1.r_SM_Main_ns_2_0__g0_3_LC_12_18_5  (
            .in0(N__23313),
            .in1(N__23990),
            .in2(N__21581),
            .in3(N__23917),
            .lcout(\b2v_inst1.N_14_0_0 ),
            .ltout(\b2v_inst1.N_14_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_Clk_Count_RNO_4_1_LC_12_18_6 .C_ON=1'b0;
    defparam \b2v_inst1.r_Clk_Count_RNO_4_1_LC_12_18_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_Clk_Count_RNO_4_1_LC_12_18_6 .LUT_INIT=16'b0000110000101110;
    LogicCell40 \b2v_inst1.r_Clk_Count_RNO_4_1_LC_12_18_6  (
            .in0(N__23703),
            .in1(N__23607),
            .in2(N__21572),
            .in3(N__21569),
            .lcout(),
            .ltout(\b2v_inst1.g3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_Clk_Count_RNO_1_1_LC_12_18_7 .C_ON=1'b0;
    defparam \b2v_inst1.r_Clk_Count_RNO_1_1_LC_12_18_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_Clk_Count_RNO_1_1_LC_12_18_7 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \b2v_inst1.r_Clk_Count_RNO_1_1_LC_12_18_7  (
            .in0(N__21530),
            .in1(_gnd_net_),
            .in2(N__21482),
            .in3(N__21454),
            .lcout(\b2v_inst1.g3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_Clk_Count_RNO_5_4_LC_12_19_1 .C_ON=1'b0;
    defparam \b2v_inst1.r_Clk_Count_RNO_5_4_LC_12_19_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_Clk_Count_RNO_5_4_LC_12_19_1 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \b2v_inst1.r_Clk_Count_RNO_5_4_LC_12_19_1  (
            .in0(N__23365),
            .in1(N__21386),
            .in2(_gnd_net_),
            .in3(N__23294),
            .lcout(),
            .ltout(\b2v_inst1.N_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_Clk_Count_RNO_2_4_LC_12_19_2 .C_ON=1'b0;
    defparam \b2v_inst1.r_Clk_Count_RNO_2_4_LC_12_19_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_Clk_Count_RNO_2_4_LC_12_19_2 .LUT_INIT=16'b1111011111110000;
    LogicCell40 \b2v_inst1.r_Clk_Count_RNO_2_4_LC_12_19_2  (
            .in0(N__23295),
            .in1(N__23489),
            .in2(N__21377),
            .in3(N__21374),
            .lcout(),
            .ltout(\b2v_inst1.g0_0_i_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_Clk_Count_4_LC_12_19_3 .C_ON=1'b0;
    defparam \b2v_inst1.r_Clk_Count_4_LC_12_19_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst1.r_Clk_Count_4_LC_12_19_3 .LUT_INIT=16'b0000000100000011;
    LogicCell40 \b2v_inst1.r_Clk_Count_4_LC_12_19_3  (
            .in0(N__24113),
            .in1(N__23225),
            .in2(N__24104),
            .in3(N__24101),
            .lcout(\b2v_inst1.r_Clk_CountZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21890),
            .ce(),
            .sr(N__24095));
    defparam \b2v_inst1.r_Clk_Count_RNO_6_1_LC_12_19_4 .C_ON=1'b0;
    defparam \b2v_inst1.r_Clk_Count_RNO_6_1_LC_12_19_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_Clk_Count_RNO_6_1_LC_12_19_4 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \b2v_inst1.r_Clk_Count_RNO_6_1_LC_12_19_4  (
            .in0(N__23986),
            .in1(N__23914),
            .in2(N__23320),
            .in3(N__23829),
            .lcout(\b2v_inst1.g2_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_Clk_Count_RNO_4_4_LC_12_20_3 .C_ON=1'b0;
    defparam \b2v_inst1.r_Clk_Count_RNO_4_4_LC_12_20_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_Clk_Count_RNO_4_4_LC_12_20_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \b2v_inst1.r_Clk_Count_RNO_4_4_LC_12_20_3  (
            .in0(_gnd_net_),
            .in1(N__23706),
            .in2(_gnd_net_),
            .in3(N__23624),
            .lcout(),
            .ltout(\b2v_inst1.g0_0_i_a6_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_Clk_Count_RNO_1_4_LC_12_20_4 .C_ON=1'b0;
    defparam \b2v_inst1.r_Clk_Count_RNO_1_4_LC_12_20_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst1.r_Clk_Count_RNO_1_4_LC_12_20_4 .LUT_INIT=16'b0101000011111100;
    LogicCell40 \b2v_inst1.r_Clk_Count_RNO_1_4_LC_12_20_4  (
            .in0(N__23488),
            .in1(N__23366),
            .in2(N__23354),
            .in3(N__23301),
            .lcout(\b2v_inst1.g0_0_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst.indice_1_LC_13_16_0 .C_ON=1'b0;
    defparam \b2v_inst.indice_1_LC_13_16_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst.indice_1_LC_13_16_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \b2v_inst.indice_1_LC_13_16_0  (
            .in0(_gnd_net_),
            .in1(N__23218),
            .in2(_gnd_net_),
            .in3(N__22996),
            .lcout(\b2v_inst.indiceZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22500),
            .ce(N__22945),
            .sr(N__22922));
    defparam \b2v_inst1.r_RX_Data_R_LC_13_19_2 .C_ON=1'b0;
    defparam \b2v_inst1.r_RX_Data_R_LC_13_19_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst1.r_RX_Data_R_LC_13_19_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst1.r_RX_Data_R_LC_13_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22772),
            .lcout(\b2v_inst1.r_RX_Data_RZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22252),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst1.r_RX_Data_LC_13_19_6 .C_ON=1'b0;
    defparam \b2v_inst1.r_RX_Data_LC_13_19_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst1.r_RX_Data_LC_13_19_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst1.r_RX_Data_LC_13_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22757),
            .lcout(\b2v_inst1.r_RX_DataZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22252),
            .ce(),
            .sr(_gnd_net_));
endmodule // anda_plis
